// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:39:48 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PABySiHwTd8qa+FnSDCSyB5XZ8shcAaKYwjff9HmZcu7lPWWg1vkNTbjVHazJGaf
4KahEnv/MjV1cJ+uepDR++Q7JT/kKRQvfnDc+6BPQVrSKRofvKNDwGzLxpuo6Zfp
/i9wGlPP2xy5IZdDq6hc2Yx/bs3LWSrwUuuT9I+hfGE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28704)
O6eG/NtLFz9s3N4FDWXH8GB7f79PMnuwYwQG9poxADJr+naO3IdGJCIajJ6wxWW0
ZhUveNN2vtA84JfUWgOT+EPY3Yfx1EPW44vMXBgEQ2XDTdxALF2S/509kkD5Fjsm
mCFsvUag73waxAgnOcOiHCkD1/N3cGie9JRAndWCLxyeAHw8XRWxIxc8Og4xSVz7
HocZ629mRkEJvEij1U4VzpaaJy0x8QFys1oIDoDjD503AgQQvORE7WjBycslft06
sPJ1hDG6W1pu7///3ogGqHW9WtjoqVNzaTFvWE9QWanbTAzHTwKSP9vq8lynX6L0
993Rvcax5eHcnILlgpQ1Si9SUO/kdelKQFXoLd6gzfCLNN1Xy6rn10sfLxbdk9lo
eE2DZ1EFqNqoHVQQSFgqxjk+ZY43N/g2vlyn4i1tZ4LIhxya1piBnUrUgZpFu0tF
fZk/TP0Y/DPM3rivEgmpib2Fe4FUA/WfIYVnCoIunWGc7DFvCBYWKISfXUZGLwJm
e2EpoQPkAw1dfe5LWvAWtJLEtKJxYbX85Uw5MXh616NkcFa+gpCDG+2FmlFtWViM
VCrkTfyaA5MolJjXv5Wi6rYLMks8j1YjulbyickedSZN4NW76GoML3AIILx+cWpy
KW2/7/x4q8g7UuVw6r1VKrf9XFpQMyC1URX4johqV2TAY9/edBucDC3CIKeT1xdI
2jiaqnZicn5Ce3L8wDBSy97DQdP5fm2TnIJYGMswDnKxu2jjK/N2L0XE5VhIbkbw
0sBnOSV206DVKYRS/Z1UJMjXWtsGFpLAZUEKQJm4GRscEkOyx8a709vW1cFqNpt2
EzxmtFOIe6gqR5mWQOD5y7Tpph/Hl9LYTd7xhVdLSfwcGdY/EqQENJZa8dzJAJP7
JVqBrL5WVz1/74RQqUwgxS/X9EcVXjllYj+MsPRuSciNSthFqis1NoFGcnPdYheP
mXIPkrrfdW5TRLW56DnHroI+whLE8Y11iM9/8MDjiS1XN6RQOTMNA6yQcuyo1Qha
kF7Qo0M1ZwQlQG+3ablt2aBodUFCfGVnPtnc7/8BHfyTg84EVUXCdDswXY43jKHT
FeYsqqVIGLYeUMY+X23WoSMPo0SZ+JjHklM/YFefuzDmF/ZOjCur5KqJHUYLNDu/
df/hVzQus96if1TIEXrKGgS+bXpjHRfxgDjo3+7mLOqB8rvF4Xxqy2hbX6t6sZu9
BLno/by/PeZDUu/OsHdzFzkn5sVBlcThCQ6xeC7Gpxs1qm3i1uXNcfCT4FRO5MFK
BgCOcZZzSQfEYPYhaTvKS648e5Ii5/+VGXqW+6ct91t47iAlpMRoO6wjjKZ+Y4yT
p7gEJEk5XnZl5VtPzDep/6Imk5bT2J9whUUsCGvnm4uWR5OyUqx3+yUX38L/SPT4
aD2bXr0Hs6t3itY/Onp/DHwFdKtrOYStKCHcvtWiqJgRxVh3pjTkP9aDrRJVX/go
WH4JALw8qp+cYIekntE0Vc8096VxeRp1EP1I6MicDquRXEa4ABI+VKf9ZN7SvKdx
JVaixLaaddtT0A9pkiwWIyh7VyM8TySnSA58RqzfMH38WQRSgRvGWZBsjWhK42HJ
1jtXzzBWNSUOweJGLjVi83Yioltgp6BtyK4qgWCqTE0BfKTJHj9QiR4YxgIU9BQS
7YDIPinKgijHQXSJEsq5nALWKF7Ygsp45+RDWDxvXDCbBQxHMOJ5ZvRFIT7m7zxN
kPwckAbYkGhGzGKt54yDRVms9O5hkAyO1bIsI0O26TXXmHTvjPoAceOcr7YEP9gN
vB7KeThdEsD2Tt1G+NPq5Cl64BsD16c/1ULQ6id4NDnw33j+HG0W5Q5xIO/O0tUo
qjIJxL4txrya6PRF1n4oeKBpL9E9fY1zEZFtYM+JiKiKlJDLFo4tDRwxAGffPwnA
PC7tPLodhGW7TRt+GrEIFtNZW+f/k8Yd/DXo/nvFeSAWzuw9cmLaKlS0jwxG5q2Q
bID5kQ9Zp2vwqBxuBszxPkEvncHn/LdxTgbaN+1Q9+cA29vGAYgMqZNKPYjiZAlP
MI+F9jKuUlig1j4XqRM4pMcnI8CPwRRT+/NloanC+N3RDZj1U+VYIS9dMHEl7FXK
WtUJv/URad+/BF8tS8V4ckNOXiKT00KA8gMjADXPvPzypXHN6LYUq0BUPurO37gb
p14C++AVJo6LIVvEZqMDmwtHMcdDf1N7zb1sKkAXFSGCIm0RZU5hJOwUacHZZadc
0bA4ltBaWhGmC/t2q5k67UBu/zok+Tkdmzi1EViYoeU/w8kfV+IEPVUvY09zpWLt
Jw+C9OA6oI/g0gX+ZS7yKrhi/hBjTg1vrS1zcp6zFtBPCYuhMH2sHGJBaylqtBGV
iaWnJFsBa1iBwzVHjJyEfYT8mzLtZ+Dd6Um0a2qZtHE3tXeGtiJ0a+g8wl7t5TD+
hKYsjFP1G+x8jOw07LGC1O2cimr77cNl+L53VQe5ElfeyRpMw384ISgj84+Dq+dz
BxTIf4F+PBcVIzBh+ZsqlK6sT9GDjSAgI+kYssVG3PL43Dp2feIXpvZEFZEL24rF
GFvNYHUHCQvYvkmU/oz36bgo4R/iZ26byakuONZL+Zo5zVGfT+sY2ED9SMxG7eYv
rroHZp8K2GA27IatGiUQ+1Vy2c1hIIywkxus0Xu6JGdhK5zCvq+9ULWcugvY+60u
He8x2WofMANKFprRFai9tToFZXGtzywBh5eoiAX2msgeuaOpcRAVGtyhjosF/RxA
g6oa+UryDLIywiYfwjRZrzdTclwouzVjNl4Vu23VrUlhN5t9k76AH8Jb+8QHuqTK
14tJPRu4reHCwYxBw+s8BUATxi+y2+PzVjb35mVLeN2REFvCcHtgJSzglkk2YqbF
T+8USch70Y6TdI5zCirsFqoWVVmpPWnryHJR1mPzsZlsNwLzoY1DINRBa9+SL2Bi
e5Rk9OO8/pMXrVUtxlO5wy4QEMHYqCNzlnOnxqI0L6IuWtRR4yMfpGHCHn+i+v9k
royMSP9RWXpsz8xayxdzGtuGCFsOXuS6wng0KBdmlFemGlhEkltMyJQ47oNQAdzy
AHyzTJxUKXZ2Blxxi9AXZcUpppTROyuEOuJIiPeqT4SXmyTWX459DP2IZOuJrzOb
iMCvbA+IFIAahWoYFpk2OL242tLr1I9mqPOlG6U7bnlJqReH2TWukYhaObtog7lG
7XnBuNuVztJydLY2jtnA8/J1zBCyDQyynJVC7HFROSrcx1U0g0VDkQgICsP3sB7/
npqKgS0YJ48Q09ZD19GvLILp0HQc8iAyBZm4iCEmyus+KO14b6d1KmvVIx6Sh0X3
9Nl/hin/49D77wu3syiCFzwk8JsdEjntRGK4hzRg7GH57oKxVmWVB6c/RJ4swGuG
xdNUrGDYPS+dm8BpgAYrM+dk2rI/JOPBsfEiNXubCJGt2VtIh8ab+b9AeSg4VlQa
XiViPv7bl83RDIzWBaNlqAFUh1aKlwUVCNF3UjNgf6WI3+yb+BQzx5dSRnAJMNPA
Q4fmjlfWi400HCARhh7CJrmi8Wt43RBwh9Mrjdp88lqVRWt/b6lvuq6K174IW2S/
y9CTRsCY7SNfM2TG/QWozu1my+i8TSodafcvRMDMQ83W/OD3udslAobKW6XzXDHE
SKD4esrRyE5hhgbBIqhPqDiEEb8spfHSIx0tI+/4cJCei43vxWqZl5/WHtUcKnk3
NphTngfgt2K6xMCBv7rLnJYPGW1BlD2VfUUY/BFHbgJcbBzaF99sDJiUvLVWuAm2
nlUdMIo8xf5ITqNNT+PZsK8lsktQCTctR1NfXaMO2PaD3jmw0ztIE9SxEvnoWHoH
v6xMZBBbN5/Yw2fbjiWhfafb1REwQghVQqFMwzGwEo4UaigAeb5T3GRzBwB/p3Y7
rb/A7fic/n6fu9mDt1JScKWN/8I2tQE+xbIbUKb38iJMV0XDYgFfcXfblFxkQKb5
UeYXSutfuGx28cp+N86QuJh0qXoLIIYRm2CeEPERVGIoDXXTIYbWepiAbzYZpWyB
GrUzpMJz01/qQReGbxXeMKe8z6tWesoSY7WPVfycbXZ+PNDM9LDg9tcL0byf+Jx8
6dFYNq47CFN02HnABkL7t4Eg8uoCoI6/nf9CQSe0F8l6nzwGZXu4ePxBjYO7c5Zd
kP4DKTOHLvEZTwRdLQfl3snfA441yhaLtjSoH4qNTMRum2nr2o47BC2Kgl06ee13
rtuchLcMBP6flctjdbva8ex/y/yaLoqGLbhEPYwIkIaR4Qn0HB/A+j2h8SVJwM3e
9tb8kbnQMKtnaJWlXxMcwiBtyrKomkWbRwT/cMOOldvdgxeeVMvGz0sfe6HxJ/1V
kvg7+3qut8/ot5fqD9AhNQ1LJ2hQXLBHe6CVP2EWCj2OCOMAJ5Vy34jZFeaRSi5U
ELbsb9NhS70EwPvFcC5/XsZECGyZHsD5mgQoYKDP1e0ZOXnkoirN8blCwrPLDocB
qlCpEmwg+SstwxIK9OJ3+qOnjnrrlx1rNk7VY0Lx985jtvRBwB6ZyM8nBVXL3NdN
oZ5P/1ES4FXgcFTOMK+lr9stHwB5C6qfpTi+hB7fCRlBic9YRN5gxOZe1JQwxT9X
Fmx9aHA44DXj+R4KPXK6b6zsvHdd1VHxy+HVK8dyht+g6k58rn/+Tzub8Kmcb9Ln
YLgeKXjDTWI28Pxto7RoFYg779XCHNLoSs/0nMjEbO6Q2ktxnljnPONXSsibMnm7
nx11VtHoJK9sweGzFBAN80IvEioHVBVwVeooF98ZOAVk8yPa1vXCZC8nJgxDp79+
wge47Khkst5xRzOa/EwyUQuwEMFJgju03gcJFmUVJX+nlHmndKN9XauUH/xGUAZ3
jvz1QydiKFCcIFJCmTF4x2WyGSxa3RB6Y20azNWIdUOxkOPgBwVfpErdCdGu0zIr
0jOhOOJOoxw/ZGxtNz/nQBTC3Obr3s2JIyvpQ9ZP8OTznpi/u0r1WfLnc6GoTcxj
0LE7A0M8NQHIRxy2iT0fFbuvUGyzmJTIB3qLKSEJw/xDQu+OAHsGGluriTHQ3LpZ
T4jsVAxmo4RJRdcROwWoz2p/MgH+eCPLHJqmLitXlX6NWGZzri83tlqfq54+7wrE
YX7K1TjMkEaC3QipAC/+ItMRAgGTs+OriMkzk1Va1eGynKw1CKrjQiUc+ItwiDiT
bZuRtEjPBOCevyJGrPbcgKYl0NhdYkkyWDPvnnod+/0NhOfEX5xx4xefvEs8qVCg
pDlRGKzjOrToJUUfdLsZsDHehWFEQTNxJ8tS+BGdnktlCoYtTNR0OQG+Y7l1sW5t
05BDCsttxqQTs3ETynbXtCaJD7HDhvAlkNom8ocCn4UWo2UaO+YVShDMmJeIt+h4
q9kvoLvP43VdOvj3CcHAUkUviEqrLn2nRx5BcURXg1MiGcJBLQY3WQpKMMab22Nx
wD+omyh//mfSSidtLvyXKICJpS38ySDEi4HDcW0rftXIJGZURGSTh228qJdK925o
82xCMZK5LYNnT8RzoUZ6UmzlXYN/iZVcs9qXfNSDdW1GIGjyiXt+GXomCvj3RGrb
6j9yJH+MqnU4J/c+mD4mh13fUjxo7VsWyBNCmvTuc5ROmOK6n/WPJz95PN3BKBBs
gpv3slZiLPkO1pffzasQC+YNdE6dQFBXJeNK4D/HeqYWQrrAnf+vSwjZpVc46kgD
vVzHHim8VeUwdULza0oM0aSTtfKwrr4CTDnXUIEiQQhF2ooZWHnSYIks5KG791Z6
eRhzrK2Gdpbo6Bzqdyjz3ky1we7g4S92jSMY1h/c2GkaOcmS4ytf9KbTZo8XTK4I
Q9hYITm+q2dksAJASZuRs/aMjzFCe8getgAu6X6Dziv9egpnWeChqTIrFvTPkC+P
mvjl+A7s3IWMuWNlgeBaP0+svn0AEq5lls6AVWPwH1czCGkiwxhDjyo8juUQ/LXx
y+w58k8FbFSXobOC6oDA+eHFl6HK4L4bcxEWErJv5j8TFPPhuKg6qGIKgQhk52p7
s4flv17bNa/kGE1ZNQ88NCCEcI+0UavviS+kwEH1d9mUUE6MxbSWkdjj6oC7Wser
T3yq3ohEqWzbjjKz+7f7EwrHgmoKJoaL+zRWm8OcSLhUH9AT2pAUB3yVfS0xNW+c
nPm1FrskryHQbJcHdP5g5VGXH51h7tHVbN9FK1PISiouy3nBMxws3sbVM4UtLd9z
u9J7Szhw9Kt3iPe0WVlHUGwDt2AegB9u4aXLkrsw5pUQpPPWNdWk1yDd6ba4YVIR
Sfqt6+kpZl/b8ygRQ0H0QOyKxzi+IgJMlfBkMnwQdBvE7poxH1aZKdedUAcfSHTd
+MFje3DMwG9o8wwYWd9xRMPp+iICpWCYVKQB4aPg+7QMUI5majpOLuMQfQ+H4XlA
H6Z1TmrJr8B7zY9FGwO3PnDaPdjWnp5Wpn/KvJBkisEKV1NQ4bjQFOhkwgI7WcSX
DZEXTY1woQ3k5tkh4l+VXXWdGDlZNPOsotO6jqbG5emCctUJnYXAHGSZmzTDC80+
sTrHsvEvehdeLGG4PwUgmBaP6c7z+l7z1lS46Ztcdp9Cka0j3SmmvULkBrqxlcW6
4Fg0G4nmJPX7xa1AiRXQTefblv07zioaBCbzIlE+CFEAUM/QxbP8++PfSxOTQrKZ
zrpLYckC7l7AbAcjMUT22FlGOKlA9zrX8CSIraIMwfYnPYEeP9Zc7jWbPi8GALbd
haWWQjk1gzijjw45TUTkedRwpZFF1X0RudiiAPKPQ6cmo4cZlSvpDehk1MGOkUIH
ZzOxNEL2jH1mjiE3nkTbeHLdNKR9nS3aDI7PlnceLlLj1WkDFie9pdqu935xue+4
jA4wNCOzCzjEY9foR+RGUHcf7AxTJlMLKCnYXLwB4uL5YW2achOTs8p/hFHv4cW2
91mrAwdEWmASDgVSgw1bS9210ZDYdoL7DRD5XS8U/6AcK4BOmCV245cyCAc7Jasz
yKnraz6og8IhvEPjDHeVu47kXcIF3sX7sMqAOApUKuTRjfdMAgpi2+vZfoNcU27c
Zigmm+5M06WS94/m1Cao5uo25Y/BB2fgi+fgo5uB+Fhv3DngsmWP0ZNyd0TKsPVC
t+QUgkN2GJnRCcFeoVFMjxmzbE/jX6Y0vKrBzBvlzbk4kXB7ZC9eqMyum8lNmUbN
M1XiWpsMY9ii/J1WR2PkmM+s5NtK1ZWtQbJcxOTC/k1039dsgMd5C+7elnlrvQOe
Gmw+NCon2Cz2LtoYywejvT1HiW+U3d4oQmE0tod4r+UCNnOTjQF8d2JI4Cqq9MEI
6F4LXUKT9Eqvacj8kNh9+xk8bK8Jb0Gf58tDJwe/IDVZGiBdDDeg1JHk2vIIUFuD
xX8gfz8QBWRDJ8AJODMECA8FMvXVQYibYX5i6bftppgWBcv+vZiOyKLrY4535SJ+
ePKLcwruooph1tHmmz/ZEFH00bqDcZUM5IRtmIbclvuYVOCZys0zL1mXFjSGON2i
TwKkfkLnzf3JHRTT6D55vQdM4RKSw14IDODTAikG+d0d3m7KpobDx1YxVWaWl12Z
ap9NgPueMocjhRcUVs/eYNM6jlk7otPI888Kj9VBk5LhpTnB2uATSaYBg0WOozaf
5crBat4AyJlaLK7jaAeEUuZYlKlPklrSKpITtupd+UJk25kgUzI68vJcgARUJqTc
CR6aOnxWnMRxa72SB9wtpHBkjL0a/K/CJO0svEVIhIR9W4TmvlxjQtVNuZ+oYfn+
otFigjJ0N6m3wO378BtGo1H/CW186TfWE1haHpQUwLzd7ayRyP1x8L6upbXLVIAu
XH7GjyfJZdMBIVBbJWv1U1J/H853lzzMscrd8h+SCiGpRP5o5UiX3zewNo6Z7WFM
q0Cdi/n6R3oq6/9dHjaBYKbFbjHuaIKu1HTx53zccWbycVo/d1xcqza6LwoDN3Tl
FvWWStuXxhz9ui3KE2PF/T8ODc9yPWNjlRMdmt8a9qeK95P5ejKTauoR+NTPMUoa
cRFUm36+hLx08zthj/TMRIJkCtdoFMctwziF61h9v04ul4Yk3OCWxxNdtdLm0/Ii
/qhh2cmctlsnDKKtCDRvy7EEkxo2Zk6nJ+ITojckpbLes0ynzE0uONPawlgUG4QO
lFOPgUeWZ/J4YLJ1NzxbdFUhXgv1/wj1keVFVWzHiav3pRtiatUM96ExOfLZoCk4
E0oIXNRX7/iTjA8iuQUn7wjD6VLg9iUoWhpUEn8jT0Kt5ufU+VWtzzhHARhhD3y3
PwWcIHjXKRqro+FYls2T+2X2uGrjFSaX59CrUIQTr2SpnvlkLEtJxYbrDrVv5Rdm
4wWDFSFvyHKaicjfFf0mLuyrUhDrpz+6TY9IRs03k+tdNqktEYOwTqLkREeua56B
QiINGYeWqPEHUCwt1pPhqiOqrhXeScnbUDSrwEhnhz+1bpopXQTGabZL3AMF6Vab
ChHOFFz8sHPI3bVzLXbJwGCrKURahPG2ooryZBPWJ/0R5RGpRrdEf5/s15Pk9xDm
dIMykqPGnODTAcAgY033iGXb1PtrLaWmZTaSR9G1qJFjxwQlUviz9i4ACMKi+tN9
7YnRJaaEKxV1s7SlgXYjO/I3PwIriZq2LhcWO7Ia3Zt0fD8xAF41X885jok27nIW
X5Jeseas+u7WEUYqFXfEpY1E2A4PWWXDIcjEBbiOvPrWPwfnepDtsiGD3QYLGZWA
S9F61zFK/tFxBb6zpmAVmKUlT8aMSMddE1+2cD8Lb6PvtDnP3RWEmmmev5OE6Df+
VJq/4w+yI4grW2ARxNfGii0tja433wYniFT5OnkhdPzhKoilLxCTe3vwQTcoJNxb
I7bl9HhaNx3kba9OctbbxjURbLkkaRN0j6NNg/yEbegFQEdmBbw3Eqym5CCX/oCu
PYmFDGtyngsu09d9Der4TyE8TfDg/xos1AUrQ33MTrET+1W6WmSVLb012OQZrT6g
kJxLxhlX+wCidiLOZeEsSNynllJq4NgwmQgueFq6bZpUSmdPmULAQA9k1yufnUZ8
LIICOE0mfeaMKH/hXyXUnAO34P4vbnFQNcvsfr3zBu+F3p6pyOA9UyxHZ0LsOEiV
fYl6xKS0ay1a5R3wvFQWbfFAu8KSQKGVTtavTKWuj0IIkSoZC2E2oHdpVO8nnGJZ
HBP0dTFdxCOQBdMTg4I3UGSmpIAIzHxeVuaFn7ieZ4yizzwMgD8N1qyDjKXFmOuB
EGBDvkS9/fkyFBTGwi0YQeO3zdPENZjp06q86OrNuoEKnrpJg+sdGDO53EGf6D7v
3QijTnhUUCEuMx/ffRQjocXgIedMrqhUWTxM9M3K3B9ETAYmDm05n4yGvKUxJj/m
b8Niy6n6eS98gmF0cT98XOWA5260Sn94uJr5P027smVWOumV9b14oQxtJy7gC0X+
R96xe/SJIDnG3p5PkwAMEHaBMocoltww2+tLTBJ5wUEVGltVKpM/BqjYiKBIqgVc
wmLJs+bNJE9jNUiPjDijx2Rg/FyFuI46zqarNDgtcdwz32otgNJyjDY1BJnTVc0y
nUqpn1OEdoFg2A+Ie8U4b4uv9FhdwjYXRRe88QGzD0LcV96AbobXLZRjOC/8UwDv
TOOo+Uoz23fo8w/YXsqJW3RxEWs39uUXPGKehFchv7Q02iGtqVLdBksqrE0Vt9/m
clnLZek7B1tY3s33fd0fc0dw13ThPp41ZMalGGdRUpzvD2Nm++LW38c8KMhclT2q
SQv5hfi2gGx8AlwJWWFI3U4edFw0Ad8SvES7R+GN/RUlM+8laPQIBr4tPPYzFCgC
jVUkvQKXHALOjyXrNkeq7jYqJ8gch27mSBCiESU4z5S+3fdWl6nM1isTvoJ0i9h5
ip9EizUyQCypGixEtAEwraWpGWTg0e6LBe0NSx3iZYC6a7LVYyP8Crvl40IFJIaT
OZn36XkeLCTEWYZ05TPSiYHHU5W53cnKnRMgwxN8XFamHwyW53xP7ywrPmeyPNwL
RGqxol1ai7V1+ShcWIITfLxZC8TqJeZ3ZyRdbvosAwSwA/l+U05uh65DKZ0RF31g
ObcTsVeMcX8C3/x2+onOyZnuozrackKv9995AACGUj0Ulyo54VyESDRiNXV6yFX1
k41BFG72cNr9F+xlYuBksBncLcr4Mz8nulPXJYcS4rBLD8fF8s8D0au8PkMiiPUp
57xWB0VZWcckqYnhEvMADuFCqKNSXnLShXS1z6EhKO1LE0UPcFq63EYzEHI45Sc3
KRR7iqjMak3xQJSxBynMx2hF4mcg+KUH7vhO9xkpYqrvjIuMsvNs6m1VapGekK/d
VuZG3pc0C8V1a+yQZ+ZIXLBv7zXN2vHJE3sObpKfSx+rQ8fGNRZqGpKDnEDvVmgS
g9h4MrIQ1ymiIqeu8JGuvx9flstRVWSqaDbOenmT6f3fEtPE4jqsuepiF4yqhuDl
DA5jE1fajFcuNgMPIEfItI1qoF7W051Fjt1cLoV7h1yQhzBBQf2hYLKa4Bu1jyfP
Lr+6WV9G049wWbPiPu2gvZ16po3XP9BjVo+ll6PjOaMZmW1+9XB3E0rrUxUQuACQ
hp2pYLTfS5VC8cQ1efiU23QxN/hzQ7KRQrSzHidwVLHckifn53rZuvVM/IKE5J1c
GmVjmtZeykYgA4jonJlnGdCgRJ+4zauyDYJ9BdWL7YKg0fGHHSFcHfrwBata0ddG
+kbOKZiIKYGqV5rLKqVTOn2Dm9h7nF+xJ+jZSjdmqtk0r52fM9OKyG2V1KWBqLAL
g4ZvncfF2ueLWSe0NyMTxQ3SF3b5q59M9isYYzjDgDCXbmmInqnIRAiOk+MH/0R7
g+uBmsFLS4nwHoX2Tq/OhKc/GD9CjNg4WmkhjYzs9ntdCoypP9RlCVkdD/dCJWmj
/qqSjmMCoJfBsY1V/LQKZ5Cz57OMy8y+TsLRjIsF+susT04DGbPlVyeMKv2sTJRb
ObVeWoSN8QxT0OcC2uWkFIpoImtmEAhOUzLktr8FykfwiGRS6bVw74SppYKaK9ub
Veci5Pcjd6wKViI0PqjzoLjTGc9Er9oVcXMkZRozIHlAD26F7dx9nR4rJAu6HssQ
U2BsLrZGpy0Mm3YC7uUhqAfE0vUcQAGwe1iItaqJjEQUF501yNL3BdArozqnNBNQ
4B7Jqm6kjeAtvPKWZ/EII9HSZrE7WEnTGyz+h1jEmEcP0HYzfIaYUlR6ZfWKioPn
DYrkBx0oC78xoXyNL8U2TVEEUbbyFtXU8tv3wA36V9YL3j75lnHPLguATwUrJfwY
PuwnJYwh/cpvjffP2oM1UOfXALWv8seKooq/HjjIlEX5nQKLIFVbTFhgKG3RvXkn
Cq06S2Z+burtgAMT0e3ixgoQbEpTsWw3+TjSeVnN05fPORKhJlujSpqKkkPoEDj2
m989JyLLhXtbwS41w6hioDTV9NhRvcDgnNLmyxW2+fHDl/oyPRwKWnbXmZztnKMg
lwXBGd2LVeLxRT682xPpy94VBxJ/5/TE8sbmc02XXQTPOuK/lPKNKzHK+S7sNt/s
Lk5VWZiuBOqnl6TWcXo65FtSZEtm0RxkUnIMfQz7VeJbCos6nccxvxiIyRnRCfqw
TiS4B72b/HqADz5C2PSauT8SV6yAa+aNl0ArtF+X1YGW1izD9BV+UmJCADdj9ErP
6MPDFqyc3kOOoB8L2NRbPlrmkoT1yZl7pkpq4vOOx0weNLHeov6muB81M6eMQlOY
RhT/mnx69VbfcTCTPXvtwHzB4LBwKwqqBm6Sh0yMgRFg2yDTfWZvgf+kV4bfAmAa
j9lxLnVAPdIcVMYsvTser1jt6WbQDrs6EQ/uwfyYDrnaZDuI73rYLxuMKObXo5eC
GJ5WWFLy4q1m96YkBRz3ZwK9+Eii+7Bp/TZdDrIeL08GzZkbaqQ0tkmF0XR8zoF1
AKRPp/xcRkwEQ/V9Z6xB7/pSGR1qSym+GuLcTnJ2K16OuVS+oe+2Ul/Us8hH8O5T
aiepIJ8Jd/VmJs4vwPHRsthM5J6B3t+jpmArJinjsNTwXU1DQXKrMo/GHLnEb2uC
3KTnVgGNSkvamMoJTUmwmRnwmpI9W1wGWcc/jwSKXSOeopMsGSA0/PUrMnGyxYBB
VZoVE7XOL3ZnsZwnswn5eonAV/TvOwlPCB46bgG4LHoaz37J3q1Ny9wGB99S2eFO
/gLqRxBkn/I9fPwR68Xk72rMhwRqS6Xpp4X2UksFGE0h3bH0u2ZJoMtb5Ua91BYj
+47qBCiZRUPVBamtAhhmfq07IL+re0K5Ohf6hRTH3/LlmqMd1w1JxbDRIqVuaFdK
tM25NLEEi6S4tXVx+XnVD6dmde0rYwx0fgWKlaANZKAJ8BKDoC6/ZP4htYGa9smW
odNb6JoAMzM/JXtKKvAI5Agk/I0xb3yLzTi+DZjRhb44qttS7qYTBTyHU2oAM5Vi
eIKdPbo/XQJY8Pr5P5b09oqYtHmrf0T5aiDr6yEk0a5dApaebTIzO04zr8BF3uVe
pZblqIcZjFdv/RirqhcnU5y1flJqEd4d2tFpyiswhwUP+2hrxBqfKvLVA0CzFxj0
eCBVI+LcBGVRsUMZqbWzFwD/FRv3qGJPgGk6y98D2S/9s6q9VMYOT2OfiCHAxe9y
kNO43NjNwxxHnb06TvNPgISgwI4T4wy8yqTnTzwrwNSp43KYPEXIFe3A8d0g5chd
nl1itp6AnB4h3U2hzaUeiK/IDF5rX6zbH2cueetcf8lRLJ3AU5uwwxpEL+INpvKb
Imaxkfp4VGY0+Y0tlwk7QsoMHfRgUSzxV9OKXxBlKIssvicF1f3PiHLUyjAEW5Kn
6mfRzr2LqFJuVphBeesIaLCzmCt7bTCeB8RN6YeqFeQLumIcDgIzkwqzUd+WGAlm
qbdb++DpWeZy9kcB7y8cSge96x8vrmu1UlkHhWgUqY11aXL82XE9WG/4HhJgQTj5
AIQJpE0K/i7i9Xhj0r3Z/LJrBuuW+efZZ+CL37PWicLPxDz+x+SCGeIZ782uN5bF
9rGiCXYWQ29yCXa14tKJ20Hgoc+IaMqNEv8uQeiTa1zQ5Fd6Vh4xprkaZ1sYFxTm
KcuLJuQvnPEMRqWbMAmpjGDR/4NVHAnbggcR8zZkoZIiAB9OdtDBpnEK5krOis3N
mMmwxcx1XcwWxv5iFsB0InJxZW3ej6jql31aZhG858Yq1DFlUck4uBl6gfQqMRct
xH4HnAw5F5R/fyGCUGi9jInuMt6YB3nCce8yTQKQuF84c3YHaFA87ivX7G5RJmVw
5GhNQwG06QNbioc2idquTMjNLaHxLbXyfrpxTjrIgai6NDpJeOl44PNnqwVsLVha
KN7XRxKvxaY/7hmUwXz6TZ5CaKnevvUT7IUhJ2N5jCl2I014NmF7Sfz2RNzbAi/x
aPIBthqbxhl+Iqk03eZOemrHor+BLkjHyORTxb4u1qSgj3K7drSKU+TooxSBz0ic
jhl7whgNykr6P72ghVJNreyZjLgbcbV1kQcEEBuADc9dlZL7qRWbq8Pkdykg/3Xw
fuFAgcWvVBRVdEioNU3l4dJYF2/eqhN/4Oha3bWIiX0Y/keTtpcy1hlZN/6OWljk
46uATLuOdknQF2ddW6/4T08ND/1NQN+mIY5lBxzi+OURAX67M5Aok7BBjrC1zZ6J
4PikCMBSZ60dOpFhFqCqah/4I6XYyrJTgzodG3LwGwt16R3qdUxqEO+tv+JqW2Oo
TUdHAYv0nfl85boeNA3jGVd9xyPMsdQwi/YXFuGMzj/3v4AwjdXJIZAzYJJbaa3W
MLMRkAmZF0DcBlABQws7qD/AjKpCV2vvMkessrFNJZ9TYLzHmK60VoPLZTmUW/2u
SBuSV4i2zOU63elKtr3sHweOrAGQxDr5Y2H/rK5fUwET1gZtfGlbdltfBw8rzvN1
Vftt/5S6X2Y6gpyXO2TqKFYokfaZr1pBjKGJFWwMVYgFKL9q2v9dCnKVI4/pZJKs
GpG2SqIJKtOivybRGpERzfB9P2waHOS2ONgqZ1k8sgLbwH/t8RI93FRN5KMdOA2i
pea2oO6W65LIzr9LKcyT7nBaB6J+YRA4t7rRdiFCzqEY6c/x6PnO7UaCiiyhTbRZ
2Gaeg/NLGPwh3WEJH9JQ9clFG0aRpSonBrTVCDPa/od3leJJaRMud6Xip+e+X14O
e2/kcMT2Ww3hkCGBxFLEROUeI+LDLDw99hdiy4nzuWgEEL9bZztV/GhgKjnibnx1
40ujrEjsBZMk+Opebt+u3IKxiCyWbmk8L7drb8o7s+D5ulNjbjeoDxhiIohJjlMs
TkHijpKekfMqu50k8wX7L4ZpcUh2vLd2jryANcThiG3bSvpTpWGdYqsxQ/Rf6TdH
0Iw8fHItWBILIjxnNwxTKyZpGNTGhSSoB3n/YfFiJaNn1qQxc0nthZ4izqWtErjP
eUj8t/Dm83SW2d5T1tlriSm7F+kegVGQkIQlNjHsgF9asdZoQ0flaWnC9UFpEvLq
tsGPSSVqSiBZ9CZI9vqOAsXK5GfJfW6hOPKkmMrRaVjzIY/Shw71PmD+hTA5W8sf
OTTYV6WJMk7Ht9R/YR3Ucf4tv/wM+lilyY7oYEIEv9gRgxVdQt/JHXrt03jeuH+5
ZJmNpt3Esu1FmD3eaSnHwrwnPVgj5xkX0Bn5h10wg7qex7mBFkkMjQaxU5PjkVx5
r2WP+Io9+nBa9wJf9fCfthGbcSsZFG70+0VR06HoQD46dnB65KGJJ92qCx8XBGHz
0fMLSoo7smliSNWiHYNY6uh0voAG3E/uTYi6cMeDdmQrELs/LgjpgqPzIsqUGrG/
MdyVl2KjvxiJ1QhraX810vStdjcEkYjLq58TLLNF/dqcxGNdc/6Gu5n+Mfpz7HH1
/HWiGxTIVitR0ZYJf/s4b47S1pcuj2gJk+2XcNob0BAVSjFYoHuUjldY6E9L+8b9
+SZTBjRzw3iKkqgYIz71OrV2N/5/bylxKYPOGcv6rth8eX9y+4j9bStSg/arMhbt
PLZrGw81COKx5KJ6yRIrtovzD/dv5Ees7RWyCj+L/1KtUuSZQS9UQme2xIEIuXLF
wFEgti9HyfjNfjQs5ehnT3mFWhqCB1palJk7+HLg8sLBqAgy87TiIGDylmjFLTSo
M9KM2vnU/mo6H9eHvYU/2C8IkRL0Vsk92aaIQUR5wGdPsqO1A9KT3TS3g/5EQ3nD
r6RqBVUjmxKKmpwEiIrSdFCm9LZ90o6V7+pX+UtBLKnkIe0KXeMpjCRk7DYaxeco
hc4UagsWyaiWnei59q1pZDbLjRG7LVyzFO/f6ToTivmhppIZXyQvVZhko1tSs1AO
jKed/BMKSZh64LNQLS+yimIMVD29l2FiE5ZnWwpBoYwRdoMd4mCkdN4xsB5R/qmq
UPYSUyqaDNOJjlND3FD8oor6iT0FwLKRf5eFJdyyo9H7ZZ45oNmQTa/nrKrDBYpH
XJmXl18AkVtKBTtQk9eeq9Ar6njGwwErXAXaUParNB29yNjWjGrQzI2ESc2T0HnZ
TOg2c/1vIQztPB8ZskfuqfwAGgWGVjUUIZbQep7RJz0zY4Zu/npoKLqF43PlomkW
AejSAaXk7Kbu3tvAefEruYewJXqYB4LTs2+Q8mZ7xUUdhdJIKyhC8FglfFG5tovN
S3BGoNYeXQmWjRpAWhjYcyATrW788kA1PF6DdcTvk6M1Ro9eC/dQYG7bY6Rm5kX/
4GsRHxBL3tmuV70h2y6CJ7N/hmkH1as8PbjPsmgCC38NjsAZUl98PJSgbWj5iiQ7
i/LbYjXkTYHt/jTd7PDe7D1c3/e6XgTw3dVab3qubkyItamt7L5izs/cT1rm5nzb
UfpysknoZ7I+iIKHVA8FvuMXCDV1Bk5e5B+0hzgf2LU+Pjo2DznZ+RHnhbTCR1lQ
ZKjeYTsvjxv+/AF2pH4pStfgySxF71oxPW37tc1CYtEvsh0dH/lG4HKMSQZXpXAz
7snZMrlULpR814Lbz1OOGfAV00dbqxIQxMqvN5DGbb288tJaC01PCKy0BhpkF3iV
bhh5u71IqoKS/GdKHrlGGwaPWZHmiW+IWFci4xFbUbgH60WNU8rfO7AhyCgis/xb
/e2D5sRjtnhTqqFQDNAHo30Py5MA9TyGXfmUv3aH0Zyg1gWWjyOByJH92DmKG0VG
PMsbrA7gHDAnsEteFhwef61crJv93U18PzbPvU5MOXXSbhsECI5I5ellCf6HTzoj
w0vpQfgwFNPfUlQ/OBiOEE+31eibRUgDm9h9gocAZi22fUjUzGLJjSmldaDTsGsw
+fY3bZkdKg4d/rC8pcldz4EfzxYWdNVvczu4Ov2Cog1WVBpWtNiMT5RXKcfrwVy8
nJY14NnM37uFz3VDRcC2Uix+oUCRoF1dw/u9D4ZC9GXL7v4gjtEHCD2/gtK3u7b0
JnBftPqdtC+jifpbTM+YjbqnAFBkOLClwWtqowMN04+w9M8LvArPyCLks3L+RgIS
lrenzean2bMhBKmOb/jzZgSfS8Hys71cds6VDMefzaRm2WFvwRmdSEeLPLL+uRKa
fQs2GdRGytJVJXaFdgKjkJjU5LAREHmEi/TaH1HFBR8xZJi7ed+iREmonm7A+A1N
KH0bVRntHTIY0qNzlZxqBA7QA+rfdrchInnJ9K0/3F67DUiBjv/ID/vHMva9NvIe
GG4tEP2vLRPVeUqcVkoNxcBoHcDDzVMAEX8iEfnfMg8y465t0iOSGu3S5qjA//79
rzV6QQtlktRIUxSeymw4vL0bfOBQcgUS69ll5+5/TZ4qjnpJeCYBf8csj8e08Tke
xGj7mBqYeXGSG115dDH1l6HTcdvxRVPrlNN19Uf87Tz6s514UPUL8qjyh7ChDz5E
UiXbj0Rb3haXGtiNGsd5nxw5DXIsuJZYUu6akwefTKNNNodcm7CQQDTiorAtASKT
cwxNr+gGriGoveF664cjFqJHr9eVFUpKFRD7xCEgcOFgAUXF4dQ5ZBvZM1H2yEkm
pWOgGd8sukqtrltnU7noalkm8sePtnAFVWcS8ov/n3yXgocIIjV1eYhUqJs/HpFc
xbAEegAlAP8g9bvqfoN4n6p36EKVplJUpJ6ErXBhzvWOAtWVziU7nTy8efKLT9Mn
XPa38SPTVjWlv4T5aS70nie2q4mxpmrGekcD+95K4eK3zcB5rMICKRD07LNORhtX
rSE+tBwm2DgUDWC4/18Dp2ZSNNDoRUMol08wquirwIfkw5MmVuJhtLinRrw58JkO
VV/OwV+/Bs2hZINN9/BS2slPjmgaFM4t5pr7EqDV2ipUwhIG22vyBsnInlfEGVHX
DVjXY7kDtT8KIWRx/fs5avhBBUzk0pf/GbDTCCOxZDjlbNleVbw0GsLCK0tmdJqh
YHVW/RuNea3bxhgzetdVT6EylccU8vLBLS+ghHvSLRk70CMsNOAjX2JMG0uoAJtd
Ipb+MVsOUH0mdj191R7/oaxKDXYWk5kL77f4J5HSd6f+amibnYnKiNVvpQapQPPd
y+OA09N/xLIuBBrJFifZLOBnfZKx6zoFzyA55KzIpfZ+/MtxKjhDgNAJjTwUMk/k
V7XYe4CRrBwugzAlUVj8+6LeZI/pYoyrjvML+Ibzvj11yZwjPdh2qXul5PiGnoI+
rZlQ4zftOnT7kmuOS7tFulErbK0/gIFZjIvNkr/jcReL9HAq/XSOnJjxUhsIW7Ah
nNuQuEvMysdT+0qOkB1GWCAQU+8yyupmOBTA4nIr83UEYeTVCAfoBElavoqO2ke8
7f0GNiHK6D67d+jQx0OxbsylrgfF3fvJlKPnMdy+pFtivhx4/ej0OL0KZjZRc7Lz
y5j4zjBXyHTPOyZH4EFvhrEJ1WSIrxtfQc43PmNfZL3iaI++9mWAbenb0j0FsTcC
jteG+ots4HSf3rxhw0EOTdV6kJCAhB85Mxah57CMYo7nmdiSlHeiPaD8rWr3Xvqq
O7S60N0i2r+yfyGH/kgKm1ROfQNleDMOmxgW087RbKXkxyddgPMYcMbrLdfEvhMb
GzWdEB3P6hWfhmbMd7f24JFvrSWGhHc4qR333R7QAHJTzwUUWNAi3IMvQPwUTJma
hmlK5dGbdURaPI/Qn9W3K1eTEzh5iUdK+sn+9TUbvW+jIdECTqm4xVmj7ACwIGmc
s6wWJpUbo23cP0zja0Scak9ny3aJ6Yfnak/L4sPtxSD5L5lP+JxMALf/VshQSCNA
zXG69Ng8b/SWxGV3nVV3Ox+Y5nchxMsgin2DAd4R8NdnEPvogk4H4NzZjmwe24Qx
xOXmLxryRDvLLFeIl5Nv8qXPaphxYxhGhlagxzvIyNnoV8LYy249U+CazeQkxdKV
iss0cyrewGEtJfd9yGq74ZfYM534Aw+Drt6zAzFVCWhzJrAOwrAYD8uaqGP1EmOS
Y8yJoUFj/dSofGZfx8itzspLWlYEVGawvj3a7GFrRSgYWd5fndX5R3ZSgaa4Cg87
BRJLzFPOam+hW6YYk2b+Py4t00p6aWZDPs07VrDC+/yF/+hD5yrWWjVD/PDFDYNG
B4aMyWzzaL9s6adCdl4bNTG3iJbIhmB9ta73J9/8psCgDa3AQjVV7N+x3ZiQAm8q
+O6M1g//50DVJgHj+5OFu2iE0VCGxuGsQiQU3g7IeexAAzozYxJuyh0U+Vk3eC34
9aOKKNfigAWZmbAre7lqEdwr+J2F+2WnrtS3ZxdbdXCO79C04MBWIk4Y95lovedd
IgdnAs/X7GdYjAwDoz9kOQWz6JbzMeC9TSOF+PgIGgIxECBDbyX3rSElhKzxqVDu
dmplApwRQxQ3ud2ZFsgCBrxPVTVkqDvID6D9PTcdROTyWC3jB59ztdR2tVVJA2w9
rcu0CfGGn97jdd6JL4nUTVwQVjGnOT6cr7bqMN8ouBIM5SqDjOULanUaZJm0aHmk
zx+OX7gLkUEgMU9ao24a3cq9aHWqlhsrnR7jbqeKHxZUk/NiD9j5GQq5epfFaVDq
foZIXlf+UV/a5YFxf56gV6gaFnOIBwJ8/2xAyEfINq1++5hf1lgZqJq/UJMEr4UE
+gcq1ZVoVoH7ghFhmZhFtg1Rk51pHT+XW+zGLWxHqTVZjuEohu9UC2/iHLmBg8mF
RnEfF6hrrlhaJePCUmo/HToE2fpE2zXmrKJL6XOY/YoNdMRs2tj/re5xuhq76ERF
+Y6NU0xkDGmezvxQXa1/IccRo6o45KNpsXvY5XPf08ENeFY0F3YNvcaHFVlvp+eo
iWbyUed9EMF5Wicv3pobXakXIp1UnUqyPx51DjbTW6jFyxLxJnQZpaihqVitzSJ7
dyCOcqrcIBsrO27OUUesWqcCGnygkhkH1zXsbm0iW9+EUsJCojhwZuz4qHceOTMB
J7/V5jD9PL/PY7vYS8OIImBBRRL+EwBP1SQMUcGcK1tg92vmntq8Gwe+aFWBsnc8
IKnUOliJVefLMX/fvqVkcW0+N1X7bR1k23Vnc6rKxjtHGAk5ADlmRwmfLwLcXnLh
3LYd5JRqQGJ/L/07PiBhFo/zh4y/kQ+lTGOlNCeIliBQlxZI1iGVXOn8+KZWcJ/v
zWcXnjakyNsFFEPYCPk88OLVow4Uesc/2iaDPU/xxu85UhxoaFn2ZVzT240gFIRF
kKwsYj5fcHDwTtnYlSLQJ0TUIXR2J2/tbQPKtTMLVe5yuinmRUbwy0dDGD7i0/79
aHPASO29mLw+18prxTG6BXSUSPOueW4Tuy7k4BLY0MsVOSyNTKJr6DqqlgoFnrL+
4vFjBBilNWHbxCxBJ61oA9U0ATb8ggUeYmj6Ll0CtBxWPHeoWaRsm1t266sb2L4t
J13Y15T9SEqu4SfrdWEzeJQrjZCLZ2OrPq8lr7hVMehM7/NJO+UTFSskURvd73yo
zSpCCa7njOCP+O666miFCGG3HfZ52RdaH6R6gpO6EFj/H7GcMB152ZAVMBLuN7ns
EKE3+v/i+o+zh5gzyjbu3TU57zO9qB+Sno4aPby4e/E+KnbMGIHCofrNx1tm3xY0
bP+EwRRMrdOk57p9ZbtKSJOle++LlHWG2WG8jvo8WhpfQpQiX05mawvBRVvFNC7j
PrE9Qlqq4H0ruqdzmktCucxnoXy4Zxbyz1wHDofeCZkX7iO4YG/6Y3zf0oHQIzbF
uOoLXuUt7bI4FQQ67M3IM0LkGN5y13+uG41GTj8Fk2ajAohGXlcp4MZopXLcM9FA
1zQ84lsqmuYvsBqlOc6DIWt55IaB/nZoVkxxUR8XyShBM55FzDB8tjtuDwTd1utf
YY5nsaNFNtEIHQ67vDE5MeKDS9UE20TVm5TURjaNR5RBvBklcezBJUrJuSLUz3zP
KJ1vcuA4yBCu069AWqglawMPKe6qudsMqgiudWW/h1YeCxwTDbjhgAJcJ5EFIiDB
qAbtwf0RhhqI1x7zXVPSk9bkZiJUWFlYaaWlM6sZuxvyhfTUzpbn/bggdbj9IkAA
u4o43XF5TJ4CIZ8t36MQwB8L4X0MXWKfJbKoMwQPgmM4l5lkmYTCoB0DvjvKruAc
XIMgDJuPfSUS0JuDfTVrUGpQ5P0tr5eBMH7S4i+IsZTzOlLhntH/nrwdsCTfy1G1
pllDZj9OjETWuyUM1wKqohxwxuSbJpxyz8FsF9bQ/+4OXYIs33dq5XvX+IeEtLXY
wwkaMwHnsseTYkRmsQWl1eKEKhVicloiuhF8/KJYLbBgv+FCfETY11wt5ZbViSih
+PK9SE7apV5QfMuHLQ3gs1plTCB6po7GnolhJBHJeYdbtQ0CenuI2cw9iXDGZ+cs
B2BrlSJRS1ux0IuDv1eXkzw6B34y5PMptpFi5ZJnKLlKWU93bzoHbUxWDPKfna58
onuAHjDICVOlulwU0rmN8M5dZ4/5UB+wY28/gb6iLXTDVsLqPjcYdgFqG19z7W5c
IedOC3Zn++HZNXTVb3iJ2eR5dMaqPRkR7LDtWtHyxaxPCW+CMJkugvpfVZMKuxpM
f3ol9H5YG57ngIidfad5Q3x3svu2N6UzmFiuoYa0ZAnScpcr3sPmHgEY7Q6+jfuD
yfqRULZ2tWnYXPZP+k4njG156AKQV+6DVCb1JejF1iymQSz/rmbgZvY60KiLVTcq
CeGJTrifm+eJfjkYB42G444SaoDwBbi3O0Azn8UwkpBSQYAWgOUcJmNlsB4tG1ye
lH6TJy3RDucvPC4VYQpxRjydbg8gKu+rD1lDYrap5NvE9YPcM4ITFrL05W7NOtvj
T/k5Ce4GOf9qbhC2MjXSgSF92pDjsSC/nwNfRlSAsQxPH6tTu6YqKdwFQvIwg+of
g2aK/cyXOT8DPYPgw5xOa4d151aLQyrCxD5qSQHm9eiH5OGPYhHj1vwRdlDdx25Y
gG7zqxp4rBVyvKx1DvH97mQkovneA3duAL1UBGv1k5NvfaB1jWT/KrqK6hwjOkEQ
AtJY6YoNmmt6iiCTVeifWA4chEbmmULA9+2hu6im4uDsowSltNkwjnwQ0El7stUY
W50YLZTqL4YTTIydmciARkVnlY8hhHWC58E2GDLLbIJIta5UERawPlajiEo/5LnT
5GZHB8VLYdr0/XA/Sc8CE/v8+LP+zZKjz+ByUEu1D5sJTy115R2/Z0fFINiLYVtj
xOYu8d+iHeMc8ibk+T8L+qeDI6S3xOQnL1eRzF9xm7q7bl6ujToMxN/MGU0Xcdwh
5MtGVekyPouzqn7Ao+88ukUGQ2PHq0NQBDPpOpdBRJgDJb5Ykvi9VopzQ5J0bcwU
XE9ee84/VjSb1tyzkUKf1qglQUxcq99B30pBsV8IRyJlZFwqPDTxHhqQt5n3zMUf
pH8kmgtE+38iSHKbCdRaskS6L297XcvRlHBRSmNJCrM9iq75Vc/MZZYF2uDhuaQ4
P6U9kG6fYofycv/iAnC/QdMZQDmxYZ8rGlvT6fmoTeiYBfngIgcmRNTjX1f+KcvB
0xLZktmtSM35Ajd4Dbh0gvF6sRwfDjsUshgHTczp+anwuSkKbSndUI6SeS36J1vD
gCVk2Ixwa21yUHdpw3jiHnJlKA3ImFE1XtKAHGVc+0qZ+IwcraNzyCik6ZJWB9Qs
jpmH5Os5K7fspntnC56wYpWLWswKIORXBwpwR3pyKieGSEpFhghFlTELINtP2fAB
I7VYC/A03PWDIvLmkEzhat1nqQjtypak0z3ncpOoKoHHCFQ64iKf9bAkabIm/y/f
tYA/TI3zshG1nPQ1I7g+zOvl3ba1yGIrQ2oN7yETs/WF4QtGw+vtmuprM9ldXq5D
OHPY1Uwg3urvrr/bP8pdXAqf3HJR4M4gl6ZzqNpt/99CuQGqJlTGCGdY3LWfSovy
GdBZp3b2/umcsP8QRTAwjpXd2nsFh3c3d9rMnMhn5rg/cEbSvATB+q9XTCcJ6by6
9bNFpDF2jSqpbzHgpbBI1/gQcS403O2svuYSsAE/TSKAE08ktIq3DqYDZAVeYDpb
T0m1aX6WSnGrcIQrf+5sYTnb320MWroazOkTHF9m522N7x/mgvFGUAHAR82S4km9
TAVYnTiudVQrZSsW2suckSofT9gUFWkVZbv/AYZQi1NUmD1YYXuw1+pGJXdtR2eR
jDlBkA9+RjkSrbTKRQ1WBVHDJyZlcWKx+jyO+NkqEY/jma4BPuHqjdbv5JjA0ry2
abNcNZ48euMI/d7Fvu2s97X6Z6l1DeL0TpE8ps3E0TG6u83lGV8IOWD06wUMAT5Q
Hombts254WClWQ8WFui3I2Ygkj9RktsU6KKasoRdK7nL27sNgHGneSulUvi+iKsY
bFXQYehMoRE1u+mwxGYxqt5WAlOoyUTK6KJNWjqGxqPdK+cB5RJ08UpKESzv8kMX
GI8N/4TrjNbWAlTC1K97X9KlmgF4sN0YyMtzPB8lbVvyHjr4BNN6/0bFadLbSRW5
3Nfk7ZzLIFG5lMF+LkWm5e6sM0wF1uu2yHLjGdiDX3RWGbQuvBCFvVveX6s+3DmY
Cw+JySvWTK7gXe4rVYOS+76OWV05M4Khw27ostQFZvQYT53K0Qa5FOVuOQgw3BOT
YPUKwL8xf4b7hPRmQdeLLpiVs3IqzgfdeEmklNeU377JiX9RRmTi41BSz2buSGhE
JQ64U02r7LPkgDpnaXQhESS8ME12ikmBtkmrJnm8qZ+c3V8vtE1lkjP+7sjaZcb9
HM0CIfTGyMUzW6wsWH56m6qUcpu0EpEUYhqmo070Ntao4XAkwN8C4XHowaGaXiqb
83buHeWFrOPrO1WNCrU7cH8F2bPqXyGP+9Pp2uLp+sH8eFJJgfD+siGWA/GBb+pl
mokbsk7x/DymBTdfrxc8liFirQhfd2ycMQTDsn0F03JoXDNmI0nvvw55tXwT3L3k
DSq84cVeUNy7hwKOvEsQWrsnPWR+XYIAkoJSVfgPxA7HxiytGhCXLTA+BexYVmoj
HBkfIvI0ubJltreD5wGvzNdKxkMH/KpWpNjKEBoymTnHEJLSsv3zgrgX7YrjbXDJ
Q0djJJihdJne9UECvLedtGc+/ifwPAZUcVpv7G0hkFG7mjvbnT+NVlb+DIakdc73
BBMHyTiq31oX9fVrU9DzIQ6LyFLlMJTuIYJjAe8qPqey3utyMjJndbPJNfb6gLTn
s4Js6TZJxVBrc9CGOBp/ngP8PWdE2d7tWZYqFr7vxfP50VgpPwm8Jpe1SVqxROAk
5rAquk2RB1q7sZKlItZqHNfAwtBidSecue8eRtvzrHj8v7tNTCTEK4HFBs6afaQ0
Ng+Gkr0SNnsygKxByuhNLE4Z5DvEQxaiD911mNzDYbnkQWitffmYBdi4RPrri3xY
sE8HHJMDmeCNX5qOCGwaQiU+r7M8sfYuOYiXa8LN+lRWAPOuk2eChUFfGuaiakky
qGs1LWOf1w2t6sWSuvMTe1mqtwr0wE87g9DXC70Igh3qIUtAsEr9meRms1X7NXhz
Ex3ilBijMzw2U0ReT7sV4izjyf5b4Vf8dSS6qhMFc16/+wRDSkVp+06BkY1K10PS
p5nO6+PgThXU1oUpfd4ImxR+zsL8BP0myev/p6YiuuS49JCJr9KoRerkJFTHEjiS
xBAwvrEGHZyE00AZeuAn3iNWSwA6kkUtgebaQQj5Q0gMRBTVOC7xrKPfQUeIMwZt
WMqQJ04sk6kO0Ohlh0H5/L1XnFzpTnN/Qrfjl4IFjy+T1qgubZNnruts8Jwfhy9q
2oGPbfIVtUgBiZ4KdWqJaRI/xXd5jjlaWbrWtgyd/N62L8otQ5go+wbc359yn9V4
IGt3FfCU3cTIdl93/T7fuQySi+6SWOHTH9+u4vpuAjhg3za41/cBDxuBeAiTD4iL
mvMidYHS5XNZApRY4qUBQFyVjFS5+cJtZSqWSS8fxkK8BYASokDxeBKCAmvMbH5Y
6udFJr9F+69a5os1aBPWYrXbi1n7f3vEo04Md84dpNhIkD70QhN872KEgcsToOrA
MbTLCagiMpGiu/9sTttySCbz6gJ9hzoFd8JX61KnHtViiwH46wGeW0yE1FTXPmxj
lshsdCDZrVSkrL8RXMZqpZCBsxGtaWpOV1xEZ0ugdmZf8zXSaF/VVyQiTDMRDeLF
sfmEhhP38mVgvh+njn37hd/vS+V8DSbcs6DCimXG08Ws/7NZC1wSHeQWFGf7V3rA
IyVTa6m4JPT7BUOKMO1FnhLZqzEPYY/X08wXI/H2IrC9QDrSvkn0VoyWPCKV6K9h
jKFIBGe9XWymNhGRhmXKtzMZY+YRSb+Jm2JojFcIxLVKiFd9XBlvnzHBRcZF9uas
I0ZzgWA91lQVab5S4IVL+MuQ53XOEq0PkihJtKmjyYjofbKx8fjZG54WTRBpC6NI
RJm4k2naAU2cNAMWU2owweOCN7za0pV5ikZheBtxEt4bDj7Qf0btEMlFPXYD2lY4
ipocc3WwxzJDPkMACNGdqpfyJd0/BTJk1FVsdTG7mYeJQddpiv8GDYAJSmPK92kG
ZofJSYqq/ypHxVYeSGx97ILGrXBL5ce918lfJbDNAsvk3YkcMZwX8B5Und0MdIkH
jOvNGju9pkpoYIjofAkUvrj43g54u/mhvMBIi7UqMyvP+HrK5zaGEl1VzwPkW6/G
prZw+JDHraEQ2ww514XPithTvII3kl4E8Nzy87o5FfMqZTA2pAWFP3q79itkIAv6
NbHwPzj+KR5nf2Bib2wRRj2Yyj4bNVWvtGKfUCJGGwpQPoW/Yqv+nTC5TKPGImZE
xaMQCgrFla/IGN5DQmtEO4qO0j/oC5c3giqyOMn2jjdhEw/uTYQ7kMxtwfr0ZzUb
4AG3bDC68SFialqs5Ti+2kzxV16CuUN39saSVDenrFaKGrEjs/LlOEKXT4JeEPR5
KR/1laJk7Y2vlvKx+qNYu/soUk4kzVpRn/HN34X8AYXH3fqa6kw2JNsbCgo0JUPq
UVAXE/XvDzbAUnfzx4GGnZWzfYXsgv8gzZuUlZzeaoZ2GNEp+zBpnfadHW0dqCHA
cXlyZc4Lz/cWWi4IGwAtJW2p2LLIvUL8xHgOQrHZ3+KFwscWe4af43ED9gRJnCz9
G0aJ+SQBhpECBd9NXfy56eCmiWZAilM80AJrXmMVUYRseKHGy29zHpzlsreApu9G
/PmNEOA9QCEgnJ4B/Zgh6QLfRqFUXCRSEIkXV49da0BqsO6xLZ56deCzbdniKj7f
ZwfTIj8vU1WQP/mXwHFLj3XU51UtmwNT3P32rzFQod84eX1/VOKfO23mHvyEjaws
XX6xOF9Vq3iEfeekS/Zf04UKmfivdCccBvR5TG6VqNQNzoIm5JuKwGfgdupn1KmJ
0/BwLs8acZj2Ua/jcm3XERl3wtYA9wTD+5YTUy1q5WMF/KV3uFnbElneEvffygO0
hGjX5ejuxcVPT4AXd4qI/S4sSNyeY/FduHl05paysQvQiSib2fTvJc1p21q703KH
dY+mrfwzibSGuCZQ1OCp0y3HrJ+gQjMdSM+QF+n3hivog7N3p/Rb2hPMNXlUprq/
vI7tz5r/tNRQdSQA2BEJDwJyR716UGkWoPrnIHrLYOVxkSCUyZoJIygz1EEDkImt
Kk7yAIs5FnljpKhCX+So7Lnq1mOTRXhbMNaNuy/15hDN9+gEaS+a/yFzxV54g2zV
f68k34++ouDu4UZaxPfPCMxymO9hSHQnsCHeoM9veGSiT1P0fEGjOOf3YNp6Jxfu
tf/XY9HceMeKAXO8Pco8IrEvvJXMNBc6gjYlv0OcOd4P8YqVsZp9Sr6BaHSXDJjM
dsTQpu1FVJGWmx5/aAK/aQfsvnrghrCOX0feqoGvgh+qEXMTWsoReOEozj7qtsUo
802tYFK6Y1LUCnICTHL/sZkB4IyHCZSNG0ztM27Jq2Bc1ls+HSMC8MWF/fBEr3Hp
iiVUE4XLzVGQDxO2jZdVM2J8/VPOHDOdlgdtkcb4L0OW2KmCd3xPfLxiDJ2aACqt
JoqI4v/UQ2AGbp776pUnmVjAC8cx2ML7wm4BCyfgc+NME083Kplf/4lVtu66U90d
T4rTk+i/uDU897e3yBfVyaxywLTA913HEo6qeJGpFoK6Vv5hUd9n4dtvNK688FU3
CNs4YSnWLbw/4guCwvUw2FfAun55tPtZ0UZ2EJEGggZiRjYPthvvpmgZXEkLsg0v
iqe4e1Oh/gNCah/48s6kDRTnaXoHf2fgggU0kXMEWSwDuR/sKmT+F/acrrDWFdaN
jW4MPkUkj3eLPb0Qey46IJlwMnz/uUk7xL+1GGrpe73mlAKppVaHnWzFQJUxMJPv
a4pn8GMCuoU8SfdP1Ed04DQOZPlx950m/qPapwQjCQowfu6teFwIs47eIteq9kTo
0qnuehAiKSkmbiFfRpYGNNoOXwM1xmhyVDOJhr+2R+vvqCqnAJh635VK36tzSYtj
g032j9nAYBJPWslzsLOgnZgPmA/Q69ndz3x70pJU/i5bmvoI+L/RbvCgk+LperBN
rJpPc4XPrB5slfiq2W9XD3J2SYfZHHSgpzq/F5PJsdKqgMj+odWyWPT2IQwpUt1m
tm8DyENIzyfoA7C5Ih79rvGtfRIXmr8+neE8bvM0aylslAol/075OaTdzRHH1Hhs
HtbkGaSaczhFltVCIkKIOZBarxOeZq2BaUbydNnkK8N2JZJe2VsL7dFNVoxCwAll
fpQYZGGWznuP/CDq+H/tP2P3CYjLfwcwsQBbbCBtaoVcK6B1YHeg3ppwTZuPOSiW
YzQcXQ7rdbC3d4Wr85PCIS5p1dszdluSP3MkMbWJpjgMdaEBrTeRLv/jQ9WR4dHr
/pGKgz1X67G9xnH48vFeqR8lY/qlWBoHCRv1sfxuMPVNU1Zpo9pVFALrDqS39paZ
Y4V02c1QRKlhlgcipLWHA7FdeigW8uYu5ShG92uh2EHsOZQTTJvtkYyL5mEhuvcx
be401nKXOWVdBCVngEXk7C6zQ9o2QEELCbKncQT1xhxXpdMdtcY5vrPHKnQSHufJ
zitDV6rbHvelKvQ33qrYXOTgL6mPM+A6lq45/8dBw/rte6DmIJxpQwYakzGQHMma
VgpU1gFPxCsqcw4GAjguzgiX3kfybxfUhpJBIlredswZaar2Ozm5+1VNUiEU4Dxy
pY99UjtMBeuAlr4UvoxW92X7osubOZ+7jxAg6daqMhc4qyKJorMmyMOu5G23ppkP
aEmzg1WCjpCANDqF6bz7PpDahNCLsScDuA5or8YdWTS7PRCiIRuHEKl40RC4aS1I
YpV6InYOqg+N36D5RQIofDV/h79xZjy8XQNymCZiBVNtJp2aHGvd9vXPRVl996sy
UM0pnD19lCD27Tt4HRD6r+TyADYVTUUkTVu2V3JnwDymSv2ZS7WJsIJ778yyxbOM
l465ny2xTCc6m8PJKfrcHV8BY8iJk6hy89gSXdYI1xAvPVRDxV6Xg6gSllqVyQ+y
3RLkiFQ+W3mKiq0Vo+gUtCxajFc4rRXIgnAnqT+p1LK9nM/34V61kMhbcIUmbFlW
JYOAIL9IxYVb4u39VW1MfhMwfazAY1hp9Aqnimkv7gN37LIf8MzZZDlMuDs0b8Ak
T87GIwf/MtuoEsv/NgTMu+vhZYwzZxHuwRlVJ3E+IGzAVEbyeOW9SZomA5XqIrEU
c1R9hlnMw7NbhofTj1/e9KVVqcFJJgA7ubbcpCCdFyqj28ScSBsaeR2vsj93BiC6
cOWexiG0Y1CyBKwZj2hut3AnpuSacRuCWecn6NHChMTXh5jtScDW/JvP3jenQyu/
Sd9PeI/RgDbwmTws56Rz7jDkRo+soQAWwoslzOto0FWK/hgyxiPiUzNkoc3sNpjE
Pg4Awx6EuNk+722NoYGzdnVP8+Bs1b/EFa3740ZryG0H2jAsDGQDgerTqs61Lh82
ZxWygNbZkaBHJ6+npLoAqry3PejE/NGGwKpNnlsmWmHZWg7TGGRafgh6dqUTlMCm
pe+eGDp4yjmqEV9NNqwz3yQPfocCPnBRnL+/FwHm881hg54pAG5T/ldsfY50x2rd
4AQyzsy0kUwFNj6nwrUYYaUXQ0hcVQmXrzzp62oV9WNx+XoNXGlYoyD1dkZY02i1
C05ohptJqaJiWrzPietJN2g5/5di6UgQ0erC2upZ8aqBB1dZ/QJe1KfM4iAk20sA
bwEFbhX+tBd3UHmJ+wDZFY56Eu+tnzoDF+h7wpLv4sGfyU2CSbQvKFpAq0EfjnWv
wjpEH7izVYkDUlPiRmlfb9OA4ytu0h/UOYJj/pTIz65uMLSvmT4yqW6Y0beWzTFr
OPBZh8hsL9QIuozguJfJkd1NcgI4zDGRHBLaRu+CjViA8uWinQ3IqJmh25r13O1K
rLY6QRS3NFAAbUC+w0PDrYDMT9vlU5eYroak3ANJV8DmkPAcAPCMkooKTOai+HCM
Q5ESrmciYDgFeLg2yjjWnrXVlz9yjCPXW2SNK13zxFNbw8ZqcSGutbRzFNUkmGLe
5w97KjXLRj5IcPnna2TlJChshOOGFc7qotOTnrS05OToPt5J6Q5j0IQ8hUjKUvaP
TUlkgLNs2d2mxEQ9c3NCQOZoqGPJjF5tZOrGN5y7abcVZ5IG3H5A6XtjfAU53/Ag
rerzR6tmPyCovOj6pPiHfjvbNWos24uXIFX2sKMNZHz3CK6hyIl3tDpyN5/gSkgj
asekGm48RPKFXldVi8ai0shN4cedshbi/7/xBI1xcm8a9zRYa3OWVlu2fLvaih0u
5Q+n2ItzybCC33uuTbgt4vt6ZzOu9+v79vbZBSuxIccOOHRkgfcIXhl8BuuOKZYw
Sj4NqzBJHP5dqxLOn1l9fbycxyIq7xKDlsPwH55jBXNE+ibnLvU4MMgY9HExXLd8
hQDNihepz6xbfLw9XHE5m50icM18Y7VH9B//CBr2YcyrKxuLCPteI/lcx0hImdNE
ybZ1VobUPBtY2USfZ944jpvcs0Nv9tEVxqeV0ljuv+3+SgR7WcJUpmZchfUtmCRb
tHFa3vLUr+1BIdUo6rWkYcob1Pznc3jtFQI7l1H30wAhbiXe4iT+AIQaBT1ptr8R
vH7NZQgHnRUDy03dU+HmTFNCURP5M5Lq0RfNxbLyIK7WckFKMh4YhCHC0KvmOnCU
AvaOnWI7RMnZZCztoezbye8Xa5MDsQxSM8cGMkYRXXblpOpPRLMEQKf9jibo1Ope
tyaG3wBm7bRLEbgAU8/rPI876J8Br7VTB+o+uMPo5YGt2voB9C7B/9idRLYHW6VK
9L0dIDueXXxnUmfR2P94q0Io+DqzC9Sr7t+RWQY5oNr0Ju/McMErjJCUoYLmKve6
jbLvPOI0VaSQs496bWtqdWIzkdG5Pahbkn/KMUPDwm9M/8rP7ZEqebbaPlq9R0rZ
ld83pNDwIPmxGyRhTLF9DcD1LKQYvbWV1Bq46Ze2iS8poTpW44+yXApRPjddrlMV
FHWep5Gb28c0oqXyJfNZxLJJDlpMKBKzDlSY0esKYWKI1spmtUXlFvtDd2E/AJ8T
et+alxR/XEYTNerg/cv9GAKb7W83UjD38ocLp2YN88fjCJttEKFbhGvnaGHbfX7u
kVmto4yxGIQMP0uvfNQmmne/AdGNGyHSt5O2Lv2Kcznd/47o4AXzE0Ga4DvQCV4L
jcu1k7R7rFO4D6qbcSV1lou6hb1KOtnjtXc0lVsgDOg2X9VxKUL5MqIdOo82fcyy
/ew6HFXca6NLzjDsyPb0y4E7cbqDMZF/AIy+Hlrulu97CnLrrjdIhfRvkpHbiD4W
e1PWweTu13xqhAtokcH1XHWyYLY+NEbgk25n9XH8F7xkwi8I1rvd5w65lISIFEcY
Dc6vXwtIWg1t3aVaCBg0579qxz15Qc8WaeE19jJPlcPyfAiMgRcWlEGK/ElBNyGa
wMK137tK8bb7MLUFF54Tyl1Fgn3UVIyz9x605DitQIlJCHszfO+Bp1hJ0t/jraEk
P1V0rp9TS5SAQvEKFYVRXy5zoWs+Dxp8ZapdHvXPpxmAH+cHEcWBfga8a/Mgwg0a
9jqHlVrvykD7kONMpGxovpq2s8Nz2+zjqYpPev5RPQyD7JZ06XYtUDkasI0MW6JJ
6BFxGX/ZOy9upfoD6jA7ijnkQTRqWhPP7hF03uDCy+TcbCLFBlQ14dHYFA+eziEM
TzgVXEFmr0EXs8XN4oUlKaqA0DcKawkSb7sgvXXbiIGxh0rK0hm3uyN0ijCYeBB2
a9JtbEnglLh97C7xAT2XYRReGBs/UaUHoz+Wg+erAI+AsY6P4tCyQTl8fBfpYBsT
IhLAHe3YmF8QKYBU1hbhqHb3O+iln3K+0OENrHT8wUpW2KZRnZey5ECAPrDcMSfH
7ChY7tpH6gArE82Xp2JyOLr1UpwblHM8fV/jfO6CNW2kD1OwoaPwzXS92j6NowFc
WjHqu4elmxObXzkjL3WOkf5GYr1Ebxy5vhaSxk91IRbhdT/pfZ/hGi5p4S9maIOa
8iXkZ8DSVLY0f/A18xYuXBX86o6aMouSPn2WFB328vqou5bOziUWY+ntapxdMKl6
gxJATR/pr6lxXGUwKKrsTaRBni1TOFMXmnUm5CIynwdNHgRZ5gk3P7JvBFc3oXiM
HpjS6cvmW4yD3pGRJw7RfXaFDbocJpB1LGoh8d6rIwSYtZot3gInA1WjlN/Pf5Dx
Kq/6iHiSdCBwhNV+pZ+m6AuIBee/kA2xY84pDseCe8EwFqdoCKDDY0pPEVKLcTII
Il2f8z72Ou4QM7CbgAwcdH/yltZoQ6lYg+BuPzpMQ/JHhW4hEPl8qVW4XXdiY4Zq
J3JSHaj7XJs/rXYittdHfFFTfJnqMYozD6p9z7V0POY8WowPKVL2iasALA+fPIsu
gmy96h+Rt/dsfiix/DDauYuCv0txVsDeEmV+nVVh+3hA/KoB7O9pyTPN2nRDQW7Y
/jxyb2bWWQcoaZaQhSCSNpkfDYnkR+FOaShmtjIcgD/kINvGzfrBAoHfxcRCVnfX
BgVT3smq1tx3kXdtBDxMD/ZcQrzRO+nIolTGMR9q0z4QC0NrVMUC0u9RkJdkq6I5
OOzm0znfFHgCA+DO7ne0GTOvyfK/kRdltpPBQYMzBXcck3DtYj1vO6Lsx7iBngSc
db/+y2tSHZrna9E/VeUNi/2B3+5BhWmo5Dyko/wzSNeK10rcIv4rIfaY4n1CMN3s
yMCXgyZV6JJDLx7LAfcu4rc+z89ltxuX0gU8QM2DlcL5qwzrDp7PUjXdAhXO6+eL
cZptCUBv0WlcgH8apmXdk+ytwMcxcGJ5nZ1c7e5TjdnmleYfk2VoFgEY+DCCFBpn
f6a+JNL/E7orLRGsBjfjNJRg0koqukcA9F7YhTvo1RuieVoK1U17V7lSv3VT2L2o
KzP6d17BbUpgZq0PkxR5almHefuP9kGs58y6ehqPGqkorMiJCAS2/qgILSqic27k
BDJxHhxh0RST1zyD/iNzDKGcN1oSuNh9xymRd8MIrQPbGIU3Vr/62Z59xRw4nbMq
bH3q3HJ41ecfu59hL6i006bVNaH6whE2Psysekn22VSaQR0lT0jBc6tSrFnTASAG
8m6yLQXWduLuL7tMzKDTFo529BhK5vPHEfZGYMsh3XzscF/X+woTOHFsDZfpe5YD
i4GQThjVjEZQRvOIN4ySDlVCNlRsLYPhoZKas+VJB4jnqBEqCNHA/RVLsYGFLnZb
sTDb9RYYzWp1+1vw1xDRKJoE0LWvHuwrmrBGl0sewqTlnkpz9yMOjh4M9VMhXFbH
LsBly9f0K+Ka5wY8q3H4UbPHcNQQGhsFttlkQAA/s9ZcfpU5W1pvb+kde97BSJCc
hQkwZheLw4UAChQVyHa6pnQLI5VlEyCGTvJeKjKqqCANjA3fHSUoqxKgTlEB2gtx
qtiPZ52wRLMv8cQ4XlilWbBJGfaB5AhMjCacOTmAaxbTYI98PgFisnNwoNWnATmj
yEQWvJ2HgNLVuhWRkisjmdpPtTYWcx5lwxdSWKL6OskN8w616KgUMYBPAEHeqlE3
HSdk10dLXg5CdgNI6xfJP9OFLnZACez9cqzPUfUgRzhD4CEjaKCTDPUZdqcpM5/w
TR21XXqgkFZtdF08RDND3gprwo6/LqTpLWTFVmJ34soqFFIwJY+dx7R4VCvFDxNE
k1tYXAzHY0PBiMxUO95rYdMJtqBlgTOLnbkPk1boj7JKBrSLekkvSlTaMB9Jcfdu
X5A9GhpDAuAGVbTkr6as23A2BdOLlc5iDVE4gISfAI7jrBq++nyXLqSpgxuIdxwR
Zqfq/hpAPJtcHEM7xEUq8sIEd/5O9+eWLVCQNiEHh+J/qRbfcufARZEQ6ru73QpM
4dGqMtaSlYCDFQvIsTsSYi3IgjI/CPfTGCfxzYKZ21Bl7auynyBkOqynG1kRsP9f
8iegZtt3kPO3I38q/M1bkm22qcnXKbWWm4uLnAKoyLgz5C0MK7j1KzKbDrWcwnhh
CWB7IJ621kUM6Y/IsnS+XfJhtQE9J7Ucxbli8jd9W0xLB/T/8/fW6PBnTeLTYwR8
PC92t9JNmLh2OpcCtb3Cd/ITMqY+aWjQ68wzKDL45cGuT5GP3berqfN68cvAaZVD
fkzHeFe43DW9+D9PnaCoeoIXU4Lk1IHz6rXAZr+7YY2tE8MR4eB31gVRj3T0QIOQ
oF9QviNh3iM9lHJtVnZtAf8qJFn4hiEcW4RzVOICJ1qs45XU51fs6zbawoMXeWEv
HPl+1/fo/eGM143S1+7WY+w1W/R8MKpD9oY/uG80wt36JP5jOSCFpu0PjnTWdLKB
e3OvuqVIJuM8wYGT5JZXhc+d0Gz5Tv5Inz1msvZz6c248SXXcbuym/OeaNkkuuZc
IPs5tdRxMra5kPFlm3tdgIbNirdLfBXsdjTk28xj2vaQ5VBlsGrcYsnpvcMrFqyj
YH3kMu5p1PVXrKCGdD9pnaiIESbFMlLFqW+YlsI43OMLhfwJtjFJCSfg32Gj8Kct
gMH2GAdwubPzpJLEc3BNs2oEJrbWlpppcTEXScR3ocmbiaW996/wJ2mxONUcxtWc
ueH800W6KZWolj431Q+nyT/cZCDG/QiHUHdbYB3692qpssIZRVtN+OMMM5TilgJZ
GKJQ1L0BKNuotlkd4L1kIL9eCUccpFQn/NzDRfpqD+hWDFryOiebfiEa8LMQ2B2K
04zzX3KdNCF5YvOBLJB9y/GXx3//+3gWicXZk2HnfTxLUJfvPV2m3XjopcBVipJ2
AOkNm4U2yD+RyVuCIMy9c/XVtKDIaP84rpoXmCLeBHgOk+3LoYXlotSXbtWGGuCc
/qmcGong6y33Xg3IYUDFomIjP2pAc5Vmy+VaQmrG3TRlzbHwPtmshJlX3+Zo4MRP
DTEOE8f5+doLbdSNmSAIxBQAO2umPBZydckB0Bg/1UHU8Hy4XuUlM2MczF5QsmBd
uUufj4WQt1q5xeshPSLmgdGss350sfr08XjnxQubXBOr14XnJvBsiG1l4n0a1A8e
4ZcHR6gv6AjbSYgy+wH4HjepZEz/c1o5rwZGpVYzoiz06Zo3RjCwtiLjrFHkYxA4
t8Ul9R0cFHVlqwCwaVc66esCb9e3MFGoszOxLI2s1xHNEtsxrhl5HeaDMXYD/9gN
CKQRi49wxbCT9gQnMiNXTzYQt98/uDx7kIMIfwXeIcnQX2gNpMlh3ya3igtMLc5c
WZoRTTGy1QNzCU3PsWq16o5VUncZ3nrb4G7Dbu0LreLDlxNnksIVa5PqAHbPuNrl
vje417ev4PsQFSHD9rRXvn7bDItUVsD6yRtSKZW/RSer83FBsZpvit+l1Hkpla63
8re/cnNlPAffIer4pHY8U+h7tBL3Po8BArKqOvP75nnD3yDRdyiiRo6xkSmqycQR
e13Nowh8XcH8kQLToQSuexgWEWm/47yXH8HbTbGXB7n0wpfNwTZyXbjZsknK9QFK
uVyv5LhLHporbQM9jIdqncEwgvJ+VoHQ85ETDuxQmDRr1TU38tX6HzmBzaaOAjJZ
KLCiYg2Ena/vQ0DtQyKWmC0t0K9DOUq4k+WFhryBywuxYDy99Tu30EPKpIYOr48e
kC18s7dc3B6vAbXUJVjl4AFVBmjAn+oU+j4rb78yXKXP8VIHOu/OYv7HzLPYBDtN
72j7a/PrZFlNiNsxYjYggAyRLWjXhrN4L5tPr3ySLKXS9dDAiecTUnMFTWMWJHS5
oV08gMEmD5TL6IP9IXl+b/BTsWpPiwApp/OXu+mfSWEKZAQePEPrBuSFH1hAt4XR
Y2YMR4w+azn/mL+eQsZg81stklHrMLAtV36HWpL82oEYfVafnsr0SlhpWaROwL3Q
bhGB4vc7CPEx6jOktYbBTDrvmBiVyWccJ2az1rXoPiPj+pFHtd2Ttd2pYX0Q/fSh
dXKw81PfFaDF2SErnTeLPoTYyQKn0PxBPv+/YC9JsbqtTJXB6CcPYLBwxrL/wmZL
k6G1BAF/EcY50TS/11iuxb6YE0Ohf3S6Pqj6WKWNPXxzhAR6O+JQy+veB4Ey/epW
MtnktBdAyA6LtTA9PRlzpkQTbslVMYsICyIH1SK7afnThFVrvVIXgg8pEC4bbCHQ
mTjwOIvEFx0KB1FFgQgy9I31H3oxTfE++CZpcA1KWBoYph2kQaefF9bJFykyjJ5D
bqMO2hiIITIS4sBiOoypUb+WXayxky3BZ9WMCQoLSYAn0Yy5lKlVm38Cit0mJJKi
AqxiyDAMo9aju5Zkb71nr8+avsymLfAB87nUs8OQkGLaW40wGsDHI4NFNgXf4UGj
6AuOWzKnD8jlXoZNpvg7hYAIKeoopZCUs+IKHmCVEKhEQt5evgh8smm43TU4y1KM
Cj8TP8tvSATn2Q3XiqYdTkg4iLOKVCXbwmKitRad9dLKVLfavFbehh8H9v70rJnl
V0CVHBwMNgL0eWwZnDtLP5dk0HTKG5EiozF09/Cifv59CNQLV82r7Stkmh6Z1Xmv
zRMfa30lfvWdkCWLC5Nn/DAODllMYqjOo8U/QYJ97alefp/2Z0/6Yf+yLG2mgxh3
l0HbMln7imxQPmNU0l6hMpC4sw6LuLDS2absfClKU/8OMf5/XWPYE1tOtGa4HH2N
QunlvQqlFneqiRt24OPxgmFltjwxFl9ZpMDKw+0e0VAsIMno31pr7M0WyCXgK0he
D9gIpEkcLSNIjv5HXJAxY+MZD1rLEG+3B79XbjMORewPQflJeoiELdU3qNilBAif
3tzQy2Y3jn2r0i9fuvKCT3KS9x4FOrywBte9p8zFq69z+xjF1LvEbZ3AnS2lFIZK
alqMdRHOxiDmSc2WklthoI0f2EonYV2N7U88EQB61yodZ2HlREX1gfoLWlvNfsdm
wid/MN1WwffrFNtEKfzpmglZmbyBPh/5lgJBgzAPfN3AQrw49pN3e64cRD6vTaqX
mtLnkKQ5s1ZGkVC9mFeBI0/cO0v/F774tkVx+ZybQZUHx24DZBYPFsL7pIjKHtn8
x5hZkigVXafhEK4LbrL9s4O10EZYEMXjLUxZndsRpiH3bwI3bkfDzFlOo3ty2o1q
tbMBz3IJHtyPecLrcl6VCMsZJlUOA7dFsdHCuSOWmg5LJq+sToY3enhf7TJdLdVk
f5Xj9TPLcFbwTNjRADghewBJGXNWeyXhd4oShaJyYBZStLJSGI1pC8yPx33La0V2
eHpNASNb3bYI1CmzEDtW1Yamzm04GLBpbmM+0Z5Qw0Jd4W6/4yNoB3vwE4eUpkxP
W2RHZqwFp4mtqgkWhRF8MDgGl+gG4PI/1rB3cNQ4t1x4fzXwmvHN+FOw1/9cDl4S
DiLqP6Q/HTij3t5wxeKE1+7pl2xDeau12hBv4PnKXOvvFcWtD5efafT1igD/yZad
dAZQY7b5L3vzQhY1p5CeRp3HiCTRgm2HJxdzovSoh8ds0kGeSmpC10mI36m8rfZd
qFA2bQdZ4dPhqzr2+1kQYiLir2MGI/+kJRQ564EjomxU9XwytGoLhZcHcitHA1NU
kdsHtTI4nMPnqybfs5JP0VmAB0Rz61wN96V7F/wCSIImQUOz03ykBObwIjBfSRQY
aY1sTd2GTq3VGLg+Wn2aqkYWWhnq2hTLkJ5KKqlMTNX4Ky+QxZ1edhs4Q1HlWC/b
GufSXCQxn0cEKJ/uophiJ8FUMGmfDE5jtkQbLslHx0HC5ghQ44qedyvkU3dZMzXK
D/pvGquZHfRcF6hZes8iEiY61bZ4vyRddgwxFbgA0gPVhDQKK8FX6g5FX4/nhXnx
JsEB/yh7ZS7PORJa9INbbyTWviuf/7/DeHaKXynKUxV05Ig7heachGIjGuKdAmaG
rQk7E7bwwXjzIbWIMfI5P28phSy+BQzWrjj7LH+iUjap4CMO2Xfae59iI6wx+qa8
GniJJ2oXRsZOYdYx5LVkVIOC9Wxpkwxurm5wBDJVP7YTtvltcSC7wNwyTK/Vam1O
Vf40wNDqhoERCbUIWpe/ywDJihzsDpca4UDeAmMimaHQGKajD1FaRJnlCxc1lEcB
APkXU12hYerEjivzxbg13SmNzJguflHEgCWgOc4Bc0sxRrlK+cpvEuaROXIEIDsN
179FctJZZELUTEjPaiifNTlIX+lBsurmsUrvIOCKSXY7k1+peAgY/plSWXQkRRqq
1KCpHMhy1Q3hRLrTq2+b5dCRjoGKAIf1sn9Wi1qwkhfDCJLppbVTvdVjJR6VStsk
g2PJuZWRf5TMPee79klpvBFzLQnK99xiKqmEM8lDqBduDqdH2OWwAsdobiL0HIdx
hx2t3d1z9SI68ZskVZHWFo7HVJPS2nVezimYKT/8s7PiAbFiKzL0cqHVKHY/S1o3
LJLEFvRj9ptf8tblczkuNwl9n3BH/6b7JTdZos55B+c+ytmPree1ykpzkHz+Lo5A
QKvLtHBpBA1cz9IoXiV5KFtGPP6gOu7qp4UMzPbW2Lyc+XgjBjurGzFZESAtG8lz
gF6kJSlorquP9LmJjNuy2HFOHUj+fIR7UuEBLPh5bcKJrzRb6RhO6vIrkUtKSy0E
rMrYJaHhlNrm6uCx8oDMksfGmy8XPVp2/+cw8B9+IQFwccNffi59yv9yDWDOQl/3
S3c6A3lHieeMf0GZo/XdE369o4sY3O5O7DMjJxzHiRt2agElGrwuL6z5c083iIvc
gSAuqwX5XtqNuMEJKKXkSjtAB6K3FueSDhEHON+0pmmBtO0j1wlfEcEG+VFiX5sa
QC2NZx3JYPy8b4uTGSWTHIa3qGHnV0EHnTrt4mW9mh80ZuYvShTb7DE/VjV8n7zs
1umOh/pk1WfIwafE7uORGDLKDTp51QpcxSQClsQMsaOXnwu6If2uBkDyx40lQEN6
dGghu/dw304kKMcT7eHQNJx0BCwFe6bLkvEbHQ6skmsEp5wkXemapPHO2mMA3z7v
HpFYsMwVMHwb02HeXLlTylVntjSjcfhHLaAZKYO/59wiVWJEGxIP+5YKmBAC4WMa
zjsXir3sqSVKTO+2T4Tp22TOsiB4c0RTKuFgDfvkaVaW6PE/nWhpFbEq2PwVf6XG
J/48yVQy5iPYeGlOnU5HoYcBCVixXavHqimiR8pMaO6MFVWvyTEp44aFE0xjG/Zw
DSSh9hvPycVqMnRYmnkLklK3bARZl+M86G/iBh3nzAMavfqLWsqq/KYh0bJKuCaL
24pbUnmXfOjb/zFbFkJWr5gfOXYMfZr8bAki1OmFzufxaXV48dCiDT8c3LeAP/+l
WmoMvWrBkzNJRrZD9EX0sjedOn4RKeF+sS/Kk2dG9eWVBx//GOIoROac8PrG9t99
hrANbZb27shALgp3c5O7ea714YAPJvimlVgYRfgyNPVjRcD6kOn8XHZM5cY33wnp
aRx8apdJ8jZ6v1jrfH6jVK8yDR6cj/gLqv2FqxSIxZJRKAX/uFdD9vlGPiI6Cstj
`pragma protect end_protected
