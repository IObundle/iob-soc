// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:08 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cvSSUKi5RYen7rgVHMlE6B+C14h0nNyoO0bWk/PMVX+5ejjksZrDwqAeXNVucZHp
lRRzxWI8bqrpVIvnxEFxNU6DPPSKJPN0IJhmJCS0ZR/3OGOSZR54ivgHPNs86csB
MDxIG/E8H2wyRo144gjAxh61s4io2LNyZFhZyjB+ZVI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
viHliFCV4ZDW8CQocL50ZBysSWpPrOnGdtX54dw+/pbPQbqkMnC5TFevT6JhUpHH
nICSH5SqTQ1LWSrhWQejvwKdzKSSEgkOD36PXtREpZblmgecfO0R4VGiR0JKNil8
al2ymvzaYRpPNtKdg1ypwBDEx8I4ukcsn6jth94/BPhUFp7j5bRJK8ZvSIQayEO5
yuNsV+EmxhmNai3/2v2hWSR4j5SJbggWU40uObhsPRg0D6BIH9rP2r7AuA/V/CJo
T4f2cqc1YH88Aj7LxBKPQJ5LMISYYBKFn8L46bDdJNcVwwU14ah+JNcwAfw2Pnu9
KTpx2m2SX8QdS0bpWCH9P81Wd80TfITRPL4Mtyw2D5TMmpxsMXZZq7oa9WsyS8ou
T4b7XBx52eauErUVqVFGx3EyaEaRhTb94jooNuEQ8QJUSms52m5dqOWmrpV9jMt0
tw5ED3gOwgSN+R84lX+CZYaEFGU78BTzV0T6u6vo5UbwflrVGGCavPf9+f0z+7cW
v+bUxZMDmGKagjw7sEEdpQJhaTa+//+JpE0Jl1VixCypsXu5xzuyjZRQ7d4I9Stm
W660Qpoq0EYWIAsPwrzZBwesTHPBymEV9Raqs+g/W1W2/doYYAD72z+JVYjYnIqj
lYr+W3E/Rml1EAIHCVQuJgVPS76ath37KeWRAnW6LMb+OfuMj9XH+PzktL4Do8kt
AFIRF5iCXRYYz1Y3vnBf43xV6hSMP61ML2Ms2D4kgGPQ/B5lhYL+ursWw4QvkEtC
Erm9snfoq4WjVPi7SRGIgZz2sOLRoK2uTo0CMHAvnZ6zAWJlt905RsF1PENco1/K
GUdGF1brEbKMGnYb/azXO360jgtc7ZKZDkLvvzV3b5LT5rO5DAaSSooPyNK9Rb13
iC9Jq/Afymv3W55DllsdwBmd7AxJge0Ln0CsjQYttmZy4ufOe/hPcm0f0/4AhbNZ
Q71zvPrP6QF0mFvlCNHXCmMe/x0eF5t3fPs+Vi3IWOpZb3u1QT/e7L+La1zOXh+q
pMvVuI52LupawYSMvybnbaWmIjolHY9E35W0xu7hVCTIsuoklgDBkIpyvZyhUlyy
EQHwRjaWFwGiRiHx22UnYHlIU1mwwN5WEKh9/J3gSCwnV/PUJ6Ry5z4ZTkKWLutl
Q/Gtn2X+D+LA34u3C+jeHBvO2mXHD0HaIGLVw5DhVLWYULWM95uImSlI2QyjF8m3
xVTIJAi0GuqiUrMU1tlQ7ivTAaM/Gy2E+N6COrwBlfShot9gMi8f6wAHMeMufhVQ
a+NLDo+tWjUUjU55AtJPgfpHL7Q079JITq6nOadAOurbkxrRkbfXT+iuCPiEv8DW
peQpo4o/MiZGJ9QWoIcg/hhaCgejdKcyqdUtrJ9gPfaeswGlX5BC8TTGKPtI5FnP
kGK/1O52poI8wSOE0s50K4avQe0ygkxgo4ld0M5Z2eK2vJXVTGDBAibiZNgKc2sT
HwITGBQSFjBasqHLZHkstXuzFJV/2DgFLgic0ThXcIVFtCL0DpDktFLQUfPL2c4g
fkMVmWSUQpRIpAOUhPovykHQlERidLIdpkSh06Tx8p1IIJbr2Q0LA6I1lNnHKcZv
2Lj2mil6xchUNH9dhCk8UrQ1YJ+a1wrAtf5yOkTsVd8vp/ZK2tVZFUlN4S9BuT+7
yyyfGgkjKBks8uqTOgYooq2yWsj030e5sfHp9TIUeFMpRFT/tOxqSZVWI2eqV6PO
A7+xFLZF73sOeA30iqS76EpFTw8B+k50k13dTdA0qkc5Rhxsd63KTLj0etPgbeD9
uxnFz7ABzztx5AYZVRnBanPUAFh+tdJOVJ94sLYRjph7Q+rpbjyurGrzSVZ2+ZtW
Or3090RsmOeh9adD5zydV+ofhXjCA9xWRusCgxOljYzn0tS11O8vrVhkHG59eyGj
icilTNiPfFj5M8ksjqjvqCDQsBe9iGRqn8z6BDUHKSijXD3cKO3frq0vfG7WVDOE
VxYr3ypT3S1pfnjna3L2wfow7Em0OF9S/2X5esspCyexB+NUp3k17m4xwjMSC3Wk
iRjKMF2DjYZIyJWn5RH/6g0yIYP+kbY3BjRgA/slhVLoym1NSeUEIryXUbcyHfVE
T8rReC9jUdGiNNCEjb/T/bCaA0N2Rt4gfkp99vFO97np+u4XwyZxWwugXIo8maWs
tzOa/maNL9TNrHusGZ8MiKCXjzjTudHAqm4b0Z9voemPod71fATzNlyjl/n7KJ9O
XAfwSZKWOVusmxYBgdIUEhNjeOf6XxZRYIR0h9bGGqPwFmUnnIq71Q0Y79po8CTY
b6F0X9Rz/8kweJ++26+e45wKZ3Q8z/eF4sKQQL+o8A65+8ncqDVzU6jX6cd8WWM0
M4SMxHQrm8yiXbiIp0A9btbB7Uh9Z4EInEg9XkhtRBYGni3Dy4bCzvYmII1kZ//H
Rh3goHeobaOiU+NzeskssYihHfmYZD1U7owmOnDE1FURsC4PLjaB/ftpleEHXwdN
SH0HBB9xtQreCMSIgvG11eKmOgi2eXcwYEdQMhJYAFB1r9L1Onj5dV4QtamdpuE3
vuw7A9gbfSziP2CEvGIO2WHpxuPd5BTGE8FipXMUwJ6DlK0Aa1ybhx5W6cuqiUkN
4dQt/6BZwziAnDaiPT1wxAdv7smjFX6TX7WEU3B9zYqRKjkz1LW70/S6dj6FksFj
0qgfuUYWDOVr3CeFgANwkimk6+J5nqTnzipCFrgO5oIK6J+XJRCiVtBpCHlHCAfl
4Pl+4trFam6d/uZ4Zt0NGswmeWsCZJ+z0DHMaL0DVya/SY+Q8KYozXZb0TDkK5qX
XAflThvQfUE5QJV3BXDR1bXgSoSG0wJYwWWd988qE0FVD4ke1mRmZbCNGTFRLA9c
uWOvJkMQA2LcahFfRJ54bR/miNhP+GkAOF4LLSO8xBV4xqmVtSdq0D/XifoWKdKh
zT4XIptwrB2e0DvvCgyEkJUnJSn9NbU/lpPSYjgA6JlxivN4HI6JH47SPMfojQnU
KyYXtT3pDRpNL/dbkHB2rXLOQc0uobAjfn2IwQeWOkH4NA+Zt9WusFpL5OoEyopt
lCZDq19c9IkY5WfDz4qyUNrxqVTm7iEUDhDrYzOL4h/Ywc9bGtkBwx9Saw6QQ7Lc
aqzdVabqh5xTcF5j9Tr8neSJOxRyU9wxku8FHlzlf1cUMYXiRVseiLiiR6cwv2Ss
71wl3N9W70/59Pc2vuvxfvrk2U5vEeNLNxZKRE5iLzlrNt6XOcXZ2r4ES8Dybtgb
/xhG6oT3hcnjJyH2qLvCzmWXBwy1dT4VLbG1aUTwqAfzrOCjaLf3nmZ4uRua4dgu
xs+I86J29JOq03j6SQCbkhN0AE/fVdo8aGW0k+Efd/rTjYB+AmdyQRTE4gR6DdNX
wDROiSrIPn9zb49NjJ3i6amFtFpyqsLTYydsKMKKWdOcIMYVv7WC3sd99yR9cb26
jRUSupZB3pD6hIVLPeAzIE3R1cxXQlUdnGm1pqovO2jNrdkzCF99TbhgQlv4QmH4
bvT0hDB4C/J1IUEUPMVjhMIX2t/F0S0/PFDbY7QVrHZ7c8CYieU3+DFSHetVm9/l
hOABQHysXnFb4Juq74jJQt8UNbrR/QpZ/PEeAwEMB1JraTdJggaGiAoyjJMQjXkU
FfDZK17s/dvyZ9ihtzr+BRQC8k6iSUnifD8M9CYphJRoSSlyy6P8CugHV0AxMxps
nS/dVXy1y2aIVGJnNVONpe0uvE//VSU8IkdMOoehMasiv+lcWoqJLMvMouWdYrQC
eUKgCaAYoHri+Cc2nyWvSsNqP5I1qNn2DNZWcjRWaZu5kCP/hnGrEOIOqk6m+Rug
PTwQ8/+bf+Qk5TudBuxf/DxvW8gDVYpmh9n7mPrT5O46H36WWzsZsjfrXUZbxyUX
yaDBnWOYJe8UF4/R3cPQ/R6XAJytgsIGgK3s05C3/a1d+g1XBwClQmqblqfliy5n
wSZLRv9eAF1d+jl221quby1EzS9LF6/1994xMyfwGiazQUPdWwkxk4zdkM4rivHe
MojIwUoLZA+5mjw4d2+6Ug==
`pragma protect end_protected
