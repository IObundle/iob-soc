// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:09 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KYqd8PZPUZBfX5vTaRKEC2kmjwxnWCaABw9I6pIAf72xLE/ZRai0NjAPitBsFDBw
O5JrM0J6XcWUd0y8+0A7yfPPZ+k61NHwG22NSSVJ9YTPt4UaW6MA0JSECW5+1h7P
jCxURWtjoH4YH2wM8sy+/dgcNlWg/tLy9qnFKvVq5As=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2352)
LAojG3wB5n4TeAX4OFLhZaq4EuANGVTKOaOkq/JXuPQPyr00MZp5MzMfd6wF99CB
yVYskczOhbcK563qqJ+7YKLCqLbklaC4tpDSpZ62YE/RWtlepb6MVBQClvzWJAVU
nB79Imdn/jRJo3xZ0hq88dRtq9zfk1+MVH/xBTzFyze71lqggw62gGeMGcMNHRh1
EiiMZxb0POwDUkkOxAag3upSdl9mUHk4pcIlEkLzqCja2Cc3vO+SdzvcYreI6ux8
xNFOLytx5RJEobKuHNtftgfi3dc17jKFUDtBESAYINbzEHTV/Qi4wtwagrAbOHXg
Ui4UknPnSNN6bZcwVU2Ryea32o3U+hoCwLb2PnwzcjcDHtvbQN5HDi/T8DbH5O2F
tXwRxwZGQZ6Z7Zuo9p7fbEwrKojNvR/YYhsTr+v5euKU7QEuVw2gcPwYDQTxFN5Q
VG+AK8Nu23Lyel6ztE/WkOlQLJ1VWr3oOdGZMYBIbqmDjVgdEWjJ902tBzLhxP5M
Ayt/i4cYz51m24NDlt9s3X4sg1gmTg4RT2tpohkFZn30XDMSsj6DdPG2V4GAwBaV
jYF8kkssMxt5PjVRMMVD+3Sv2eBMKaJwXTAmHdDAzvbx37sCSThA4Vji5bMMvoo3
x7Tw7XvZxtc8/n6kUZUyU1G5GsVFRkwl2n8BEZhuVGrIlKJ9sNRNUfEYDAPwkeP6
MXyW0UefBMOqqSRctC5wpchvd5Y8SW2zfB8S8omgHJozJQ/VXimANjwXUp5aLPUa
ctGcxkywDLQEW/anZBEmfy71wT5wLxu5+mwuVVQkvI+dlNa+22DpWVSCiOc7Gv1w
FuSlSfNs5oDGs3Z8erOQYDc27zqy3lGKhJo+/+Y9OhFgsCVpuNhLlK3IlFm4tIrb
OTOROIfqxTUrhJYYAAceowuc4yEjxPJFaklV+kv6qiO6FJhfg2yZlkUemx4kMLAy
QapsMBw/Zqelc0huUtnIrZS5tRroeetePiG3WW0fwJldxpEvtxI9Kh8jqP5r9wEX
b4Pghi9PrexL8w+woaz0VvmPtdaeIGAF7Dxw55iRt2/YiWQTGkNIfUtWxAW9UARk
BDcBc2kyJctSeoGzeEln9mN3bbezKu7l64UQ/7sa4q0xPbCrQ3cXvzVuPMDhk3CW
thL9CefkpzHt4G2iapz571SzcuIeZhghWkj7aP8D7WnnL6UoVB2eIN6OaNh7ZSwN
ZaEM2QbgiNQT98j9K1WUa+CARidmLjg/tCSTOQwZ81Xmoitp3LvwPZXobb6gu/qb
shVfkEt4yIC4z3QXsIfvd6a8UYuPXqGebJ9n34CPqL3NW9kXE0k6lSFmxz39jWa/
pWnA/gWZqwDYZpXzIY4MTbaYh17T3otiVdjCltUDLjAKV3qgQkdJ7tYCbw+oPf1G
dQ6SXysy8ZT6UC2Rpsb+kJmNq1ZrnaPaWqQP+NqP32M2tRVhVicBPz1LEy4yFTMt
YiELJrAlzTA3Zpzv/0V3fgmEWwzmilAoM0YS51kEN2LLah85hVy1CKgEadQQ/YJ7
5Y7xDPZEvIQ4QwbqNLCuXblav118pP+n0uPIyA4Y0o4Zhh9c3Iu+A7z/xX/EEcQ7
F3eeVKlyiQ06YK6MT4iJdk72BKkU3C4UPTNtL3iTXQ+8ZGqxFjIlD2WqyQ9MK7N+
DRQ3dqwWtKoibvNKQBjstuV+EFZFHLjrMr3XrdBg0Qvgd2QRh4Ixk9QMej7wVoAL
4nqaOgiIAFAYJyS+vN1DPLpxuJBULc3dTPku91/3opuGZzIKCIuy6DdpTfzOVim9
+zVeLoDlMG/h1K5GOpKn7Jct/xN3NEx8mDPXD6WVAIKGS2kn5nvZfLeB9rqRwIig
gCmyxGwFrqmyTEqoYnVJaE2HycJOkJIjjVuFl88UoNiqSvG74j7dHYV+nNw/j3W2
hGYU9tNfbg2O8t/KxAz23/AUxi6R/Hh9V+5IKo3xW0fBT1tGlnN59/teX++k8yh3
tBg+nMntvcpq0J+n2DlRpaWXpfFHKnRsrwahuccZ+XI8m00e6U/OyA8/k1u5y4HH
D0YAuLsxcyEsK9dWrL6YIinSttZ1nuKwrmifI+jOT3FWsoZnZeWISGVJElYNdGRm
7+/FbcYMrmvt2NsADRBq501dS4e1bb6yCIpv3G6B7PWKBMJcFDlPhKD8Jp6arhzq
sHy1p//CDjWZi30MKJCELHz/nC9WTelMhFsReZRknoEeKmbw41oAZ2fWcZrodpgZ
/hjsdqqAD5WTycJfCqJoajlF45DFBESX2CxoGfs+aNeaBOcjzaRaIt1U7U5LlAMu
VHSEIt+1rGmzYpu5s3p7aZ7aLfwITZvUT96ZTLDbMNx0DLeJ8VeAdWNCW1UhO4pq
g6uYuifvahM6IzpvmLRh8BzpTqkpswUkS2mtOnE7KC9w2py7zV1crJkVfIe4C2jZ
VL0Yw0/VmiTrTN6ztLwvV9KKYhCIbkQEB/ecgnvHe7WHS6A57vn0WWyaIpOn9n6/
FP0G99Hq2o3oac2aOS5o/jzDIUCcBSRNFEqEz18vTsBp0qg4KlxwlPEiPJX0UloD
nyj+I98vpGXR3JRNNOAaTvokDD/ET9XdfEdyaphozt5jOF0NlO2YePpqFXx2eyDj
GwY4DNUWGlORGnzaexOArhV7YrIiYpAXs2j/kVZeYNtBF7rMtcPWa9z4IirVCggn
AZdliQm/AFMZt/og8U5JQCt2PZH4YqKhy0pZs0PxUv8q54uWzEFKmFgf7PQjtk5j
V8KuB0jVNLFucK+zn21OcexPTq4gAjHkAS51ZelIB7/llQ+zN8/W9XwRbQ33iquU
mVbpVpyc5mudvQCI+AFlyCcnfiugY8KiGCqPnXkZeytHyZ4KGAeXpZIoqgzmi9Db
SRUftzNHkvi0roVy3dSsYkNJxddxR4do+Go2HrNsEhLPxhjuyca0QJ73tpQ4IBxx
ROKSUcv+MFmkRXiNbKeeaiLdQtbuwwBR05HssoiUNjs4+Mk7m494cZBPygYXgoD1
TVkFKctwfcipkVTqxAVlc0/PCyaAClMBmauDadWIODRGEHFFR02TBkgs5JiIRMqr
CuALdnWqIbcBzsN6cCv6kh+lZPTaFuNIoEJpVtYfGEUVmp/bDQMNXMwIPYjCmGWH
`pragma protect end_protected
