// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:01 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CMkw5Q8DIcokSB0+zZZjBit/YY1Nw/japQ98LdQTG63kxdy3oeuIP6TMC3x8h301
GJzaCHfGyIZ13CnyTxa9r9sxOz7jxcyhd55crU0OwMty2j543anThvHSu/triiYA
nv0yTn/tIBBS3DAvdST7HzPguFCCVMdcYV6ePGyoCb0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 54992)
zrz9zE87JYhDJDb619zgE3gIdRvdYqtHRzofoOdvg+n5qcCI1fiO2iJD1NuoTIS8
s4YMh2ZJkTbjrrVWmMQo7xZeS/FQGxAVAUKg2p0mm3qvA5I7PGB3jNUmZaZZlQYf
J7B9AZ07h9ocrF1uWOgLNF3OWnQ1ySF2E0f9SdSnwHvGEwiSPPCIQ5P72LcH7dmy
R7BwRsQaakLq71lAdSquipF2bVp86OC7JN45L/kho3eRniTzEBZkthp9Kz4Etx1w
61O0jxgfwMGeW04Fj0HkjN+eIE2k5Dqvx+HHr6Www2m7JkawiUzbTmKURV+EYJx8
IGtBPrVey8VOaA5cPprJIJj7iT7C2V5z+Jw3AKcV8+xoqNT9TScGZ/I07+EWektM
TopwqNNFZaoQmWmLxKxzKpmWzQU8nwg1OGFVLn3aThZqcganUrHbyd8afFv5FJx1
EPeAJZbG0qklZbOSmrn2leRUbTBw5dsc6Duamfa0uzn3AKRefkDxQlIBGgF1n5oB
QZhnCsPDLxwtIrSOXmxc4hJhR4J6a77RWrFksiD6SGahbGiBvAxfVndsl+tCs6ov
1TAAyfpp0iN5Ch2yyqpana+HuQXHSu1aSGCixqcrdb5c444YHaaRPNRgNq+k60Br
liSDTol3AHlbBv+6SE5TefThcXcihDMpySljtzwvKMZQSffBUDhqFzlJoUw/rPRW
xhd81RLL5kIQch2d7N4C+4e8Y7ZOgGVQMGslO5ew9cN9HsWCATa0jAsdxPc0Ir3o
EsfbXtv8fe5xppuw1iDdVSifjMstu34SuoJIz4r+y31RAPEz9X+Kj5uJG1kPYuCF
G41W4jLVCS5J8JqbATCFssoxrODG1ngEokNA2LBTF+X9wGh2bB92seaQ1bQX+pG0
BRwhnN9M/oIqjwUw8GxMNhVtlX6U6fcSvpRMxAnK5VqCYO3dT0UE+rU+5GeUvgTG
PVEj8k16BXxgfecic4Y8HL/ImISqJqT1bDkMEiVIC2ViODQqXR/W8dHpoGvpH3a6
0PbgukwgwVVD3ZSf6rof8B1LdaZ+y/cbr8X79P4yVk6TaKFc214e9e2nk6PwODPQ
feztRlieNy4vHtp7aJxh2zANCvZaptBLIIZ3+c4A9XlxK1zkZER+yXSj7A8Wtbys
G1D5xKc3Fx4J1ugK22nJDEqds1PlgIqIc/vNN2mUnZriD2Ngc/oubyqk82QFszdx
lFnwj7KF3Y+gAAXepo9pDZbRf2tur7nh4ZGlD+sBfs5ijF2tTAjBoNmPjVD9+e4p
nuX4hWqUYhoAYGe3DcuNkCrj6LZG/0VT0nRxfLkUzWM4MMbOh1mmk239NwKWF+fD
5zt2Np+i7xBzL5PQC2ETqF7bhQ45t/X/DJhlLDbhvPpwudpnXpVDvuoswAaKkNC3
eYqbf5NfcJIK0se1L9QwcAFM0VpNpYaLfl52je0QrBod+snyGM9b6P0eZRDhegJy
PHMFp+BJaXNgM70X3Mfb6egZ49kR953NyAJOgzrIhkP9RD+GsKmNjJgPFVwLc0qC
CEQsS2QNlOO/pyXQcgRkIXf4F7iCwYuQGGa3Y/84enfB69a/4gua3nSy4Twfd6lB
di5Jnl6sONs7O5PDXbyvFkAjH9wpcDOTEn2t+GQjranoWG4OzxNpGwmowOgiry4g
Kzs7PzQSy2lW4rYi5JJYesbKxaXMGwpxdQ02EjgCQT1Kg0k6jV050dzoLKeUSqQc
PW3j9xNAVSlEKle/Z3iJpUxgp8F1sIgQkImPzv36BSgdoBmqeS9945s0zhc7VzNl
fvSme4kW/2VC6dzoy2+RuvABf4ffh7Nijvx6enlBcA2XasCTwYLvrBok2nDwV76X
OsgW+WuZamCivGQSwxwiI469WyBKBfoPPnP34ARFhWkpoohVBeVnM57xWfDIdsQv
YQjbqo6wId4TLrvqRWOIiL12e5fFxvzWTYSeH5FLPbb/8WyGmj0MRw9MQxUwl+2C
iCDnj4qL0Q2m5bMOBMkznvcNQeN08cAspMggWEr7GE0o56nBECXB9ppgz9EZ8F7Q
3YAyie0/xcBnRkw+kmpBPGZJJ6ltS0HJfu/oDOdBk2fzTfqzRwIT7S6zMe1693cL
4bXbocUzsMpa/ozoWKh2y5KRjLsAhXhPikVEtf1aSykEkyPNV8v4uCfiVrewDIxm
l7aQa0SJ2wBBn2MoTrxNCqmg/1VQy31lb+VXV8zBkfWIZ8sX9zrcHHYSgciNA5+Q
gJgJPkDnETf9pYRpF9m5haQvO5b5kxN+I8/RroqH6xgOswXUJVP8+Att3eRDB6wv
XKTd7mHO+aZnMOgqBLwpw06u2aojZ5V+fZ2EaSB07zl5+QRX0stpEYKxbcJKnsmv
7qwOUiOrNqtqL+fEgzufag3kzPIoiGErLV6rTzTS5sNN7Yr5Dk9NmCO+/hbLgUg2
z1h2TncVHM/8qmjQvBiiFpzcqsRJ2YyRNc59GZN+vxPFKD9mtcdyXaSP21IjGC1c
alyhwETuSN3QqdNOWW9730mcWi+dLu+xuL/iMaz8m38VnkRgno8C5O8hv6jt4WgO
q7RPFfypyzGs5cJBuA9OBYNaYSzMzBGGeyGvouYP9KBire56jtXxOjycKRnzFJpQ
R/Q5ufO3r4UChH6MqXSV4k/fFpfzc8B66NS9ZWMb90v1Tob23PIXEvp/3G/KRt0X
2zckPJ6tZF9Cek2/UAzdCKpkMCKG0K/brrJLIPyt4IewfP5KrBuzekSd4BhLhvYa
NLyNWiooCzPzPmREGOGPX8frdBYkORJYu0MAM05x+bVYP2c9NFBUDx6FB6sCEdYb
L0TI+Oa4PugIxLS1gPNcPWPFJ8fz2KM23JqtKj+WWzLOn+ffNW9Nd2WP7bLDrKrp
xBeHGp/kR+bDoO/846BZAv/L02CW5TS41nBcXxV9cvyqS9z4wcop/fVTSPdEAQlZ
1FbNXe1uLXcS4LWEy0QGBikeOebDXmASpBS/Ig3H8YSuNmaImw6lT9Ksi1JrMVHX
qqk4447TxYyUSspK605deeiaz6ZDrkOMz8WBCqzTeFK8ApvWq/DCtr5dGIuKzUqs
LjlMSobyP6s1LrbidQVX+1zDythPh8tkfEIB5E7phHJ6t6IAfyo56BceQMIC7e+T
3MLonozAMGP2yu1r5X3ZfmMswibAXcI/kybqxQINGsykOUiY0jqj3CmSxfyimAjJ
p5GDVBdHAoXIIGWcj/FqmTgdOiAWlZYT9dN8JVr30KZWUrhO/TQIoAwj8pN69ntz
fCQQ8nTVL4lv2TScFSQIX1FG4twIuk6Y/EXcsB06xGwCqwLCL0cnOrr/2K6OT14O
ulcRI+Fjap8z95kn8cjpmzs5Jtd4EmYIGtVRagZD9NDD+3yebDYS/DorXB6/B39Z
K3WIVNqlq7Ba9bIgeMFdzxamOrrVWcoXog87rk0ckQohJwPHt41f/SlrTGIlmObl
qdIA6Lgl079W2lRcMerSIhMwLP746JrqXo/WYEVjKFA1XtpXwSFh61wzXaSMRNJq
PaoWqhd/RbSrWK0//Q9qDMylN+NARIkzUCzzFTWe9k9039JBkXRq/pLhrwTalMq1
6F1RW0kayK1kd7THwU5xOo71jbkag0ZU5cCi8LKw4954gJHjGG5mUGV4eei+WhK9
rA64k/KIrWgNOclKb3qdoor0LllGqocROa9nybgqk97bYJm2eDjE92BuVVTUrI24
LnPf+2R5OdAwvLu5MbOWGQh+gSDuei0GzP8zMPZQPFlZjRjjb+u0tSrx4Wjlfyd2
keukDhnu6NNYK+f/634hfSE+G0Ow0jVe0xB34sDphhmHA0553od0jXAeAxeCZDis
4GYuHRpAQKztQttG0czL6G1ehlj/mV0QgnNC7NgknaECTvfV9uWRaZu/0LZD19mX
+JjnNGNuQ9VBPul2izAvALUAj60ugUHAIxhAXbGeFMwqCJU/yYDDsoB3iHZOlcK+
sZADa+ND4RN10vk2EO9rNPbUQ6PApmzmikPXPzgjaBk0zCNESueZtbQEA7v9yVQP
NpEbfO7K1Xe7hLKt/KUORBNQVC65q0OxdX5XilyPV3mTYmGv1wNaA8WkLQlIJRTQ
DYyrSq3zxIj1468nrZkJaqNyMNhH0mKsbVBPyY2K2rwHee3s/XukqnvhTsrIfumZ
g/IyAmeoSHbQe+bpb16ttGAbC9JgBrqy3aNuDXpr040cjnlMRQ7gg2Ut/NeptuvB
BcsyQ+3PGMoxCoU1eKGX6InEzErxGKLhux+77iNhz8Mk0UuusT7j4i1dWFRrQh9l
ZIJydulc4Nh0/fWwSntxy+6noDUOKUnO/8O74bcytKX8aO2iLdWNtmrro0ZEenq4
poGq7QkLBmuUy3W4xFEpvcuTuNF9S0h9sYTvv0LbctqPOOVA4M1eIfNmt1684L48
D1MaUX5MMZrLZRo3uoRgUyTbs81t7xboDu8nzS+grcGRZoxAgYZgJlnRsLXH7DYS
yhRFXWjSZ2ipE/dNj2LZGxB4lA/JUtiJJWcMoEMrp+2HSCyKgkFv1Bm8L2ciYQwg
eCfKMtv5Xx7PM/oLmlTJ3TEOXPgUr7irkNGYR6x/DAhpYsnPoLhAiNZ9Dg8f8BRD
dDgSLYchWpAW5wTMJB7fs2P7hOSbfZ/choSQQtMAY983IWUXXCh6oZh/C6552E/y
FamhkNam66KkmYUVDdQdPbBZj7I/ysvW+SRFtqrUBlGK0Z9jW4ggyIJFu5KUxp9F
lsM+g1k92C8vkzrbTgNFsRvrLLeAbRURoLbKEDIq75WdHE3sZXj1jWo2HZkFWhoO
fkU++GnrAGOl5FARq4tettlbNs4mqIRPTUmTYL43g7C+6PyC3kzbOwtd8piNGuxK
z7FgrAAkPoxJs+2svwLt2gNcQCudJuxw/lvcpG54RCZ/fMxyADWpbiY4RxQO1ct9
kD76MD/vkzj+HxgqKwwqHI0H7bkXGaLqGmP24FG0IW7xYECW2ZjtJg8a3Q2M/vR4
hrouwbICE0h9sVXRwjrgwyf5paBpNwP+LRf91dN61vZxesRbFAWvYOfN+pd6+tDb
1ZJ2PiEg4GzgdXnywsTen20KNDc4/IUcgXc6Z+6I6GqAcqqUTRYuKry9Ah+W/z7e
wNIslE6VnVElnd7uJoY92qJtWKkjDwYcdK8gq8/3h/YPicRvrq62EWco3VxQcann
AVjxXSQUKYec7l4H4Z7Dvx5bzDa7g2ZN5KFy/hLewEWqHAvySXsUgL+ioySUdF8E
bNbZ9K/zsrJVqv6n8DgwIfkLT85n99kRV6ylQfPBeq0E3LxhNBPHH3Vh+pGEH9nI
nwxzuvzpcRg+nYIayeL73aK48iIVf4Op7eQgA/fU9dJJSPJ3sUr+ZkQbBECy5sLp
KD8wxU1MkC2/v1ZWfEpg9lvma4PzYfQU4VUXLTbzYA4NjTXiyPqb2PKtjL8HYkFW
VFVsUoCO7GwRjZtbTOJJfMwdWPKzR1xcJEyDb0A6OJIo0rw/s18IDdWK9l10ql0t
ipp9mPUHp5t2Qytti2md492NbYpytWNdTUpCelC4t5eEnd3cCvYwYwXXJz0TACWp
KagfbfcvaJdNSf0I2Oh9MZNoD6WNn3+yYToZdounmdSpHKwH87OFbPgLS2yLHXFV
54T7R8yR9USr4g7ivMiIOq6PU/zwar/IPsZlTLoTuDkWtWHWxZjDr3c+OyWuSjEC
3vrihRlibAGaw+oulx9mOjy9O5bWBrDd4H4CROxfxYhHCU2hhCaLrqbXna7/q5CU
gx61BubI+1c/G68/f7fjSe4K855TG0tES12VOOOTiiD6o4bCKIGX0M5SFXogrT0A
Z/EqyWETdn3j9dJkJaI5ZLennf2jlFRn88gRx4CPUao6mQ3WXbORZUefMCt+aqHj
fI6w/G999oAtkGbGb+OfERBsQZ5GAf2cSzqyHkEKypYwebzojNDih9+2fiZum8gy
Maa1+Uyye/6zqbQvOoUcXkEPL7jaZn5/kLnCq2+DmHBTiiNRiohme0/YV6adrQM+
R055y+dpnhOunP/JpgVHR8arTWfZF87JmG+1FK6Ls405qNc2rL5CUOAXRGgzAyTo
zo7t1X9EHIdQ/R2NbNlFb2w3Sf0wHgGJQ6OkdGDc44ecwwhw9QqnRG40bPRJQuTN
WCSBjCt+M7D3UvRF6+q3jNOD8JWGxm0WX10b//r5BferwnvG/ILTrhLpuSqEiDXR
KYGjOfvjShy98UNSd46A+6yRYAeZiYeBGzGOzEywMK4trZpfSkpPKgydQ7QHAacK
8l1KJMNfr3K9d3eZfZgCVhfQYGPvpQcu9EzbtcWgN6huzLlFguUgtxKhEmlstgtC
Vjob9FmYiKIijOgQAVnrbIRSjq369fQ0ymk/UOsDMGxXhad32Rvw9lsUvHqh6ipZ
TOcyuTv+0WFXwOR5Sk9EnQaYh26gWfcD3mYbg7XvOp9N1GnMX0Un1HXLzQd87U86
lmrN46cBBQKaDMfI33NAaKBeWeS34COljoyJRSP4no3IlUIhsEMP+o5LNkOEspDF
VTGg9sXYNA9BeqI10p/g7mzuBFT6C4OFsCnzAsIrEw8ylWxxBxQ+IjYCbnNaRMg7
dZVocR4Ts8IVxG754Fb8ukBdklY3QmBH8EhDNgrSx4XbJsDbS5OUKqWwJuLEm3nn
MYggTAWSf3o9PkChEtcAykzaC4oGH3e4ExUoWNKX0lUBITofAlFiS6cYmseMAyiu
op+gBuxyLlFuaEIZ5L4/TrMrmyey/bAfaheMTb6f1rREki6s8k3kA5eY7Yp3ZL8y
6AwRdwJ3vgn42M01D5zLtrHdvq1xZdqtnPrrzcPtueMRYXbJfNNpis7gYiaU5lqh
2xrgydXB2FWYtppF04QU3zh65QHoIwjB/NFHCg5LJjxOAAE+cdW+EPDlPdvmTKlm
hyJasOxHEt3GY9wwJHyCwYMWSRRSmVeq7h7NtHVk5pg5DIDeZB44TC7UaYVkCChO
LOM7eEE2ffSawDcGXhsAvhgsrPAKCazPkIzKmH6w+Z88vLctzIcDwstbQxPXVD3i
YfRkkFp3nuRkvJxPjnKdagxQzY0pt9MmxLbVRVMQkVqNS3mzHpH0hPKkAzcpsQbS
yiDUj1JVEiN/Fq/LIGwWg9WOCYZItfRUxDqo+B84PsKQwS8Jsed7KHjJIQkai72x
E4CN10Evy0thGPk3Wp+THjbaLnI1NqjPZUUAJiEMrd+N3L4f3ObvpfbFcq90+G2J
M3j2ar9t4LT2sodAy3lm/a9TVt7kyLO0YSFWdVS3YDANrc2tt0rYuOCet4C+t2BX
In980YNK3VFVAoTRrIVWLRbxUX5UYeCk5zc/I6koi9A4v0XfrC3qoUsAYnBluXZ4
w4epmmPNmwOJBxwM9+SGmHQREBiGH6FNOWnGxGCa6B8PnPcKxhNDjhZrJ8pzHH3B
DEdwb3xuwZbUQJQy2czeWl9ieoN5wAA7mlBmF72Hcn8ywcxrl+Fj8vdLC36Hr5+I
m9nuGuUPiiakbZaJz5ewbAbsrswP4qS140SuORU5ONTVB4VJpynUTTG+uLIY7bvZ
hZH+6Ddz1jiHz12vMy5gL9fbQBDbkLBjrgsTVLzs9Chy4Obf6urkhzPNqmplLzjT
YkWcj0/MAEkmkh1g1WGGQqRC+bfPtoZWDtdgp0hdgQArNIoiogn1ZLO/N9TEjUBk
fvIOtNmJ0gDehNREu5WowT4ilbcgo4JbgoBfCmbygVz3HaZQ5D3lolGgMsolFxQE
7OCxgwkSjsrAZraxAjRHf8MC0sm4WvGqSdkBWFS/L3EZglCm4wD6rrba1h3mAs4f
1JVB02jZjICefqKaQAVfzKnPgx32z9iH7rlavWHaGftrOHwHaS9jsAopBUKXwwZ3
/Fo+aKuh+gOoRItB9gFx3zaw94wS1y1beDTxUyZZk0RTiGKKCivmI9uwnBEA8LSr
K4s070eZNMA0+oGWhiAsaOwy/Z4HVIVnEGUubJE1/mCE9tlSuGrwzn6ySsdNR7ek
e57IdYntWO26m9M53+OAX5A5A5rZ1UYmcri5q+YE2KRJZqhzLBe0j6RewOmGf570
PNP9Hc+zFHEhqq3b5WUPvlVW2Gx5GAcK/XBqBrthxPsyhZ9t0ROoGnbU2vHmY6IU
r7eZo1bm2UcObdqctbjK7/zOhHYagAQLNkFRAWKwFwo4id+xmJdC4Aq94FQN7ane
E15ENjktHrKcyRY7BPyTj0v2w3C3OmuhKjtN/7EfhO+31Kq3+Mw4lhU6F5dETTdK
xNZljSkTcZxV/x9Ruk2SMrpyDQmh2WwjF42nTEpTCJfD+dTHEPpoKTlPzZUEYoNi
C/WiwPQTRbuJGzgdlXHLNmNsJ7ZlJOPsjEFy6mQ2Fe6bQ19cVBUrMZWZekTFAykR
OOABJNJg9107kH5He9nd7ptVPt8C/n4r8cjmjcgyYl60B8FQy/N50ayOg1qR9FAi
IOvjvvw8xvAtoW21+xlq/D3gXOvQFD/xRAFOjs5jsmGggd3x1+gaECI8wc7oD7bL
1w5cQHPxLn3xJ3/h2HXlnOLm8a8pA0kJg0GqgmUt5Y9n7opWPDs02Ny1M2uVBizR
Y1m41LiG7toCGCUxdONcAFJdzA4XyuyhubWhzz1GlzM07GB7jGPFo7FJG6nvuYxG
PD60nRJxgyWlH5sRLi4G2RxQRkOZVZoKg0q+0y7lrL2/qeUI4ylcCCdAhIKyH3rw
x29dIjIW26vhNvx5oBvOdOJoUvHSmuvQjep3RKbTuPBkJV0ZK0QhDJdyBTkQtrJA
YUJaI8iPjRaYbXD9CUv+8IxrPuoqV3V0iQaSMY/maIpadctq9Gf1zs6DFTKISI74
sHxx0wqbhFBGVAOT/WIfFKGWBl+XlUfXmIxB5JnAcFneBdh2DxZnFVYf5oSpP/Qc
89YY11VPoXzoyrT8R7sh/+zNozcphSl/zL4A018O8GKvLW4ftZzc7+KKX00I8VOK
2sPtaDHlh/cvAkS8w+PF4Ea2LiAogaHAdukVFO6iPzbhN6vg0nsm3jIRzEo/3yxk
cFBnFQ0xQfn0aG9ZRnvcuxrP/9UAWVxUHEz/NDbdA3dKd2jPEWbtcDQn72lvoV4N
PZHWgd7WtAkpx1nim+S8qs29YuyBRoLI51mWRiSP51tE31J/TDk0uTNN51mgfdaU
CY6eTKB1HUk25mFCoMaFZplhV2UTFx7bSMXsrVY4mVGtHNsTis90mlZThhP+rcp1
XH9xlCG7kxFt/6sf1a17zv1xmSduDn9gAVrUN1dHBYCP8TD77geFDfgofPufX+zh
R3vxgYg8lXK3GqdtWzWtotq1H2VUyOvsQdFdmSDRD7eJiI81Jqlfmwl7ZF3XK4kp
b6nScFfdWbjd0aXpSbQ6iJ6rQkMloE07fvrc3y94iP4R8kwKSpG1mFGMQ1zNDXjp
EZmJ21On7xnpV7HXSrGTD17B/gQDTCko1yTx663nFqTL4/a7S09QXEsXBTnF9feT
Tm/PNL3vO2p/3pW+wn7/ixwrzmTl9C8jOWqeIbnf7sK9WoNmbvi3rPPoe6yXOWVC
WnEGt0agPkIOtZVzp/uJIESuGUSAqjOuN5Ok6onqGy9FBCjJSWipnhxeC23qWa6I
fc/nBN8G0NbowNODprhHf9IGFXorZrF52x1Ge1aMnQLTioLxWdcHSwVOAkpzUcCv
M+eUbler46iSwP84b2jDA8xsWqAPJ8pdToaMeNZelNcB7ig4MrHe1qPNdP31TeFJ
PvzmAdbF9TnjnJvtHQ2jRaRRT43hCdonz99HApGlIrOP3zc0xpLaLw9QxueDpBnv
AB0Run1HDZDZYBF6PVEYLwuQPmLcCwKSKMxf4WPw9kWEAD0mnDeZDnLT4mal2dCf
QeDR3J03nn7KCWdli7105YesJb3LW3pJRTe8ghsn/tDkeYL2kZGT09DgQeiT/wo6
1dF7oDAARs33jByfNcuugxb4xnMcn2R/dS7DV89nzLbVJv9WK6zo6qi2efjVtfwj
wii3LyWsUckMeh7m5UmOJuRhD0+PS88yloHNguAqZrKjdhSNxKvAQbsd2unIr99w
3/5O3Qgv1pmCPob0u26dnSp0RS4UhDombGBGK9F9h+TyoweNT05t3/+xQKnWilep
NBJ3O1meGZuKBlQA/1BDijF9Al0+CES45XNxIE7Qg4ipFhD5T7JuHYji50hGaANm
7YT5sQxvrGMgllh2Ponc3llxOCRXbUyKeFNGS1T6FJMSjhXtyuXnml9vzYSLzEEJ
a94KPZeipeMRBHgSeSIwtjjS5jLp3nZL5OIpIGylVm/zxYWq+Xb3ZoqtTzCXfaPE
GwkqpWnVlH+KXE87tYLjwktlFQDdxo2w0PMd0MQqZsh8qc/VrbvKdFZ6wM+RwckN
zUdJyLHdNHAFavkKFttS3XstQZ05DIvTqhMAhuHVala9QniFBNe8whnPqmTUu9LR
Hl5tB00IYkm3zxF1qkk5sb2c6kYQTFrfq5CEo1AhMIlDrtpk5Jt8VenycQdF9ua8
hS8J+TOS8nA/TEgJxjuAueCNC2ag5LOSeaTiPV48WkK9gTI/obd+6AREc/gxdlWp
ezzuvvQ92t9X0fTjUvWzE9kdj1e1owepibX+zvUrnfUrZbrOYRnp3TxWFAqvWKVg
euy2gcGuzmaK1QTN4Bqrjs0djzJ8z/ygfx0IWec/eR3ijKxfjHPEwBt1GuAPXIIq
ZwlfiAonqx7kOr83wFrnkru+f81t1n1Z9xCc7gtqbmkDLC/Mq62/rYu8pqU51MOB
AoJSaHC2ABaPJLzM55ox7LoO6+Bm+VxStn1f6YkA7J8lDg2/5f1w+jHSVaJLL75s
b/Pr7HwBpdvsKkjlzuyJ07PjbLBr1TCNxnaaOqEHLw84twC3SIF4ooLpViQ/YRBp
cfpfV5ywKZbdlbbhS4pj38yW59N6w5ZEOv1qXXTiq8/LNTf3cp6ll6plgZvfVIsz
Adb9CEgN3GTjPy4JZoHFs7iUy2mDGdp+NSp2rJZOsonGk2UZjyP/n+t9Dso3FvJh
9gTYyY+tiIUgYMaZyEYjf+QTwdr9fsEN0m7m8vWoFY0yrdViX5y3r21P+kxUiWgf
qhcx7SzPCb5SMab0hlJhF/afQJY6mknfP1q6CRp9K5ZJFmkNDJNFLy/PvB1xxjmu
vXbioLd5ZBbyTL0K6I/W/3Ty52uU5A4J0QXaVvBY6NafHYtaXkXfixVmT8QKqfqV
lSIK22TsPsAPN2svaES6fDJ0+EmM6+78Wlr2V8qdVPGf++8qjWA7WXEPpxxkZMQR
Ro7QIoNvF0kvCWIFcHehXfHjgKfhg/2cgKxLVFdCosTZWs43VTX7h27CFfIBU2Zy
UUGSPOI6ttaxIfr1Ya+13ZygZB7FpRjFDZuMhP04+jIAhULEpqctZa9T5P3/K9Gh
a26i7hXRqf/klmdKrG4vNwlvQ6nKdyHy0/i6e+job7YAkmjP7iX0la6Rm/xUDB0W
289UYJYpWBArVo6eqZlxPj5HQE9W7sWuPyMT+SKpcB4mo998tNpxdp1W7jnc7Iq0
0RZu1EXJ9HK1Z8V6eoSpdxHFL/OI58x9FX3u/gryuokT/UNcbg6IjzspvdNT0LH0
2W4S5q6PQyJJgepyxD//RkTJ2kly4ASpLN9ndYDipjKMZ8LgHpBvra6g24deRvPa
sp4bwRvgKMOCahe5ujlGNgQZno7C6ESVs0YcgOlrnjt81msee/+ocSwPwA/UgFQv
n+NH1T4dqEyVYPerbKv4siN8fO2LjTpOEV/CL2vrZtNNF3NCdQt+nq/HorMrrp3t
vMp3FnMc4V2saGftqwuK9N0a786DuiKyDNXXntROyE1OxGU5Lc8/SuyLQ9nrhl81
TTb1spEbYL7OMgubIJUaWrvUt/fChiOa6J6iX8TkRrGYTkxofn/G9TT4WC7E9jZD
8du7o8lu+k+KnQW4JVK+H4jc5BD/+G+RmAVHOxUSDyKY8b7MtV2N3tOJ1KVod9Qk
S4f127SulUmnD/lcnqcWY07UqEzoKr5aUsbNjWtOzHcZa6YOdmzOTIwr8dLA1XHB
/Ez8IzQqLGigiMscDjZzupCEIEF0hVTXXo9u+MdZDQTW3vBsiDPK8kN07fe0PjH9
09sYStEA32o7p76FY8YsZgNTaHb13Jfw3C+Yrgo3YeByh4EB4cbhIBh7EoE4mY7D
ueB8LCnpg9XVy09/Zv6+b9SBH0+DNqslvzyf1uK+hfG6sxZ+Ua7mk/TsfhWkUkjS
GZ1GL5Ludd/qqxPPM40FDEx673EQMbR6D8CEdSBAMbNBI0T8IeGVzwrGxQ3WSYed
q9HNJ8LrriHCbYZ+u46SgCBZ00J112Y25HAOCho9qfKQ2HIJsaUeSkvbDCjRuUFq
1PVOB9zAgDGAHtxys0vEnQoPuhd2ifzhv/p4GGNcaXBksd8JO/WZZn7/r3K9rV6E
EOnS5P57dN+09OPv90xyPFeF75YXRRnA01DJYeIkWHLA5xaIQfAFhW9khJjtwzam
lC29uy1nTBYoNy9iLdEM/N8G/YdK0c2IXb6IlzNxWntFzam5YlE76ZwYtZzPzFrc
fNYWO3aC6asxq+qU2uRnQR4RaFVFNtjajjcnq9MEkuWCNJOOgarThAzWoNLuQAKs
rJGv9NkVULMlySyGo6F1zWXfVBRv2qETEKGojvgGFc6m7HPj5Nl4FZxAO7en3O8M
hw7loaa3deWcsCNL3OTMxdqGlDsj5i4aMJhE1wk6cubPb2ENisZcUXW4EiXLdt0D
NT8XKAqHbR0WA5ZH0F9nP0jbeIKG0Ihwy4hIDhW/CEEE3hoW6OrAStawX2CVJ00w
OPVRaOnn0Afh2QTCuzqsh3OT6xGEtlIdxdhd+wERkqM12GJ7Oj4VK7e/KmKlVxi8
XMyE5dY26mixsPfWzpMfwH8lgFXBEWb2XVAIMYh0zrPUutEPsDa7UE0MYyRnsJDn
NaxgIwI6bI7kgVYFtm3ZI/M7RHp3neh75pB5jsGcUjmbDZ1z5Sz/+CDFKzGPWuNN
/qfMVIP4KaI1EQ6Ha0m8CXhDO94AV8t6MrHxXG9VjNl1TNtjf+zzmL1s2lQLM33p
IwatHckyTD8s3WP1xOhBs5E4pQ2z9eEUZS9oLF/py2GjIw+NvgVQrSg+Y/50GBJ3
558RGZUffpfKrgGJ7oCdEFSCaULecC/Y7H1AJahkPrzANwGtk5awReLIdUSqVLrg
QaZK9GXLTzfslWwsBAiyAcIADkpyMB85P8VpyzVrYsrDg5/ay2FEENmbef3Tybtd
mAjs6PHPM9sqyQq4Xb7hM/fjM2hLTXk2+S15p7GQk3LqdnzCBPnekH6AyM7BnmkV
CoFA0GiJYRbn8+8SXxmc8gnw35EeAIvBS8UItOTzb6AimkFeUpx/KeBbXZ02EVyp
o41ODgezkMbMEcp+1PZrUCkkKKOHNN2brDJ2Ik2+yCddSxVhgek+L2A+KAV9EoUU
YiipUnTM78jbmWlr1zjyAd36St7KCxyM2hPRsvwTPb1wKEuujPSTREJEV/sE9x5a
yt0A4wsrzz8hkfpwBMqwiuYKn+I4RLZYhOwvTAVsX1bUS74AFx/EKPAfy51xrfhQ
wsszW3XSr98C7uf1ljsj7h6M3ZDajbMOYrDmlbGvtG34OYKuTmSuY5kXnfTR/ngY
SGq5GXa7jcDeOw/ZA1zEx882MI8yAN4HgOD6wUcwFj9yAVKw5A/zh9U6Ex5IXkeG
tfI0VBWn8Da+lPh8x+gNg39/bRBYDJQpLJErr0q8/v2rTtPl1CfrS/b+0utKlAtX
exCH0OHPQhsT8tzYozctO4cWBnsXoRRpXggEqneRg2MH8N53SPpk7bzGpKbMyz1v
NHVUvbeCkrXzC2inSINhlJD9OZf9B8rfxN0YDG6ojxe9WNjKiqZSI3Kt3gBRkUl5
EWyURblV4BPBzquKSIB9ERuytNda2KVzXU1VdlM8zv97DzwoyliMYX1oPuVXwqw/
NWYXAigAAx1je0EdyncoS2qXgIQsua8/d8qgTFUpXKtcwQjxJn6jUHtpzwukAz9m
NLNkbPp63Am1FPbtTa0UbMDjqlMTCHTSGiKd4ntQTTtd4LyBBy2lQZooRrst7gDy
/LNAZWY1Uf0fB3I3eC/IKUClOrYQlSRrEv4wa0xhXodiAL3zM1qz2rdte3mZX9VJ
r1Z49GMA8teaL/hxRbgVcn/Vm3eUnwiFDfFItj9CQ6BvFpezWIqZhCslTrO/BmWB
aXon2IcSZxcHB5I0k5mHVgp2sjwSFuha7eRxppPXL10o5igj20SmMpP+3cZ1EqgY
J8G+t6+nC38NSNdmShs26Ldyzgov4ejsVWXUW7Dr5CtJReXPI5xnDXAUuasYDWNi
kBgMe7MS1pfnc00iWl+rRtNqYLkUFxwfpIpWyYIR1nV1BVcnFJ/+ULBG/Vikovgv
SJJ06sTrBiiT19Aq6x3oLK34h+4zGdkDVGeHg8/Q0zkaEA9koZfSwee0BW/n2v5q
sExJjOXZHWhIoiBE6dhp6mMc+qb/pB4jo5DA/jBzc0Oi/fNuqKQIBcvzvJs4fs6r
tkllds8AhF5Fp9tJ58CgUCVCijka4wLITy3t107/K556s7W0uJ7Ff3Mtx/1hFOrM
m8CBZw4LGMWN+M65byN/NlWfIcftJrzPlucsB0Lg+vBCs8vpBMccCxDAXHlwsVOL
B4Zjc24KpJt6pFtfpkrCl+GcaN1banM1lnOsd/RAFCg9ZmRZptCFXPmdWDpdlOQu
BmAKP0AFVqp8wQ0JfA+Dyqit5n0jYIg0xY7G4GHHcR8BL0TiUlo5HzZLEjc6xZHr
/mEZQU7SkzuVOH/237u7EOoExcBnPFejsRiKRpqeHB00NAVMG/ROf1MstNZeZ7iG
y9b4hsQtMiulersESnARbLn+ncdqpVa4IXlNMA0V1iZSrUdwI6yFS3eZH7o5HFyv
a26QgqgZgj3DXoxJjgKDvPbF1z/Bd41UWGpa7WP2TdkhTPnIDmjhTGAt1VFErfMh
lHOgeKDkKbG4Q9VXsBzX3ufL95jLuk4jnc0Hpz9gvitGE0lq7EhT0KiKP9IJAyC3
hgj7GGU+Uk29dZcRmyxcu9bQQ/dks3+2TpYToePiS6Sfr3l/KPquQ9+l+XeHJKqu
r7elPKw76zz5ZPk1pULwPNpBbK8wnyK9qBnsXaQTU9biOJx6lhAncnQjOCR6kD8o
SqQsuDJM4xnv1eVT2bvioo6mFDMEA93xhQ7ZtkQ44h4uQsyswDsCEmlsbuPquDFd
y95IDx02QpOuKfcc8KTtWbkdsIUdiZlubPne1YaZTwi94OpLG48YxB2YQ9VznRtS
ZY/emGEFFs6U0HCgj2iFk3v8SZ9gnAqHva44chOHJxkGYz9tfpwreS/LyP50Jr3K
XbEMHM30BRRfWkBoM11WS95CwpRo/UaSlort2EhxtT/kyKCpBR45lK19ne4mbLQx
PjCZZwnGJJ2POC/NCmC8Xu73kaah7ZC/5Mg93wuD2xrvVGGFsII3jDjm48hWgYDm
sqYo1hIRaf8MfbO9XzLSdFb5z5ILe6oHI77zOlh3vNIdJjb4ccMXX80yBTDxZc7n
lSd+RbmDfgYo4CU+jimlcUan8IsaPqbmiGhP3B0xUEJI+cfOte/4AcAGKjgOH9yF
G7UluOeaHgcBYxllx0VkSwYMstEmXyugSDD0mSHPoJjEOQPgusqcnjHGa5c2L+an
l4ONr7wr+NXYkyn4vmEVOym8xVGvmDFMOBIZqvqOF6MpicM3HuMr2ycoUKFwoAnO
k/VNI0FKs1BrZTZrlYvYTFVwzv+9LF5fd0AVxW23BYVpdf3/0VzD6hxJJoz343bQ
I6ATZv2HYFWAwsEnje+eF0krAFGoqB0uKN6vJqHVNdmGrMhmfcqi4iTzU1yMiEt4
ayrpm+sKxIzA0YJSjZuG+MAawJtG63FVW7C30M98qlXyjE9xctVZ6fxFWVhAdNgC
k3HOo6FNBQ2XB7TmvMLLKP7hSQ3O9NI+XeXwvMh9ZzM6/ZkxA423WOrrOlwtVb1c
Zf1F+NsgHTWSvefOPNB8fudFjKkoimpvd2RXzbeXgFXc1v+BAZctGm72Jl5G/gd8
2yghj4KiPX1G8a8VpJJk9jKdaBxPyyAtc6mnJJMbE/tGJps/zMU7rSfgBkyDBBCI
9QjmOLQvmL2dCgDFl0885E/rRD2lpgvH74sTB93yrTZ5hPYVlxxlm58mQnJR6u3d
x6epOUiZNz7OxNtaVJ0XV3vCK9W+GLZsxmqD4LonPhhb7TzbtpERd642YHluhAbF
+Dz5olAgqLFLDRxigTx3q2mrpc6/1xpL/3ukaP3KJEoXwUnYhXxG7xax8hmA+g2N
kJ1NO7dmTNYXlJZd6Vj/JYvQn6UjLDurWPH82DR2fKQYGVcY+aIRpk5+FirZP/0O
3hAkpUJrcwgqsr1/i4dlArFhqdAsp6K6/qfZaZBiQUjnDNRRXKs1tkqnqIZJZxcS
ZXKWuox6UFjhBZ8pLOvaSyN3drh9RWijrPAf+TQwT7jEOXZOQiLgYRHG261h2Zaq
AkSMnE3lvprKE5hU1GNzNOJcBHfNxpLPc4k8tz0N45C+EGuYMKgZ9OMe5ubvr8/h
uPqxOzbtYI8rH9zRIpW9q/fuUlXGnl/OCBC57D9A3K4wTwoeZW5ZK5Pu8oiza9tM
zAEHypvskGKPOkDO7BXKu1aavSk6TPhZtJ2Ead5UxDe1bcF+SWUHC272M+hrZU0M
k5OJ2aJ9v6TCgGKrlq49FmFubN5Q3Pi1mQ9otrecjM/jrd5ptdfuVKXcBtBQQrY3
bRGwn0laA03cE7W1AehpryZK5DE3p3e3X+IwTdzCSwNVvTYDFbZqUNrK14Q/eNV8
672LUx9eHMeylZPC2hLx+6pkYx8+RivOBBxgFxxtlOXRoe02pMOuO3xMpRkVGQhU
S9Q8QhDjS1rFe6Yypp95EC42kSRW3NtwGMdVHDMDbX49HeuboRG/SN7YacmDGlJR
bQ8OKssXJP5IoQnTPxvb3b4Dj+FX3zOhXmOp6HZeynTYIHIGjJzQqkn9iEKtfytb
8d9zTsr1wrAQBTZC1LuSAxYN+ZQwyjfzLTo9z2Wd62OUBB7VQpQtWYlggI8y0SVb
6WbP8/dncS9/miLiZgn5uAaip+k4iQOj5iAh3d9etwuYAJcSYvZGTi3DKOLblGfA
5pzcOVDylGTCVXgR1Bkq8waa4yx34pe3RWuMSJ3OdorHAr4/QmzWs1tB1+AM2eNl
5lkswr+/Kvbfj267po1e58dae9T03wlJArQqsPobRk/aWbyhb2d2mP86xbR2oI+G
bF0x1WEiaz4uxP+Hphwz51Seiz+XuVD4HhjAnajVRa/ct3mJr4VHYwH+tH+4T1Lj
364sqiU13YjwrDuxTBGul0UwGBQnNZtv0AcmRHmYcCFkZQ6sJkG0EWbjTodhiJAd
XLt5XjPtIQ6Gv+miiJftNI2z83OkCJI4AsEtJAoxalG4TicDpNousGp6YncncmFj
u575jkHqebJ65eINF7GeDaQfTF4d+/5DE2rpAbUOpQF4nN1V0B+TXP6raGQHT+7L
G4CXdWiSL5AlZSQ1k6srrw304znsH3xl7rQAzVCbCWj1iU+Bg2ILUzY2xFHOjxl1
nAjLBLq2sxFMwzfzdPcrK9evwirXnJlbQx2DPH8P2VQihSn26+E5A4Zz9pXihLbU
wu2Tk/dxvCPBp8kr160XpdqNsN5U4xMJYEl8GW+r2HX1+N6cfwuDUil6ZyNEhjZ2
XuzjKntvQBTwRPei+anks/w/unXpY4zWapfVRQjJZe60ED6OeIIT8ZrQl+fMJa9n
BTaG3h7BSsjAtHj1NNGs1eXYWddMNlLqtcNk9eSmlVvfq6LDbmB9vzYXhmCtNNvl
dFLIZIuDtrJrRRJaZXq4ZrKrXMTCeo757hlIMc0TTAydRu7TnAJttyYhfyNhPN+S
aea1xnVeXm9WHEWytSPBAKzRzdPzfNOowLfEpKHi2eE86+Bw8yJr43TxlVzLrmlQ
lc1UJt3/v/dzcp6X4cMbbZyc6qGAPKy9CAC6Wv7O9LDk4t7B4IxqxeiJiaUsJGEm
1UsYITiRfnsoEmcWh1d6rSD1p9Gypxabkr2pVwnxj51qCEei3/QxMu+GGdPb/bPb
dZfEUduoPbI9CP+/OorAkeTh33SYGJa8S0qCKxf37ukdXccj33EPLSFXkcmvOF82
/vmeBaLA+8WM3mF9gRx8azsoLyByqRzjl5BOrRMjh0GLBWyUP2lIVGaFKqmeHaL9
mxIAyhlXDmzaogewQQmly75dls4nslDv0WR5QMf8vSBYfscaQRbHoDh1Yz46anc6
qll5KCQHPtVDLu0YVcBRw6qlnC/hRL8/mLNofmvzPJ4D3jDEuqM37VJFzisbwIdB
53rUzsU3zXUX2KxX034KJU08XJIoZJVx19DcLatqKOWIcsFNMmKaIFNO49rSj2vE
EdwYRgvcHpznsPATH7Q4SN+miBRh4T1NpB9sTp2Tg1mU0KI4SN6G+OP+DXnyoEdf
JY07XqkjaHO33ZL1mPRe/GpeUq2IjIROKsCogOUEcvbrVMD9/FFfksoFoEMbz346
8Kvc7oFlsNtss5//mclvO96RDn983Ag21FcMWOzQcz2uSTr2lrmGALi97dRvT2FZ
VZqe7lC0qiV2H1GxkSX2COqlccbYXbZn5lSIV1yLvwizGpnGOd4VM7AXy90+rQ4Z
819sHvCAIyzJLon7sx6peOwCrir/1TC6+1CcI2lngS862iLIRRDbtptWcOZdHQxz
WhD5aytPXYOQi3/GfgoK1OnkVMtq9+5uci3hWGtC1QrZCoG3hrJMa0lLK1kxZPh6
6/xT67iJljxkVkGMlAdK3FMk99/++K5rFSM4c7GCZp3ZBSluoilhr/sV8HulyMXh
KMGI79p/Up/qWWH4nwhi2J1b7WEhiBn0NGkYu/ytS/1hzZ5BvJMVPu/3bfpsbpCb
CrUhQpPM2Di1JFJDsxI/n+10bipOiUkgkCvFtv+jVKSPI4HQjXW6ZJvF44TcD7Ui
CyrzEsd30zxWPUgOD3n4agzko52bx1vrByEHe6LC8biXLnyvns239I+9gbbdb4yx
6d9Sbxa1+n18SQIeWRidFQa/+dGvw1iddtjWz1oGMZdMtzJhSQ99WbUwsJiWI2AQ
lez+rws7RJ2VvoipO5SHum2lbbYh+dDQO5aywV8hlaRGuGZkyHI1ps0fVDyJTKLk
rBcDi0kSBjSMNBt5PKM/QUrKdmzxVf7J/XXkhbrNspIokmAyOgKLZKZwMwkKtWA9
BHv1SvLqFYXOQLGn41hHXY0qq71qdyvsHrp9vGD0unwPh8BjyKAFePx9p/RC88l9
SSMJyLp4qCDZTSzhhQfn7N8gInSHPjX7JbgGtqT+8YYhNL+7mDWORr1ZLqXzEQQN
oGgvXdgAfqomG+zzwYHPWXBlsi/yI9pSnD/yfrpvZlTlpnUs2mcMTf3QTUjctPvD
q9w69UCQ8c6GinG8hMljEttCd/yLcUs7JkkETrF6dkXIt81AGChN2XmyJY3CYldA
WLZVcJbARfB/liJYC3ZKgPrdBEQJicQQFor+j/RKIVXQ1aPAgOUUMKIVzPyRj042
bfUag3KuZWRm4EqVf3wvLzDTKzEta/josAX501X0xcp399D5S4Qdl9K2+q+QBIbr
NcwZcojuTZF9tQXxRjq5IQmezy3GBp0+SqNdrT41h5mYzsZu/ZBO5LRPG2+lL33t
75folRDP5xg3FyOK10xR0z+he1FvDCtGFdX7aNuSmzcuVbSW/t1CTGka3hbjnV0V
gj1Lh/2keorPFlvON/fcnI3W8j3wscA5K8ZSaVF4gH+dz3i4U0KPFvLfJmV9GYw5
EpiyfIHRIrwo/K/o/0ftJUTzhmDWwENadPW+678+5MvVxl8haqTVMAAzpBcENjpC
aeHFGM/FNgHPdsMxALowJJK75j1FdRFZ7r8g1jBVk1r3N5YGlC3D9WOZNDvyPdwk
iz6CZajcZSaO7ow6bGnzQ19gh7qHFIvmbeWApFojuewmnJSUD6kgXa28MVCRscX/
KZNaOH9bAjSRxKoMTnX1PD63Jx4OzTiuW+8eArSp6msOFFn1C1nSDd+ySVDfYQlD
jwgHXfvmULjGlUUzvdF8LmZoiwvZkuyzFxt5MDgl1ZNILESHBZQ0+KZHHF9HwCDU
U+bjMggvBjPmS3xVcyiJaVbj+cbByDmTglgGeYnKQ5Pu+jYz3V7i+2t5hGox4YvI
ZEBVVwj7Y6eK48YOi5TegRGFgTTRflP3g3wpa+azA6FLQMh6XfHBCHYRnf6sNT5L
WQ4JYpjbnvoUUBUymLS8K8X0/qrAlNwoZFCDKwim68kMKwWJHNBzpxo82VX/n6PP
vUONlvsx0jFVEpOED58KJjM4XaEI2+9Fi0iHfUsZ2dbJeEoxNM/9zwpU0SyT278V
lshA0PPOYm45XpvOnI1e2mbBPPboLlfNZU3nNc7uf5J/p0+i5wHJJfXuQcIyv4vD
Ybya6rTrqQHfjj7JtVJxzGEBA/GASg+fO+11ioa3ebVlOizyPuRI/rYxGp9vx7SI
aqg1xipJ5rDpJ0QYP/i6QNCeuUZ77ydFJ5aAmqnlP+Lsc2powiDf3irljI5gY99p
xCbNoRWDg+0q8fZvwd3J3hhmu5vRiqSm9x4mVMVXHgSfJDOWw5jIb/q9QeR/L7x6
tU6zHmuDGiwfAfNOhRLfIBwZ/OLmX33S/bBqwCNRl39ZfQ5WkgAotIMViSgn/QYX
37dn81587T+C5goA1l+X0EZIuzHbt0YQpAA7hqkbf2hRNVaDTq5fXdHeVu7M/n3w
qLnlGjtc7n9u52CrLavYWsOdzMmSmxvZhzvcDY6iKYOmMSeJtebSdA8yczR3WiFX
6SiIdhn7HnWWbNLdDJ9NfAijuquHtZU42OyAKkHtczdZSbaNj6Dj/wPdWhX2d6UF
muaBCJQvpbXyGA3nDuNPr2HHzhk5mNGL4M2TQFcDGfhLf/DZzTNyUUN1A7zVv3Cy
jfqUY0ZlYgw57P8GyIWM0BbrziLBV8y/P8YeffvMVVEyZQC4HdzcCd0rMYZfigYS
al3Y5M5nXpNb/osXEViimbJpNnLPPhnIc92YNZz7Ba6uE+TDva5jf0QbTo+DFu3P
pVtzn962sk+8J9kA9HzZPQmSKczbLCXl5vzIfULYjWUHWv19t7z4HTiYCQdTOGea
m63kU5rbTpzzjrX7K2l8LDBlxNaHuy/UFJ0Gt0LwvHdaMnN1GOOn/9pAN8FP38DA
DIHJ+TjonUaP4Ys5TxOXkXpRQSop/Nz83a9pYlHjLuSUQCv2B6Phh7y4JUWX0EiS
Kw99qREqHb/qTT1rgZvj5NloAFZmI/vkvS3h1TAVittEvHKIkNGDGNtfi/4FWM9/
z6F6+GmJYXVrJ1rneKxBcaTcI7BOaD79LFPN9ocA+Cv4D2mSakRT5g+Mneixdqs0
ADVjt/VckxCZHEpbdN/3he1zRPrts4C3aFROzdUtlnhN2FG78lXuWqfDihvZti4p
Q1cWWwl7Z9ZLkfgvZni8SmuwO94n9IKI3gbUqcTKy51sACdb9tJV3G7gM5vkcZUa
Scg355P5lFjJ8htDdtNlHL9XfKOqZ3cwdk1zA+q1P5Lk9OtgNiFdmNsf2rpC7/kc
dZqVPXpLkt7wCIhyV9jO16UooFXVXL56RvPlxPeIKLnPd5r1IxB/OlQVGPNn4AaH
d20DiJiIitzr/KgXLg1sxkdv+J0swyM+UXLIH3XlPwnFoexQ/5VA9gfKjjlTwJ5j
0aQCF/aGjv0+jmSJtxAjThZSd09bOG9HMAbWMlmUXblCT73iMsWvR0NG7qxxCW2L
70aeGWOlOca55i36SHlJG94zPkpzbK2ZX1pwv6+BUeak32vMdtMe7ja+oqY8YbRg
29y0zHtqey24cHZty7Mn9cU8o8ECzYNMLpjmGoNRNCcYzWASz2HsidYfZFCaKZXK
Cln4Fr87pSngCG3HdX7ZnMV4NiruObnFDzFjgGAZPDVMgUcpmmpDl2OsiJNFufQn
h1SiMPR/ZGuptTztZCOx8OJ30TWoef0HKdwDa2DnoZvtYYXamqPAbJu2cAWdNrXR
Wq9lnRGb1G8PyTiMiWrioxiFHHCrwmw3GxbG9ZipsvOqKXrwyI8LI90YS0rP1S62
HovirIFqrquBV2SGjasSPOaZPEAiZ2pivwI/nysaEwb9iFtcTv3WfCYsoYdFeB7H
hVuqM3oYlD/rIfknRHthNHhwzAqaPmqB7in+i1f1fJHLxwbTqzxJF3Nataiezy5B
jhkAXCVzt+pBOVrmKqm7W/m3GDBcC5VizybsTpaxNPD7raNfNFE4XLuVxxy4WyYY
+kv4m6B9JaHxxZ/KLlcaCvubaxUyx9fEzj8+95APXgTGPkcDySxBZ9Vk1VxF++lt
19blMgvccSB5vDfUaStiHKn7S9jaMhS9pSslmCH9BHmXeyxZuNQGnO40iAen9Oi8
EhnnPTtXFQC1H9uPT9ws6bHX7C7hD/vH2+66/oOERLRZfr8nP9ZTZ2A9myyse4b4
Ac4VkSbvl7xL4+RJct98FFORcbM4OkSBiOrxt9MeLP6a2iJO+mwWht9fni6bYaMG
XEdDQ4bsOQKGTlHAlqzU5IQxRJqCx20AV4AKcr883/f5qtv+ZAcMzyxEFugBKwiW
ZFV2va0kq7R13YFnmJ9ae3nydDBDGma2T6yySu/TMrpmtY6zBxyLk/lO0Yu9USPM
g2Ol9AE1llZEbP03LDHCYZmwxjaABK2eQhgMfRL/S42VIB+skujIF96AG+Zop+2Q
YXuMiVX/+ZpE+PHaTFdRbncib7GLAATiQ6h8qmmAKexBc7mqefFVcCsn1FTIkCgw
A5G5QkTEg/rMKUvD+j0doStSQQU8Ur5ZuvwTytaIkPKiWojZ2t84Fh57zKDTBYpc
qVCbxTkQt2YZQdfjT/+v57G4FU+FWgOnN7lJOUDGUQGLjiR3qKKww/I4W4e2kf/t
lVQ5KOmrNPxBvI/FhcSQZbMrlaDmzA6nbOj3ypWfcN/zWgMJuDuWngpJUrqVaK9y
GoB5iZ9gAUgA25qOhnmaaEs1WTCoWuZUDHBOxUmWR2VJPmNsUqJCZJLlw9/mraSV
hIZxGUvlQBOn6aLbrDoCGCC+RlNGLzL3l19tR9Qz/cuvS3wnMTZU2EJZgL8uBVSI
R7IqavA/GCrs1D7w029kVF7gRroqbnMEDteb7RqNN39xfkxPH8wawMiTMC5amnJC
zc5upiZ9tCuY3lv44/VRPjuuBOYd9roED6X8RTZK/Yi39t4HIeyeK6wwC2WUgpkd
snGiLapluA8N/3HicPR+dNEF4K+FJdjhMJdyR3GtNGQ63cZJr3DCn0W3mKkb1L5n
czMOY+IDJDs+Ds2yOmZza2LLdgdJYmtfyXN4IegZ/2S7CYJgbPkyHYK64NyEofPI
c/EPc3lnqO72etJ7LxcdCBuZdKXIQayZDAPQgOIir2Lqlq9bcwZWXSuHYIFA1Q7s
B1fxVyued2qisroU8WHP9kCM2HtSDaEdv6DICsu/DV2K9nClqpo11gLzWBbIryFw
RDtGFCiH5IkY9UE1ajEHZhKS01+Wfrl4iGdwHhsk4w4nBenJuFFnJ/ruJXYE3Qox
pNNLQ27nQ5PPx7N/ztjgnQnDiMwWt/+WMhP50X/OcFkinvpmvkdo1ycC0TxW6+S4
svPzklgBAaKxFORwI+Iia6pQqwTeUHqp+T6YwA7tJhignCjWh1WXIAcdUlTSbvl+
zNAudm5Vk4kjiimlHsPKKLRmZ5v/eFurPA7jQH9bbVMKghw6nGzD8yHe0CI1EHCL
DWFOgaDVxWQJcMiO1YelsCz5QKMtv3ZCXB2RCorzkCXg7S7EmdqH+zT19MzyoR8A
N8xinm4NtmIGv2PJjJCsDRnVczf04pef6fmQOoLmpWuHSjgd388CwnnHQLoUIcF8
/GrtuUjmRqInvdVE/fi1yNIVfS+njzMX1bSoRxHoMrB/gGr6K0ujvo6uwGy9T5ju
8gtn1p42Q1bixoudDeUEKzFBWoOcIERS6jEPv7odko+gH5ovLzd66RycqVpL4jn/
VeWX8cqcl10ZA5IeweRLmZxoYLQDqpFkpk6JQf8lEWcp4juF69qdnfQ8YxtgFQEb
y2Y+k1amb4dhkciSajUo3khMJTRMM0m/PakATZUtueYN3ucQKAzHtBxeTTeuxu/U
DXbMN4AnNqj1hiG2P4ZCqlC+0Knemv6HmgexWC4a2BlV7fe8oP410CfI4Qw37Qqx
zh4IOQ0dXTmC0OOcL7C72PFYQfeC0AQa5PfilrwvyjBzfmNcgPd5TE6otRnxmh3/
/ODP6XIQabkoMHH8BY18A3m407zLTSjhNwQw92BEWSePHF2h2sl6Tow63sdIlmG9
cwKnulV0tO3cQJJcG1wp+eYcRR3GzaBZLIL39Ue5WI+8/1Hagl+Z7U45/OaC0SzW
mr01zISkZivYQE2+efof3/QnzhjpvzYVcN2Pb/kWVW02zA+BGYqgv34RyZhADOhD
/WUd3MRPPcIt55y48A2I2DfM/2uOC++WlNnaMjjYPPOWjLaHONzOy0kCecoCJ24Q
1JRvC5thR9F3GOZEAidC7op2hsKqO6IszwL7NsrR/oZ2kDWq1nNO7JY3y5sBm1Bc
lKUldrjcm7zgam6WF1ZVWdUoQAY4EOO4JQ56oRpE2CdxOaWij/RRw5ZG/Db2qLo2
HzdjgK+zxJ6nFpmJ5OjFTtDAX9qiLJ2MejNgdFzxgD1fSLIk/jzKnP9AH2U5tAbU
+1OhetAYPO7TFkZR2P/YkL5PRsi4MQJrKI2OMYv01hu78GKGRYbfOc2BShz+T4/W
zM/cmalzeJJhO9JvhjLcifI6gq8m67G7/tsfa/a6YGPIbWAKZiwFxunyV0Ytxvsc
rk/1dJuAZ6zngGJR0iswss4WhkIbHYGG7TiYB8iLPTeV8VdFRmypBqTy7GE4VDPn
Jp1PRNP2+O8pTZ/gUfy1l4vr5M4JCSBXStptpbYx2jVB6/IhnflzLeacNsfq9HwD
btBiN2NjdG8PapbFtSeqWq1bYpGWp+CqBZhT0Blf9fe7FsocPtD70v0x0cylVSqB
fJgMhG6ftlA3GOjBiCMwjvuP513flH5zTlB16Tx+l7gsttyU8nb5cAwhqonGK+Mj
Tx6C63lIryr3gkXEhRCOd6eNkIGujAiSEvqG3fFh76mezl6Jylve/dqPCPbiVvyb
axxNaCEZfAEVx4sNY6bxtM60mvjgV+9MXfyNY7fVxgrsCxnkgA73mryBGja9gZr0
/SH58Glhf21Cdl7k7pwbbwOS7P9X/ZZWLntNmGsnXNQSzc7B/+l1wBJhQPD4bVKh
yKOKB1B96O2AjSMXZAeVjGbnUbrXPUEfai0R01GmLD/DQ01/l4kXY2rIocxKQmsO
hw3jRJ5kpGWFbt3V5h6J8A40XGXwD0+04BA/lt+EcwG4TUAuu82zZKUxBOP3yr/i
StGicRMHolih6c7PDB7MfaFLryKF0fq1QEPDx0wKNGcDzjh7+8Yv7szKY//6oZyb
fm/GyyVB3Y+DeLcgdSvQH1ZIuDKSkx2rJgpenWXDj9zmjRT57bXurebGXWwix46d
GDTHdiXOkEb9soNJ3YjFjjx4VEB9hFi3yAeaYcLibn6Xf3uoaaexDsG1Kyydf4zn
iGxz95e8wep2Db1KfZdjhjpq3LS6JmfL/I31V9M91i0oSRNgtFTCPdotJAoMEsCm
1IaDj8hkb23+PD9FneX6nuS4gbmGfQh4GhDPiEW/ef3COXqnwcbb9RGhS/HkLB+l
R0rhKD19Hss8NgOAx324/NzpJZ52N6Z/pg9bAzaY8lg0rmKrSlngBkQvpwEvgasv
Sow6Nu7r2dtJjifK9iG8c1CqzwCLb6PnGI588eELAsRLnlOwY1uQ6A3x2wJoa8Hv
rNLA1uM4Cf2wKqYfBTT4O5cjJBO48fm+o+wD3SU0Uu1tlAM2UWdpkAuXnRU4X5F5
aSriWDozh/hOeePy4yHFYKfue3MXXrgYRlZUOcK8c6UjjkmtNdvJFNApH9c28vwg
86VjNOM1Gh9kxgQJtm6GQLc8qReOZXqbsqxBYQKiCxSquB/WI/5vVYuM0BT5sWxC
hpyMMYeFHqjrYIc8Xvvt78vkC7giSuZiAIP703KuvwjMPw/7tHKZRAm7faRpGbh+
JQOz33XEwWZXSPb9S7KNNlgMhQIKLAXKaViqJqsmZNR9fTkjICBSqINDIaW/gW8u
bpkCpYRxIo1K1U6BJB4WPi8SQA9sp82B1NrvIz3kfG+dUHg105txui99c0KuWdkT
5UdUMYzsEvuf4OOWRW5SHvcYBu9+K7y00TKN4++abV1S2d4qsYG6dWI7aJTrMDrc
nNDG94L8UyE0DR82pandh4M2F8T7vJ+uwzY7CtrZriamYGA6gQjZajazkel83ju6
am1y5j0qNKrdOxJKDH87E1mpXLeExCqLKtucuOFctrEGfuF8rXUnCanMEJsiKhad
sdAFPjugfGy9R4KLhQfnaYJpoMCKU0PdCy2BWQEZhW7d/XI1HTalD3T/Js9bZkpw
Qt+C4FzJCyNxpsyUFQVVXdWiMrBmu6cfeNnRn5+p+tSvsaxATHmDI2JwQAkLf7Uc
CEmy6ytw5it4eSLjCmboty9WSuxqayDLgxoo8YvV3J5kU3rnEuJ2ld8VtHSKLC6H
+v00G7GzOM8ZqBPICubXpZ5Aj5jOHxII1P/mzLiJHWTfNLEWTsR7IHyxZ8unYOM7
65Al0VoA8WwZW7rpDTP96NKgY0r8r3xfcBD8/oQimEXPjTD56yjOuL+zm8lyJpud
WvvUi+v5WIFrfntqhwno9pIttW/idK3R7JBwF0WNDCXAFBUhWzKTPZu5HOGsdSdu
QursYyxg1SrY8M8cnUBt3Oh+mFPvVgVt7PFgml02NMDa3gBwX94dVdxymFn2Gd7T
h0+0pGL9OSp8pCs5MtUv9vu4ZPzTfmlQfXgNxshGBc+Q8xUzlaP3S6hfttbJtLla
3uHLN0UaVcaYh7RChmXftHcUI1PAor7jufJyjFudywnFVlVeNEWlJgznVXQ3dDlR
NCXoffI4/077oxBzOG7Rid+jeqok2+chXTgrt/spwrxgDOLsvWKKBRgNarhapwCR
VnJHTIU1SZyjNz6y90BorQhxhkML59lJEE/jynmBQFelaRdQg+sm+wcScYHLqkWX
b4ZhUs8aNbrew4kaHKYaKJH7C+EkUFsHyKs651+oopwo0SlXQPplzZZ3od2/WR7t
SbewAPBeLj4iqOawJ0C3eTANSxBuwrLrrAGknxMiRbc+uN+XlzQrlN1Ceu/4k3KA
teNvFXjZnXiuR0ycv32dtAqHhh4H96A8UEwkw6XyxhIjrZf0puHK4EhDVhkgFE70
zBnTjejGRmFtjQsqOcTeWYHM6pbY5p+kkHs+7ksnRH8VIUQkx7SC6TVQH0y8zs2j
1tlCW7P6Fod4UwHPRDAF2pr1cB5qDm6MqSUDkk2zAtc2cDnBtxtpQaKMJTMbn6Pn
ilPfkA0mXtq9uTiy8Z7FSVfYg/5GZVnIBaw+NUpIEA4+HLQjTuqiB1EkAroMxd+B
J8JM41TLqAxtq8yzIBjIylsVGh7NEeXdlhBS4HjEvD+HKkLlEx+5DrQ6GarfSLIA
jgQUcMjo1fKGJKWo9Fywvked9PmXD0hXtNManGOcQOS1MaXAKoJk6Keixp4Ol5/2
q0pVfC3ycGtUgHGnGrRRLSTshWNXPt5TYev5khi5oE5MgYHQu2/xj7b+r/Z++0ap
wEefdtyQFy0ag761LbkA7TmVqWHaUfccGxEHEaFtl5SQHBtflJcJM9QuXmUCMK3N
/balUpKxZUOcmzPR6WlONhrURwZYwZy+ca6Ox3xdxk8guKc2lA/yD3y0GRtRME2/
zEd8cjObqBJCov1Kby3FoDL/YHXMkJmdrM3GDpjuNvuz0C5HAFCOqvofgpBYp5bm
4nKwIVGCk4GE27N0gsemlvJDs6KcqH4mEjiZBEqJS6ZCuaoJmHTm90vlQPOAb2Xb
VBfsH/pieFna9GO4RzIXPs4PIBx7Ukz/E3mAvEYB3wunrbGnCCc0DVylXaAYpp7j
64/Flmsk58moQaPAhHMm/qDiosX3RGUGLgLdRgEwUYkUX/FNek8/5Os82Rvqj4Uf
iJMn7H8CF0bWSsLMapPSFpAoezurBRkPJh0EUP8cBbqieWM12IlKdVGO0hFfqRN9
DBwhsZHJdimADfafIlaPdOcsGA8ckOsW6LbXPfLr6WYZ4WN3fi5lkG9f2aiTf3p/
Se2bcBZseyj+8w1D83enOAGtdKaPCHdjkmcmjWbE/T2xSgy6sI4SUBY0P5v2nLST
cN7zvnx6hOL+zo5t9vLyRl/hpFvwtDlJKZT0YtjH0iB+5r8ULL+7f9PVFio7/D10
tyGYdHWcpHsHoNBagCjROmL4t6EVGiauwrHminV6kOTXPRRgrsgfRzMC1JH11BgY
/uOk1Tw/x0sgXTN7j4TvjV0ncAQYNfwRGC9d3sFYYlSNuw1iK7+9wf5+PHw2DdPw
xGO+KnWxa+L/3iJlAulLChWuqbVa+j13lKtfxjNvGA365u0ppwFE+8T1CfuQV69L
rq6t4e6piIohOpgqdDDCsWrygAztjKIrmgXWeiNioPpc5cJ1foF1rxmMLkhJDt+T
oGTQC2+QHCsdc8XXoIC7BLFw+3e+O48nvLD7jugwWO8anQ67ZkBZoZzKpO7ab4/j
lK3AcJJPmQ47ORtf5oih1im+9/tjhxux6QYqtgG41Ex8pWrbi4RXuDwzwCPSfRHa
qCfHmBnTLBD/3Vau9vRskFSnRlse2Wzn786fCduKWaTwM04V+AgEKjZApjEC+VHy
zQv5qWx1IrwkL8r62vWz+paMMmQQNFrYDsg0h8PfiltDwtzEoAR5+eCORTBsFiOm
OnhBd/80H4lXZwQvA8It/IMqmdOM7LBbR7gL7J1QndecbiAq3ugraYm2c45dRjkK
Q+82cAZdTyHtgTWhMyzFLeNiqoKzAbJOtWk/j8hJ8PK7Xa2FlyNLOPlGfiH2zNoT
KaToelGroUamCXOjdz04wKdHgGApjVH6nEKdFA0mbAfEA5t/+4y8f3UHGX+HBRPQ
QM+UziMUTNBNo5fqfBL4y+6/Vn5ehCQDQHq5DEssEDNTzkkaz8C0XIq9yaslpBFt
No5rZhamNv4VMHPRh95s34up3Mg3Zkn+lRk8czGhp+BJz6Y7xmyjElKnLKY4ME+t
OOte5xeMb/v2X96fgcB13H+7/dcMGDdLjYJoqCQMfYm5AGEQcVK4DAJ2bhHqNzZv
tPPGB//0ycLM5GngnRAuQbOL86SSBc5Ws1ug6ErgJDEjh0/rlk6bdnhKoOD0Cl2e
xCU5y7OgNiZMiNjPiMSaDM9Eqg3JWGusTiLR9QdJbg5iGbKo0Wozi6kP/2XoiFfT
IjUSudWTVXU2xv9a9sTErJhAznPnYOC+yZ9Dyg9QoXwZVNWLW8T4tT58+AmHnjJt
ZN07JT1wBBoYouG11qx9aJEhQhCSNGKhEhZ9F93dkFryl7b9STzjprarjNfHDBHz
Pl53Gs9hDi9T/T7fthi275wpa8nxhYqwXcd9jWTnTa/sU9C7Bw17JdqtP3GerVxw
YGN3fmuv776bhC7XblAAjnZudWXcFHix/aLZEhyVET7BTh5R8kPYklTLL5sILeTB
ZrGrFa0WYvRMI31zZnGtKGWBEkbHDuiPzCRclIt8jqXRi4ZkMu4pVqlUqrfUoGxA
/GBGGej9Z5CwUtsXY8iyWL6B0SQiW7xZr51pH94ZDhw3BEFBjqVvnovRzO6bimiQ
MVWuL4EbW0rtirooD16fV8ZZ8zZbNMqHPoPwK8oMf/QGCGGHCNWd7aHAJ7TJO/ZD
7NWyDoSQZho8+m74Wwskxc1yluH+EgWmc9tOohoUYjbH9m9zKcHBr68XLEEVoW/W
f6pMBWLCYuXd8bUJSaxzMWEX2FbiKhpRIkDVpas51Fj8YDZ29jiQYU9DD6PXeEHt
ZT4M5cS+ohmG/X68h+kj/x6ENw4Wt9MEAnnYloZVUSiAHE2R7NY22ETa8QQIbzV9
VFSDo/BVFZUvXTN4u1U9J1hu+H0OxQ79Gtwb580tbXsis3iiEc/t0nPoCL4p/PT0
Brq1umGd8zreHmU8D59GfRXHQlzIpEIcDe/ft22yx7cSCWuvbrkBLxCsc7pQb8Gf
iTjVAIBevvABwLOZxzc7CRvKN5TGtbmNldbXVpHXvuP2CKA4tfEdY//WwfZXR2Ht
PZxOGQKBoXZM2eVSNvhk6Jywpgk243w2tyWipn858bmG586aUT17KRHzCdPDGkU+
BjvF6Am3vwXdHR/nZsPHGayYkBpQIOY9agi6HHsYsonmpNhJJAjct/3MksVL2Grs
JW8qG8e1xHEdlwfCR5WYVHkGWiyl9mDe2Tp9IKhy7XyO63AvQ2xMdM9a5xW8Ra5a
lX6xeIvhOtu/5y9BDgjZdKx1Z5AGjjoTpdch/inYGclYmQxwH8paO7gj5piM8TK6
IH8bnuGI+xE6fhYJeB6mArPMwS3RXyQNt2olm5OuxrqyOkpWzXAFF5GJrdipCzmN
XDFG09cX/dzb95FK5Iwibjz4NnyrMa5xY6o6KzMaoZ24CEhAYNdO2Wet2dbqIfkv
wS4+icTr0oqxN7zX9p0svzeZ4jJwtmi2GydA4lfqwGRWdTCsHaTHb9xIOdsgMVvN
8asGPf/WvH3x6/aJKMv0lNTORZWcJ1+h9hR05j3i07KBWFippFIn30goErdj09UJ
KvC9RRSz0a9C9pUKBMl1SlexEyI1tsyhO1wDJlYnDxUJHjuibmGyxaZl0M/Dic7I
yxQAn4OvGFKdsKevZnoOcPTYCkXz/XjZm3n1zPMLgPeE+xZXnwfG1N3iR/l1LwQG
hB5u5B2+2ds4NrftybxjZU/cwXyiHbAZy6XaNPVM7DT7WMMe5RvBn4lxKqOxE0kV
JhsCCfNNkTLTi0fa9MK0n+dsqKswFt9MNUmJTJeNU2/lZpG8UvintWRk92a7ZQ62
Vs2WblLqu7M6knw7TpHOWZBLrADJCco+pYA4SBLR1FGKtmwk56wH9fs/D5KERTmg
z4gr4BQ7gjW2sob+AMhwrsgs9oGVJ6uF/b7MX0xOmDgAHlgU4Y3KQp0HITZCsjps
PHYKGXP6oUSYV4uWaMS9TSgnty+gKK/OXOgvHwAwaRhdsNyJsHA1M5Un/8DsBncC
gfFRaRQp70u9/s/coVwmyGf1GbQv5GELrInOw5YrRfFj3gbM8I54RinCQKOTfhnD
HCn+JqarYM4ugAb05ggB/YVPbRnrtsDPzPwffktwHc5oKH689iTkj84IQvqFzzPX
wycKIvp9Bol5d03hNwXPs3Beko8mcAxALwyqRnX6Hoz414zmkbIN1Ur0f2bCNtEG
vzceIuwBLyN8M6SHuCwPgT4Wof1wc9AvuL4M73S2TKqT8CNiDox9a++NWpagDQ0d
n+L7JeSJcJr9+pnYH+iULCCf6ZCh6mq7fTxT4l/DjBo3U/qhPNbtFkpxFrUJ7fvH
6oz0K/g10G+sQmWr14kN23xhjHVP078eWobJJyfX0HfMJ9YsZvFOJvxeOLWfnFY8
vjZqKfCNo+uDuQwFw9AqLeAnDRJGGqweKGxEyAxDcSAAz6YhMUQyqpHCpOcDLcc/
4cyA7QdHxN1fHrdbOnVmIT97Qlhme4pZgI42chzmc63SbK5rld33nlpMiO/RVpYo
B1EolEtlwNo0ht5O9bH2K03Rt+5hhWJN77OJI57v6Xao2gP6XCNzTPnLpi5xMOhA
NovCHE/uoFLkUgIYtcYGphSoiKTslHCfjGp6YpjWZmY4ZUvIS6KNSO8uS3YSw3nZ
ZjugO0YegRICXfmsrmRmyNuKTcMbWhgVSVa3TlSTV6FNP4hYsOGmPonwzipqOlA5
a6nj4BSheHTfyfOG58ZUjlXJ6wdwyJdV/djpd6LLkuFT7j+ZN6k8IrzZ2eF3g90f
ANa7aRfMYvCLDwK7UPIjCqJ7MKXBr3ud/AT0ztONbXDck5hxIHFr1E+QYlCSeIO7
y/4Ei3JFgCA3Byn0hRlfJ1lMKVRldbvSRCXnhWOLwHIAA2uaRZWQW2+CVoz1LXVp
wQbeEY2FwqCgZ1Y3tKg8mbNyPcpOEvmCE7xMNZ0zj8ury+LGgx8sX2JUR3B/y05L
nxhbzc9CSm3o4RR3PcTI0raOIYxvqPrSjRT+6uQ+T+Ndpt94dcIS0CNgzHNYLslK
SFmCGAHc+u3RzN+0eaRGMZ3IjX4qfsmGJbGUcPGsUXgnPJ/k4nOIq7pNgGiT0lqB
0oX1STQI5bhmLG96BCns8kW6gujQo6ZX3ZyEekrROQePcAQo3C6XMcrvzX+ftRQp
E3sfKh8arPvC0ecayX1TGV5/sIIn6PI1gADT/M5ISCxn5Xxnc/2dAML7D4+tlImv
XJt9wqoa1bzo69NhOgLk1bHFn3UBIquRmXYd45Tsgj5nc2xvlkRZsCO0kRtfOJo+
A7iMLJoPCJ/tgN4Wy2oHb5wJeoL5Tl7Ef2Lxrx65HnS2xLrTX8zNfnUkjLHjps/U
ns2i2jWcpoc0kED4pZbKtBkLrfqKrDb0+JQTQT9yEX+VkWxrTv0kjIa4WcmVVXUY
WdUO1NW2GxueeIxGVTkxslo+pLNjZPe6ub7TCr7nmJ+r3n8n4RQZxXEoeWmKfvVg
zjs4kCTLpsXhDwXRnHaX2iP0+raaVJSIwU0qAzg8pZGt8mSOnaRiuq2pX92nqWVj
LcaeDw2fowCH21FASQq5qgvQPam9iKG8WOHhWnu+nvT5kK5gxsxHkPkZolaADYXU
Wmvhc+D3iNRZJd3xIvW9BWT7S4XS7pqN7H7G75CbkjlLyErywm9uJ5Rm496XA/IW
LygHpHlt6jtOqibmHovofACHnvUB15Z8ybGfpopejOXI3KJul1xEkKr7nd5nn2S7
bnbzI01YygMW/WLyuIgJ14r7TIEhz2At6bxhhfSqXyl0lNwu0IJFarDLu3Bf52u7
mMxmDQLSEckEFkDvuJCWfFRvcc0V/RCq2AxGZoh+K7vvVErvTFTIMnnlF04NfVFq
9cQ20JTbRqWgy0axPI0Xg+W2VVqxObSmRxzMN6FH2LRbDcACT+6PywrLafHEbndF
p8xRvHnij5N5ZTWK5VxNtyg62x5mSIMufVBp4WErE7JMoMm8pcJEB0VBLZzEZZfY
O6d2syli1TsAz0enFZhlaucUVE+nk8606jI54GKmgvsvhRdijnnFXj/bMAf+PaA7
LR+5h8tZ2fDazqChB9wVqZlF272Anet/Exxl+zTG5z4SGdNbu3NQ7jAmmeE0cSST
QeQROTEe+B4YQuAYgK+CgIRIyW7LZlrvNPNK3atVUpUmJba+8LnA2AA4ojP+QO9s
zDRQnOGst2og7gFNuYyW4Fb/1pA3FyLOF3/Y9GZM6Hofsttg+y1K6HgJaAGZ/A5M
cg/Kqa9Giyktt5C7Z+BL/56wvnaM7rthzxNGovg3lgTw3w0UY3bLRSElXGlcLry3
gslvDXpxQogrWtC6EZ1xbzs/XFsAFl6vwuOWUTqLE43G8pYKiS2OWONYKUtvDWK7
jUQnPcjTrNKgXXF/mBmiyOcz+G/ASjcixWLpz/2Ccq58fsBei5l5VdGU3UOgdE4O
F483VplUkFJpFzE2XY/cgBeJvkhPgWiN6b0HxcrO50wrYUMkJ08CzxBFTRS1ltzA
PAsH9+OCeRtHe8RViIURb7AYW9iGzJH41Tu03rUMZuTcvaTFA2Qs8EtM4xikC7tz
7qdGtHXpgh+s30z/HU6gJKNRn5wwnLBd0RLTiQQW+aekEHhb24JrMG1KjL3/0f7T
EpPX5nqVP9LeOahm7mwNsz/vPwhOdyLdHoqsSFSUUH+bSOK86CoJvQWgG/okc66n
KB4N/nzRDaNu27TPqPojf8hylQWabraBsKSKV19p/MNDarCmmfzbw9nWL50mZA40
vrU6HuR2rjSM0QOIfu1A+/NJde3mJSQOZHCTeEWySiaXzP/IIWn/x9NayBbcQJgL
n3xm9qAInx57i148sCYzzMqjktX+NVxpS652KYpcrO5JlYUfiVxF1mspUoaL39xD
7gDDLmz+FWLINtUA8PTm9PYEYFwdFM3UfPvKGIGSNYQHkBBcqdOSNJm7GRzhkAUl
GEHOjb6FOmPJzeHB1WHjd3gHT4jElEorZI5aMZBhNiIjKQs6no+B+Jl7aLysJcfI
IzgaD1FNCXiLnOecvEp3Fr9kh19Kt4ly86dI4YsqJshfdk5V8iei/rFk/MKFvMOi
fjS3GH7J/9Cz9M65+vyx9bsyq5vrZe9T6GBEs1HE2i1pJFMS1vxBZt9Fj3G9+Obj
LLyEnZH8vGyLduWSMxjCYXevSC995jq96yOXXTBwR7zi6k459bfZrjihDMUD11Xz
URZ4PxfvVoKhrbPxU7vja2wtB/4TjSYRPgpTngeMbZQr6p/nSK2B2CfE9Yh2nx8D
kDRLf4bg7AC4ltB3vHa/qKqARkiep9f5prXWErWOkctvQKF/QEtAHUEp5Dsnn1Nb
yXDkiWt9WqOcOEox/WKFuCocQuZ+l8K25cYUfIQ8HwHelFxbYYz3d2RkKcjBwHLs
2qBgiodXLNYQfO4583P6z0FkUY9lQ4v31mvWhG8k++gC8NnB/Oabqxjn/jBE5+E+
3bwzMW9SQkAnOXJFQpDOpiQbzN5f2V+bFkgBsswKKgy9iuc3EH0iQNQvOFAiJW22
vN0mYgRit+9jqHr2+RHlXENiEkrcq6wIxiCjJDRqX70tg9qKddLkK/KyX2ffbHTU
EX2fAQVpkQ2HkSUGTcFV1bRApn6fdit14Eld8MD9SSCCnlyYevhVp7T7/rDk04RH
1V+4wSWw2SmjTrc6j1TUOB+FIlJjHTXiwKKFsbCa03HroJhF/4/ZYHuSfPNzTdu6
uFpBbG/hyfqdtX8h/eaYiQNx+iGi/EE14/IFFPFCe8xOApbMNfQ7bZZrMPbNOlJd
BIORXPqrK4hX+qnEi6gpaModctrJ3U6d/rV40pKgcmXNxD+fQhqs6kduHxJ00RTs
nWvTEq8eoxJRsdOYbThauSdpSTthaThaYC0sF6gA5H3IQlXyXl/886kwz9KI7voH
/BEYE/c2ut/qtAQtEOzWt2CVOkGI2BCtZxngFsdn6SJg3dmK5jRnEqATnOuYbYMc
hWxJTAMLZDIKE8Gp9NzE9+R4i8yNl5SJ/1+Q21lAOtARuy4fOR8tlklnJDLMhoXG
o/018ZgVTFJnMyb2dSQRtvGdT/BSJKfCGLPwQps2Y3Mm90fB9v0us+cN5mSuEFMG
tsS0aynbc9UcCiAE9EZC3Hy7TFP5n6qQHVZCcLDRzkxTzaG4xpKBRG3sFCq+YDSP
seNwmO/Bim15AOlwOnrPchW4kVD8hXC5tF2p+VFjpiB0pNqm32OH0IVJrrG7J+V7
g/H0+POu5NntjiLkqYbakNouaDklpnM75Y4p4pDTBWz4FIDvZmQ7j/TE/zqZg++U
N7k7CqZKCSbvtuiPFGWgLQLJQZHIKNXsXufsIh2LhBqDQDTRobFlPD/gVKG8Qb7y
cZgmof8LG84rAk9pwyDgdbY7soq+awZoGdo8qfPmGdW6a5cXtcsmScDJ2o4N07vn
CLYn3xU8R5+MPcEmzaVLZ2l+agKbskzpPOyMNy2bDQokFGaw2Q8HgZELDDDdOU55
8IpaBr/JuVmkbZT6/JCwdbKDbLd356F55rxMi2Lo8594zZ7Nd3dv0TSvq0yGdBqx
gnjSjieffvzU3dWqDg66YVbQVAXLzJO8K2yQN3UmOKFRZmrMLapFPqm8rUCyGIne
enxkNQg/0ynQkVU2w+wWBGyprWVPqZAKy0qEM3aTae4l6+OoXu9gNtkwYudg/PEc
H3XQn4pHkeO8rO760JkR4BEFBV9WUFGQICAXJLPMQijnxOf1NMY4bghUEAafH0ta
U5TyrC9Nu0ua7m85oeYXDItELVAicuH+g12KrUvbweWFRBop1kTX4KX7obh4QJW8
cx/OOpclOLMiKCKSI6+Vgeq7+etPKddHz/G2b13zhD9W8JNT5OF4xtACRDu+057L
A/lF9auqFLM+WOI6hPL7/f5fmkT8y+5SLBMc3t1MakChbskfeitLzcEREAtvXOwS
qf2bS/tepYF4vQqdPodFX8rdDI1H7WzjxVt+S/kE8GVRU5jMAP553ZpB7j9hlJ6h
REwDb6tiq5NZtJwqorK7S7zoI/sot32ktbJe8gYhA8XWNqLNnL8NApMB6Klk47Mk
7dvuPvXZNHHugnZ/hq5I/rs1DNXR/1WbpngR/UF+g7NOQIXW+B3HhqtQj+kuyYml
nP8UnaLIodEoGhn2OVFZsK+KpwNo55KtAANOWmWUHO2D0sjgSS3YfL8ISTDbR5yr
kTsUKwqenBow4h8cxl7XLema5w+eyYAUBZWkSGmVpThY+CVKhLF+EUVTzfvH+YrB
LvJQK5XRWdwEXTPusRnPDIjOHhUbN/Z/4SZBZVxqaONvCXB3Au0TT+MdxIQB+0Ku
S9KleVvYPF9D+0dJudcWu9A39G1IQDL1/6IQEpbyfTp8xc9zLSVNwEVPqQsuLSoN
ArXK2nFwa3jUn51IzuUs6c3xJVZeCEKiEWBpjqjldoHd4B55LNM9fNaFbQGuO2FD
7EbvwBW1FhsLmbul4mJXzqes9+It97eQw61CFKXZojMgCIhDuXgeAM17ROnr874R
+uHO+ua1EakNaeX0AV5nn86hfMxTuuMqQkwTfBKXQADM+ehQh4AzmPhvg2yUQ8Hw
Lbn2x6vwQ79qgRYmqhr7PlKiCBpVwkrFupeGz+qOFMWW3HVbJaSXgp833p0dn1QK
YJsnjZTgDSbea2Ot0kWyS/0VU9iqrSco3enGeqatWmw7Oazteuit0KDYdEeuIemJ
4XLCpq41UgkGRMT3+QOUMlO9GgCwB77UCUgYLJGR5ccf67wP0crCJkyAas5ESnRe
y2zlpAfnkXQarnR1oewQRPAExMYpfSDXV+bifxkbk6qcAqL/Sgz/xaLXn6DuFWiI
Evzuhnt2bbdz1lkWBpwKoG0qaInEvjNU+fdDr6Lsr+v1hwYlmiMA3KGQl8ftTbjW
fsLq0UTeWlytNt5kL+/AyVt1FoUIY/dXC/9PQ7qWAK8BH8yYUJYiYabGlzfi0lqY
bruO/chnZKsBH4PrH82qzC/9IJzR2gTP8N4wnJ9J/Q5uAUuZXFViCHLESGbVt4wS
F2knmdWZTAPEaIFiK4Uww93/N9JamrdN9T4DT+vGFW7C4vXbe1jYG5liw1UglYQk
x01da1/OiTtvQi4xeOID/OBebIQHgyJOapmllznLAR5QlwV59YamflQff1/UY62o
nXC9ILvEIMR+xFKLlVG4iR7kXuo41N4lBfTegHaOOGBjL084bOMGE6Orzl+PpNPE
2IFP3+CTPyxOM7OnqQfh+prkoY+3gxhL2j3cfXhR53LizOJoDSKC2WEjW8nkwokE
9gZcQKQF7GFgfa1X6B8EJrDw/463PLjprt2wKctq3qAXW/q7oitCvnajdujlu31a
gw0XJ3E3xevs1yVJAX0VFJuzufU8ARyKoWFV4DnJp22ridKwHUrt9JgnW8IoNisV
M/AqPmxV+GZUyuKLoeMchoPgtC4SD9aho9yDjdf1gL1wIODziDNkZVRL/aDAv9Zl
MRDt0tNsmwLjBrIG82bdCfOsuEZ+KdIXjT+uycFK87VR8+GXhB+TdyZQ/BO76lL+
IbJ0CzurfSpANDR/dFGJ1GgLgMwauc8vJ/SNAHeBx4tmm4D9DPyn3nQIRRd7IQ4h
94GicRJDwNmVrxSb4Fo7Bp86cGBsKYMY3aBzpRaBrXZ6GsVRicFXaRSkc+sEnIOc
9Xz+katGtZQ/yplpRqMM0VmG+g46nTiV2cme8gUXNKwNryLOmRWPwFP1RDm7fVU0
mMCjo//ZK7J1tYSvCvrgP5a/aaVwK8kpLE3/95DaDN54eQiCRytu+iqxnirIFBtM
qLuAdDQDIudyKjnh/ZMEA6EW7r347H86vO5aMcAVgbdGq66orCskBfICiL1eLQkO
UBRZP0K1Oo7ea++q2LUQqurwq6hzpbR6unB0b6OKMmGV+5zPiAnvn6O37bz32C4L
sIfcpjTAACInlBarjAzAzGhSfYg0+vCZAsI/Qgo6XDZIF472+imsm+qepx7t7kyE
cH+uouZARtGy3WR/+iG3/XHJLeZH5NX5eOGL2zbg1BwiALLlRhMXMnIVGIlTrbu0
RDYz4vfprFzDnrMPg3tu/K1Ohkc7Neg/0N+4GS6gIhAcjICQ2wKbwblHBs+BNqKg
NDwOnUM30ZU2662Imz84TIouYLcQTW1YVbZHwbuB89Xx/w0JSV3BHfQaWtPk+O+F
ERv1u9MFcwfiHSdMEgs6LWeVlh1oTIMyBjzSg+CYl1sQole95LRyTQ/3gLC0QOHm
MjUx5dfb5kODYbHh9XBcUn4TUzsvJvjYDtbFCIvgO8Nywo6s/CpJ/9C/olQ4cVpT
3yGh0EOO+EBHbt/TRTAKEOVGll2NESsMfvwv+MlNnAN8d0N2t7NQgTWFOd13+60N
VfIJD2RWEkzLVIdq437q1iWTUDohI7kCUc4wVyHq483KO8V1StVUQifhrn12EFv0
WJMTtr76Ds5lbzaJ6QX2+Xs+wjb4GIsQT02b2l3ArbB1tthyvOWj6h3NSd/guv2y
N+8F2e2ys3YkAErOtKKndmXsCaIxNDUpgEwaMvy0oI2A9OJlLqhaBTThudK+o68r
Lw2a5JkPM5v0FwppMyoDGPoW4u9Yj+jlxA/iHsFiUBQXiSPO3kQBzX+wlY82UPOq
r4O9MnPRkc+1s/EosJ2MXsaCvk9VxYTv7lrej2q2ZfKgeh9jyUXziz6WFKu4+WKD
CbQqsL/IcVnrMlfWWE+hPbJT1hfTygEgOuv1BBEQOjdZ0DVnBdy+wJi5AbjklWrw
kdNOBsIwWWYAb7TW1icAWAQBl77PKxNH/hVk72Tu3Bb1Jj9731sQLXD+mB3IQBo3
9w2V5LxOysGGaAYepbJZ+8+rrkhKNHF+H8nUrbUiN1ums0+WoS2cztI5eAS6FPLd
amGTdCfHZlY9KrjhFTlhUsRy9W8cq3uKqAflaD4XbWbcxqavpIl2jeynIhK41Nus
GJfYWfPUbm4upuVbR1HHE4FNPlkezxFwJoSjIsFHeggp4dVdxpxpWve+XQhF7Cld
YW0TzTjWFcdp5aKLtXSGA3P44YiZdfpmPi16A2fJzzlTTLQKEKFPrljJzEgQ/GpF
8R/bbYzsDyaIOAi8OUEZC/R/2eKiyI0w07Dky52q/hjSHk9A+TZ0CsXvyqJvyWOG
HqI9VwHEW1g1uIrd5sTMTAxHNdoKwsUOS0iMlKE4JEv4a2kUquvBBidSy4v/fPdy
qf58lRUTBALmo7kEQpZy9mcVbyuZKJNFmWDG7fVBd6DW9QFiqMFrAICO8d3T4cWk
hLuehY4GGSuHU5/Esphc+hJae5rdSgL3wZpukG2i6SEpetcccPn2zpx26ENWoSdg
BkalwEEQkWczy7bY+hREACJoFVG07O0yAcbjZgH1bDrgdzO507S1C0cL3l/zD3Si
Q56HE3ymAiGFNCPWYOoE+8BnPI21crPMF7wmOpK6N+vatzNpK+Q89/JrOszd8Z6O
ouU2ba4+veIkUx4YXbsp2OL74oT5SdwMm2J8ePLB1CWmJkBLyEFIFk1s+XTetCpf
NkuFqR2ocTxIVz0SKE2Eg8l+P5JmtCoH4Wu/8E/YEu15CFNyOW9U400hxEhuIFl0
Tvf1zPWrdCOEsdcfpHl7/0OLlEWLKXv1cIABytHUlMo1p7lc5BNBVqg/FlNoXWqU
fUp3IYXHBXobncmTwTc2Jta8omGLgbERAcVh+J/Pfy+EVBK612KVxww18oIvCSux
TZ1vjZHM7SBOG4s0WpU993un1fCgGcdjaPvsrWlgocrW8JaRnVr+i/eHGWX7w40R
1YLsRp3lBz4xfeYMYB3DplpTnsN6o/LRJRymDkGRXqsEeIPc0FUI7jep+kE+MsfP
7Z03Bu5iLFl5q/dxJ7zBP3jwZFXmil88wVSXz43NPowSwtxzpLgdlnMKk/PV3acc
wuT+aHPhwBA2J4iq1VlhFyw7RbNI5dRmrDX4iDJRp2Qgp13KytkMJyxWmQW8E8t9
TBlaN0qqdg1tScBsn0SHO6N6mUbWWejsrbLSck8mnTBv6sCZ7yEEcYDhvB/8OI2z
voAp3xkmGeiJgzs4STcXl491kyuzWoXCyRMTQ3bDosW+zxExC55COYDdJi2+FUR8
cbtKm0M9SZFuNH78f9EHhaw0uL/qKdmlso4TbFJOij6uybJ8D6/BwvRyjFsGAovX
JTfT1eStC0ENrg1baf2iE0rViLu9xiX6IxKBmKluYAhmh3o2f7H0D8jsiqEdUXUg
csWQ8yZs+8SaSIIOeTim6UjYU2dsTbY8tBXRLpzVlYDFj1YbZ+IXEOQRPTPGN04x
OLpr6E+BGc+0t7aUkNQREYUufSP0Blf+XJxOv0sN1CZ6ryyvB/2MWodO/2TIvwLU
nmIfvTUj8sIIlfO0pbAa3Xe6V9iDtbTA1MLtsw73c2U4rpyaXLETNbw7x/9Yx7xN
RCN9aZpnhhpz1P7ZVj762HASeDFg4kZFuJYiz3SejHIfNIg/iRbl5/mT60Q0ychr
2yZfrkBVkAfua/02EHDSifkt7ntBH8DazyuuoNLcCXyLJWwLIUoGW3sFRthunVbP
Mmef+FMZjFXibLEWrtoXHH+GRygSS+1F+pbMQmHoTazXvvDG0+KitEttS/N31pl5
b9GZxHVvdBZH0eP6mRnIAn3AEQ9oc+e9nW2jiTUbyOvBG+zuG3iJSJM2hVpmw5Vf
yaZKb59RozE8nDpGSy4QmHV820/4n5vqVtel/vuNqRzpKUVoleo/Pp06bAzF/gKs
nMQzB8cOcscJ2zXQ5nQAZo4SnMah4wRmSAgXLwBkXYwfTcD4Ouhih1Z3bvdBYJfV
DOqVEVbFu05KknwXtX8UeGqWo5JLjMcD4+qxnTrz1OzvI36xQZdeu4mWtD5TjvGO
0XHd02eU3r61ka/60vr9nMmh5AX87iGLVSwm6u4ppL8ZMkv7DfBxrKGhV3JRrS46
6gYZNuHVwgXCmrna3ERDTR6m5EIiX0DRw06+YxZJz9k4LsqxbV5itBHZEVRVgMKx
nvvkrEJLhNidh5wXhHXg/SdXOZGyRfBPT+JuHv64aOMuhe9q4UXjtR1uWXZE8aS7
3hPifqlpLXsbVR9PUajnTrOWMsp+LACJn02le8o8TQaeqMwbaEfNxWYc1D3eGppo
9gPkAnQ7w3kCH1g8K5HWWhtIPxlt6TMiKaLTOSR/Y+N8ag8+63jYF7yhl62+Kj9I
QenTnInUk3Wtp6IC34nY3jc++xHbfk/cdjmKBLv2XKLiG5roZ7jVVpndozJEbxyZ
IzYSAFJQ1Wl1b35aWMu1KpEAjBLf8hk7THyHWbfch5095LWaLs+NI6HHuaoMJ8uk
bk2CWWa+98yEhuPZHVXCcoeQnjWcIkVv+sFztGmJW0vgZPxl3mGkfDv1EjqER/LB
NRDoBg1tERW7bhUzjlvoB1LrjtqStWIB/4Xc+xibhw46oL6/8Os22MyzCAWJvXqC
xThC7Y7F9mpAhXtcxubxxRx3nnHP/vez7jWyQYj4ji6/N42/os659USl8XewCRXa
T6ZjKRFQau9W6+PbEZOuHvsUTNtkd7N3mlLktbDbE1RNZiYIy5jBITWiQGK57HK8
z2EDS4M52emcIlsPgUwgDa13x4Dngstc6+HW5fgZ2jV/wus8PnJ6m4SG4mlLtUgj
Po7nB94RnUE4te3UHZMdqKj7Z67qItfL5fdiL35lecis6JIxkj+ar4COn7zgn3m+
3wVZB7wraoDrxsfIekSGNgVfVcS+aP9lUo0mD3bkJmM61aPjVBEdQ2eph8KNsYjf
vD0BF8p9wnt/8YI5KAyO0eIWeoF+nH7A7/pRoKt53MZA3vth1Q94IQqLHCiPvJoD
vVrFxwvnZ/Xb2qdeyjcpbnW3NPgMnL2hxpwNRXuhvBOOAMvyWI0JC0bKpKQB230Y
gpuKXKuXLG3g4PHzXGmeJJeTscpVcfJq67eYX0RvqUFnNsgo8et4kADxzWEb7b3K
Viq1eq2D2y08qqY0qvT1Adi+5S3UtOHPnOhl8oJd9z7//Yz5j0Umojs0JJPps/uh
sEiCEoJXV8DJIHYx6fy8KrkWcFQuhQyOtPYiBCgp7UAgmQHTqwtFq+kIa3ZTxNus
tTqjGJMrtTwDwV6m1L5M0yZ4kfDolvULwEhHLOltoB0a4rH8OwKwCclI/TVRhAMd
qotm6fUKORkVez3qyNq32S5y5VzkHAQDoDkGRhWiycChT2VvJJ+1u48qvHDA2RrN
N4+KKBTQasJFG58SKnsy5pbGFb3Y5iwfAdqn5sk+YORPlqNf+gDafbBC2bLFw0N/
yUjGXZYg7ALRoXp5z1cZ1tJYgXM0vd5alYT2DqhYHi3093sv2AhQt+8TFz8DQls3
HpXbwTou9aqQOkXYRv+MKB2GLdD9NrCvcWDr0UU3w825F1ETVFQo5suaJdDJjqLB
xAsHmIXA4J46QhGkfJO0h0NfXUtCDzx0Wa1MM23BPjaSwAqVqUyplnw4SrUb/LDn
dlLsyjgKpOBHVaFRBEYalOeWoCf1IO1XOGjBWEXol5MK3jtzX3fen0ciH9PeWAjW
1tq9SbYeLNNwHje36dQEOqqBJnq54KjoN3jWXrNXNMTdE1Qr3rsF44amqBCeS7hs
ChAaxe93HpPJLaJF5QKplukEfus8P4lWXmxkAuAsiIRLsZl0N57Pa6oteeh3A6eS
yo9pIaFbKvNKUhm7D/U9mfiIXelkjv3zzrCgLInshj1oIqXmzWRLwCJRVWNmoJPi
7I/aMtFIGiad81JcuPKTct4OGwxQIo9a0TKtJjFWTU5ZOyj6ryu5Y0uznBJ8J6bj
ra75rE1mB/MiVJZn4A11HF+dOUuHTQXeYXac4XMp2AY1DpBIinRDtvz2zkz9o2GJ
EHm+nqe8wRO18JgNwloN6MPs3CGG+jj3VB4jkdgDMyeu3h4hdPqTZRG7p+CNmfup
DtWtzsXtSU5sQWWA4gGVY40b99f1uR4pv8u+DDZ/EdwrbytFDyrIwH8zCEMUA6kR
xLVwKO+otAEH+SJ80TQfTQQCIZrjo5NJ0oJKXzjZsdrarR/FVouz+LxvXnM/YLRr
3ytui4bCpX2g0974qqGPAfJnfP+s27/gnLqdTKEMMl5O7SGNJ7P9f/VHU8uH5T27
oMtVOgWi1VrMMaQDrHfMHs2M1fcEdJyTMQ0gHcuULYHtDYCV5K+qkARIr27CwvtM
7gqsVFePbHthMJ71rMYgiCyQQFKtLgp7TZffW+2AyKXI0Nydz5+/QuJS/BX1EWqB
/CmoJWEXjC1D846cr4hyhHJ+Q2xzx5ss9JOavlk+yU3bKZ2vXo1ClHLevom9bjNn
Qh0FxtIvt/T2GwpsuxFFr/+rwzwWBdNUssKjXJrImlBd4EwppbNNzBHoAegd8R01
iBUl5I/zTqTmglza3zs8y4UW/z8PRpYOuKysQHKpwk+4tqq+u8sY2Z4TdBtgvPMp
cZD2eSPV7PctNTsAaDDo2UzFxeCNH7QhB5eMKMwLsj0vWW2r/cbiKQS1U/SvifGI
B2tbDwt1s/HyW9G4v2DC1iwj+gBTCNyKBNNsEeypSIdlRBJadQophGxSRTw7tR3k
XpskCUxWGdxZtP4K2dN6pW6wwhympJ3GFGQ1ddnDMoe9BGDIxzwzV46T2U9hd2bD
fMy+FpykR7fCECqMCGOQUIxcYHlz6aUavJjqc7EDmOoYnzBsDjOOtq06y6AH9nm9
VmcQJC6Dq9bpwaqX5Qf7y1r7cmBzNq/RaIXJRj+21b+ln+jGi1nwlfDrmfbQBsKF
uyC9EljqVEds2/aDpodYTqSEvSJGVq8s5tIOhfNTPmY8bJkvXFqUdy/+2BjxKWYF
UMdDxqWdo5JRXFwQNNfnkRhsIL1pfgQKw+LH1uyafQj3EI5z+Mq+NVS/J7JLpi/B
86Piz6cWOEHk4/cxFQXMkTj5AFJqYhbR+i+/G4q4nuza+F3lIg6kJi+MN2h9PIys
IxekMFpmkGQ7nCRDNkhcgoPPvymgFdvUDFIlFdWjO9zNK5YAfOUEEHmZ38gloViT
fpsW2yqxcOOhFIhhhhWatn2WXHidLJVTEDTeph3VQJDAae15i9yetrVR7NtXnIl3
Rm/zfxFlVdfA/rq/8csk7goT/krQfn3U/ExpUYOGYTxXxqpzMC60c9w79jiT/ZIs
CGPln+sIHJbhqbukdUXT2pUfCOayXnji0ffYlM2V1tTN9TIqodSNvbzg46qQEmUi
VvS5AfBWwjATx0FZy09oXy4HXDf4G5C6SmdxIoGaCpcx1I87frV69XgnqbQk/zuG
hmuge0NtFtL13vhJttmYHBpX4+p8hgCqSN5r8eHrYC3t+G1AwLYXEmgyWofNezWG
PyRDNaiaoZgZKvoVMVTnpCpllI0p59321p8Am0ltGO/UNV8ND7lc7FzIQTeyzLqh
UHpkOQ5aE3qDvevHgvs4LiJ39w2DPslL/4VQw7KS+tU0bQ033rliEIC8ALCQ2LJg
JWPPMI0SlwJI2C2k5BRM5plkN7wtd3jIbdyuWpSvVH5z8ucWS03nWLm3sqmB59cQ
GGn/CVd/RpopX+GbhMewK1+8ZjCFaAGFfux4CtBRqASYwQlWMCew0el4NnHZu8l6
h2bSpWAfOVcRPbWRn8Gtbc7CxtYJYQcDUYqFT66lAMwY/vHW87Ysb7lQRbLC8y+z
i4Yf73UNXGBnL/rLxEJ+tdZoeERgSuCLLo3f37+sjQV2LH9sz7DCIm9WuysQyxWe
PKW+WTAtid/5SaZhAUgigXbn7hqZYZDaflytfNqAqA3uWx+cJS0ZiVdqnE6wb6No
kpm/kuQQyN2uVyzveUhrtvmceua5/U35e9cLYcZyiwDCgiy2O6FGH9zPBe6915z7
xSy7zHj/QVLWxaYByN8TnN3HdMFBOBKOcbs+Qfhhr4u+EmFmgCsspYxfK2nRYj62
dERtsHS3gEd7MxhXXsmCklisFup16hBAW1rZ0ryp6XD7qgoxdJZDv85+YGxrNtSl
YBryHsWb7XCBTfwFyQsPcjfT/+DFMHUMh5/eKzmBc9VmTwGjjMk/EhNVmQArlRv7
jwZJ74i1ZKdlOzIxcKuUNz9HGWKnYM13UOUAzxk9OY2ADQBzIobR0DCB+ND/hYPq
LFfqLx4ZGa0AT5g5d+e2am/newU5nwN1+f87IDFJIBHMGhOG/VKo9fweunTtIGCS
69KP4N+cXd+GSw+LxWIuJ1+5xsITXPKK1m2FpOyPFHfJC/Vqf0cvkpJaNCsD1M2v
jEcTxebeKliD780o3QrWpAXv/7xHysvsmVtb0zt/QlGLvjm+AydTyhGVW9L/mFDN
y8p6ZISEsFzyIdr0fWO/aA0HSUF9lCGOj+dyZdI7KJL1orXX0utjI+2VLAIcnkTj
8YUbzKO1R86WYiU63N/RDbMFiuj0aMqM9x9/lxsOH7Mpy7tB5tZ9K/VkXKO6Sb/o
OOSUK2w2pUnKa4SUJnE5NIctscOCMN8PSoE3L0iu59JiZ9skovrbRKyBqNMZE3+5
X5fF8UIwNhGDQvDKHa+IPnj2Axq4OcoPyM8Wls+3XUInDtzo0FNACHhH6ZUx3U0k
f3NvDRTB9xOaHt0yGCWHR59xnNn9iDkBDr6UNTiWDyQEd43XxPWTbtZ4WdTX86za
MHiY/xVsWBg3kq2gk5soquZn8NgFZz5uRBCEjmDnrYoqC5Iqrc7PMtfh0cgieYWu
97URV1/5jg6FhkLxGFZttEK/JUS0fqRAj30T81/v7u3LKHQ2/mKkhhG7l/JnMUA9
Idzu6RbWCmnFmv5FbpO4EUpJL1l93ilK/XkQtfu+PgC22Rm5sBYEoRjWPE2FBRPa
MyhyoQcnmN4OwYfnjYXK+XrqYytAEphYl1FSxnz7PjJME/XTfbz/ZIYX7spws4Eu
YZEl36vRkxPovyt1bdyMOB+Gng4vXc1cl+HWZBhFeJMXw/WJcDCgvcyTXgnuWWRn
Lt3RhC3v23VHR+KQDQZOUui4lncDLfKjXWMQ+OiGWIKdBMVzQtKbUysYA85hnePp
7axAu2zBTnPCw5qmOIDCT1L6kHxwEV5Ot0Hz/XrSdaYegEascwmI0REJYi1Esl56
C8c1IAfKMIctDKTp6JWFIXqEGVyLpZbpkAu+j4+yxIbw0Arz7MRFhi/CRnGBjy3J
Beb5S0MA61uKwpTlEGaEvNyifpSPlrDn+AodhYofjR4/RmxxII5UN3VieJ9wWrCD
1cg5yQrDfoCu2KJEQJ1ab1/lt+cZ5CfZSVojG4F8SmuPB58nDrLsO/VVVK35hJGd
U3+EzpU6Ldqak56uCle4jsUDrOYNZzQBtXdjP+t/u8jzAGyABTSmBQgZZU5QM90X
1tMFWst1o8u0qjb2nVrZHj0/w9/Av2EDF6VcBw4NDzYACIPHq/oHmVfdNz2cvDev
fRqkdTgElGw2QlqXw2KuVfivfpMf5163PmO37dlVTuh4WJM/KXUf/5a3TMq4BJ2n
yAf1TZj2whZ5mZr0pdviWPYA1d2COzzXRaN1uasLHAtH3WWoJuYYFxVegAigBTRx
TmF/SRwZVtq3uBF4A37Ehg1l7i4OWA6Vz56s0J3Y/jm24IxTHa/WN5zglYaIRFFq
SgC/JMn2XM5tUXPAQ3D3IJbcdJFvhkDY9TNB24DgS8SV0cB3VIwzL92DAQcjpKzl
0QKfM9MUfp6R54xJkarGkZnPj3PP21CLSQYmoiAD/Wn319SgUamgGhtTtsh+TpiA
Rb1rtSdc4oeh/qI+m0HwrUnJtQmUC0SZbqfOuVroxg/NFX6f0U4XvubMIjzVTKKz
0AhrZEP6QA7iF5ufwuHkXmkCYYTKDSW00+IVNCSOsvjZvXdtSaxWXbcNpgCkKNmy
I47PFYdib5b15vG0v95a85pzz33ELXh7YNse2h7sW0Kt2R9widBSs824tvqy3xrM
fQORIeeuDeOLEy9qmNc8zvCukP6GtYQx2YSJRKUVQbZmst6xnwriLY1l0L+4o6r0
ErzTvIo3kSvezs6O4FNqOz1BMv8GnvPP/Mec1WrR+WT+73hQrAeDN3x5dNBawqkf
vo7tYeSkYQbbR0xBGTELCDAKfPrFoSD/osJfJBAk0dZJYuq/lVWLRwX2S+qlt+0Y
Ebm8It2TeniqLGZPVJXNmr1itYlHm/qhk2ol08bG4lngJjc6akThxyK7zNJyg/IZ
7Q8cjj4B5dx6Li9/wi4TtTRa2Tau0RqHCr+xkstfaYtVuLfJR4+ExLpZmGWOoaP9
HRNh5M9nSm02yrx0rGtDMQUjjXP0SrItWOJO1AVbvaTnEAzkvxgFVne/iLnKEjM8
vIFfAhSNTHAQ+NUzinVqkKmPhC6X/KNVI96xZVn0cNhmxiaZukJq5dhzM5vgef6i
6XfUKBPOUymO3FEwjaag/if1fB8Gv9oLDUfcywoBk/QdLVv8n4eYqrmaIaUjKngo
qiGKHeEPoAFlRqdbxQ42FGgh64pLlhEaHOiqL/EAKUYhQqEDJznCdTO7exXUBRp3
lJxJhkXyfTMb9dqvpnvuWOFfh8e/hDuF1DJKSe2egKCqxykfBSSlWIKXFAJWdFIN
obwiO5wyPuWyogw0LtFTsT0LiQtoSZfZPQ2tm5LgCnBl24UD1PqT42G6PZZXoF9z
oOH2rS7W26Yg+s4A+JGmFO75Gy7Hw8fKPtdmkxyYq0sNPYb+B+aeTQT4+8uAxCcY
gllc7pC7cc4bcip5QnUkejWu7UDCs3sMppTkMW6kvIIQ7eY8LeWdp/QUvFuKs4b+
fVWtRv+ZW+BAXog9n+rEjUV6lIe/De/sxi1B6GF5qHZlH26r7fvGlwfwkab1IMg3
ZcREntWbZuNkFTxjO0Ek7wdh3l7fSafUHRMNpQM/d35Z2wdbz6a+K4RtHPGDpyDb
2M8lNsLsh+tcHm1dVwecgwVq5HI8nB/PlKbUJMi1g89jqz4zSGUheLUMNkMzqLEq
MbJTYEvTRneBjQ3uOwso9CM4lEhulXmFt8ZUMosBExr2RxpD2NNO/E/w1l+jhhXn
QwynXT3rxmqrzozJpa/CAU2xresqcPUnFWSzYIr+UI9yJf3kt8WFIHkNZ8Qf8vQm
JQYorSTraOhn9pXI8moyZuxcAzdsdpi+iS8zLupnmykxvKF7EPmALpD62JMIa1c6
5UhDXnNhjqoLdoKuYXEToD2ib10ikls+ysWHFDp27rryk44aklnvOEMrsmW5sMH4
klDNr2Na4nAWW8Oq45HUQXSL6+Nkrqg3530NUPUdOXHQBAKJfJ7PS4HNSsM/O+km
DiSepLHcRA8da4qjaurmrMI3z+pjLu8zERkAhYd1KKwj9PA8/GSQ6/TPvBhMguWM
kOT9zv1jlZEGEjEdc2GzN5+XGbYNJdljkbT5oLctMxOkh05Yd5W3pABEiF2HpNY4
zUfoWX1ihElDH+xr95N2845ErpiMtQZWc82bFMlGgljoP4KAr+sOjZgFFjjhU8xQ
aJ/bvILwy7/V0FIYfkBHr1GY0Ay0v3B6b99RwTUThjDZqpo8OOdVY/QUFBakcnU4
1+mwPYSDdCE48jh0QxiCsNtJ97iwaQLCySQOVedcHHZKsc5yNz38SLnRsMK6WMIJ
bbzETMVHEfzPwQaTduQh2Scrr/3M15ezF0zkvc8T+jZrnFjBlzhfZjzOVN2mB1Fm
TMJCpLtjwDqKJVCieSA6Qq3e4KR1LWtoFHH9USzV9q7tWZrzAyJtqAxUSx43sGuS
/BM3Kab75fAu2wsClI0P7ehNd6qeW8zJ0FXtY8NtpMOKxmrkOsQLGFLKSQ4rv//w
bM0AvwlStmlSRV+1eYcfqM/XeOYVbk6oyZAKOxcUc9Ej5c5X/kanOlTi9gckXrWr
3VhIOqkUlonzWswbyeuaXir3CetW7qoI7EFpFfGYev5LMBFN71B8AB1g3rg6FzXg
nDtVuJeIr3/JJiuyj9NAC81en0fjTIH0DkY95jKbuE7K8cFXgOpprzmTEDXWCpAf
TS1oNbT27hfKFOWoQwkP5cwNALGHsHdgjijDxvRZKHS264LnpORMBxSslF/zrhwN
Gnz6NRI5A6Gu1Apvviy8ITuBEL5N2Bo9AOV72aXlGCoIGu9mK6Vl/oI4CbtOmQO9
kHWBJ767x9i1bOtaQZCJ6vEwX8I2Egalu0X4ph/vBYVRVk6pGuzEzqp+18T5kWft
7fjB/pndtYwXaXglmF0vjB8NPX3pRpIlf1iQN6z6chg0IwUIz7EIJkvX+HQztt4F
QTjqyjSUD7jIETAWOoK0Lfxym6ZNf6EB9uhQcH1zm0ILQXelGtNRGOd09QTWN+tp
lQf1KFcnmm3IVBAtRnSTncXJQhtdu7Yo1Xx0TnOnmE3/mtpv/5kg0F/9wXm+Rx/R
ZRUaRMNUTIKXaCeChOVA8jAC5+UPdf8F0qEybd9dPErrPkigDrXkDdddqm56aSlt
f167U9AxfotAK7KlhVJ0+edtv9FrEmkxjGzQk1p9gPf1L+KndnrO6LsB7JLmERng
DO675MOwBlDVtdh/H0JJwnOYMAJHx7jy9m1XKwT5YU7/br4ca1thqioDR8TPQeTa
Sfpl0cVmwLnzwo2vn4VuBwK0a1Xlp3DvUA0dmEzDk5mbtEWiZIUZVfjO+vy0qemF
aqwLZaZc8aq143/pKnKStpcuaju014uYUNg1BVo3YxpShOiaQCeRXQLGGvVP6Ry6
ArYdbsIJ9wKFAGBhzrM/WxtVl2Mfw+YMXR/+FG90Yvt2bYPHx7DGyFBiO4plITZF
159IKyTi0OoWn0X1O5Be51gzIotCtxUHrlBZsuo5v1oiEASwAqhNkLCWJP4yU4jJ
UnnpuOSGBGbjyr8k/1VuhbWSDjf8UuduStC1BMWKSaHE71cK3JCc7qLVGQ5sEF4S
28iTfDeirztn6bJ61m1myV8A2S7ztuLah+7WLLKJp6AT5tLYlUojT9TvmxVjnkgj
SyIs5GUUrfAOlc7LasgybLRdOEGcS+X9Ylht2wAduAXGGZdNKvlzAFHjX9N31/dL
aqHYmPLCs61o2jsO07OZAVdr6CXvWDCyn7oiNgkBBiVcIPkSOxiuNPm2WeYqGwNW
Q4V+ooPqH6ckKSwLTIeaQDEQXCb5shmE8xfWShwvr/1G0nB2kCm4laJRx/023Xp9
pTDjyjcz4gGf/M+G+cMa8Ww5biMhLMsMn98VL66H03ar92ElDHZDiB2y8y7RmaQT
thyD6uq/QIOz+q25L/w84Dv/VjNGF+3NVTM5oyOr1VRG1D8qW9eDdZThlZK8qV/f
x5OUA5IfJUqBN+qFQ4PUENVNjdCQ8m7d4O5A/8xhGBLp1D4NXeCqPS61btIl05kw
ZzszObFLqVoUFtcyrRjJ6F1YS5i7I2hJzkXgYLA3Tww13PTOnbWaL53YjDVcW7qw
1NKPuSvcUB9gO3v+7W1JFQX0dLCbAylN6upjxutLuNmBZTF+gis7mwvl6MD8fZwM
pEsIidRoOZ1F7/iKL4HnMBu2B4s4NgLd9ZYgtqOprz6JCznnh7pMlm2IvzUvVX52
wz/ky3ItUOJWM2SZ14s9LWRLT9bAeTP0pUO9OV1BPhZfAfG7FEXvM0g2uKZs1niX
lucDnvd91wwRSdBAGWHg/95mp7D4mOnC3ogyb+Jrks2Uuko85ZY43P9wE2dra7Kh
R9OopOM458+r4MH+7J7dnpFK1dGPWGxy4HNFIkPaP8kmzKp9LVpMIjQdEQUgCUKb
XEDuuAKhteC5GUDs2FPBT2L1yeiZ5uoSDRWYZisBWivIV4rm1nrWl2hjJQV7xmHL
DHf/h037eb4vV9obpnHcH6DkPBVBldvVNAKAuWX4kgyU+iUhjp0m8EYzuJInL5cf
lyRPxpTA5HLZJq3+w5vYpLHqEsnt6JpYr8aD/rTg5amJKXJBOB90FPujvaGN3bhv
aLLDC2CD+SkgjEFx+dZYhVONGX2M4+ec1BAkHx/hsLVAQvNy8Xuhc7LovyW44VQX
A2A11qOzPa3PemzRXE6ftPfB7tjS/HXrnwx6LAXYsAyGIWMieLK7IyUSTDHGSh10
mCJUk3uDGZQCam4YyUdvi8E7Fx5dfAEPVRe5izvvwhmCi8SgkHxOt/x+9T+TVO08
49leW/hQLLP3JID086qIlH17OsNKRhbLCeWK2+ncZrFt3OUAriT9GFGO0UcGcwRv
824D0fgsDIW3YALmCAgvRQC8PHwb4dimLv1AxLhwdXtjlAWQjexJFvisDL+dh/hu
UeGSouXPc1zFBjjE520tU0x7HQ8Rgyswl/k2iTj2KxG1To2HVRz0xW4I1vspun3n
kGPKyepOgSchmOIESGkAnkFkP2Ldu0wxZmc3E1Cje+VZorgfIUyrv7SzhExFGTTn
dExJ+lmFMOjsbWAusYz3Uqvl4oITFZ34YSAKtaNY/fepuTwrwii00S3pONBe+EYU
nzfVQTUeaKoIZfzPUdQ0k20yTIp6Erq4wVtZzgVEAAUZIENYLFNFGqSh9lLpQ3BY
rXmA4mYM73O4VrE4GWJ1g0slixZNhmyqAyolHlKnL8x3wl5i5zusHwy5mfPCeHGw
XVLKbMOMxhe5wyf5PqmCw4gg65SmbmyWuQfxc54RYn1sdQv3ZI7MY0tRHsS4B4gE
FjuyFq4WqWftbF6y+AECCkTNVYTUegRm+QXKX7/uXjw/i86DNVMFiVrhose1IzAs
FyGkJhs4Lb7P/H84pk69lASho7BwoCUpU/C5D5ikxlIT8X7+nG/33H9paQnZ2DAQ
NGAf1YiWJNJaH8xaf0BtlUfrQyzVfwMBLHlYqCkx8LpH+ZGQV4n8VZfjcDOFk+bw
uLs2qCJvbKSMLvb50lhRyaaMQcmtw7ID5DTJQ7MEFSCylJCJbuZu6vfyOKieS6f1
YDUlkZBbjpxNshRrXIOcRNBpJcZadTqC9aAzL2JHRIlPh+2e+mv26wD0PpBg66YY
hK7CFLGyldkpLZ95BQtBDiW3F8jG1zA8+YtRUdIF8NgQOR+ky37pH2PhA4/5rpYF
78MU29KqBp5X5O756+e1kKBteksYa+JbjUfgJ8PfjezeeZIPlRFkg+pd+6C+ar/X
9nwqGMGBrud3ICiDTR2Z1nYlnWB2/BTlgxuYpcGs7mfm1oo7IafSPYRoFYSeEjT5
EtD8aHSG/7Zi2Mx+PymRWeLm5PYuaEPbrcQik5GjP0jJePHNpTs0Gr8hYQIqRC46
I3mU3y9j3AfhB34GZTEnF+Jt6DjI1/qG4LWggvjYPIs6y4JCMQD20dKXQAsmyPb5
p1Cqg6XWqgky/60dciZ2UsLjAWhc6+Eio9w7yvDpMkP7EZs9EP85Gnaok3ozytAK
KJ3VhHdXQehQgJtB7vDbuGZh4xYTQUp+F9eBfSb3ZX1JPJwGbJBTlIOrM2JyYGCo
fOoJh9Z5j4ImkLu/F6wZRkb9k1j/mluni10FBXZ77lxUiOfQ+hVTuZy6RmfEX6/+
ijidN0TE3Kd3OPnBuQQ7/PRzCpiC9BdYdLNoFE/ZptMedrXBpavj84kxBAYHK4Vv
2MkEz3PLZT/FnfB1yRnpOtgna6t9zTGviB+wTVCPYKF3kx8N9VSHi2x26VimZmLt
i46w1/uMXcShc/9L1BXiXbarpI8ArY3SBxTBPpBcp9fSE80FxMTFLbhlsMPTq4a3
9dah6JmH4Z8q7C26eVgitPDsV1sLI7JU9s/XSkfq/jws1gWDXzl8m51iXnUSLh6e
K6MBKh7gwQxOB1zVHuQ0OswaqXVt6rBqegfq/592L4ks+q6O0hyxGfI/67cYz6Pa
P7LRL79KJCLPjIl6QFARkf0O4XOfnAA2Af7UZ1ilFplK7cC1oDCtgW2GbDiMKQWM
rX9GiWaGDVKG3nwq+W4ICejN9QXbaCThMrI3Hezt45BHDr3NFbsldjngUVMo5/Xn
yB6yu+PnBdO5MbQC2/HEUHiyfzPYpPYr7lPzvfeB2iHpFxjGMukgi3J6+eSi1Q4k
qvp+uSrIjVrUpboxVaFxOeuOLUP5n5dhnS6GkHokL4iJPAJr8mlEPo4g24QDjZp0
QiLUofPaWAqynjjKTTwAc7vE0D4hK9eklzJFv5qsG3w2rDaE6USFDKxRl9nd3nzs
YqImGwCQU27SmRPM5s0zhCJVzNEkSmGt8r6wqAOcevkVZB2mpxpHP4hmHtb9yGW1
LA/v3bauV17juOuo2DsmOwbbQqrsSXG6YyTJFvudcEpBDvtO1HdMpoDWYkSBGC21
iPGKpaZXWEJXTnbwQ9/EZZ0Ba5616e7C4erxDJ83ikkh/vk7zpb/2Qhd/eEea9Ou
5jifng1ZJPVIfHQ7ARZ4QJcwWuniCprhz2MdsSzOV7Us9DzW18ijI9OSZMwBdVcF
PNFplrxLPhR6s/cQ116PBU7dC9fkDegebPBs3WMp5gOB1X9pMrzXYnZ+Hkjgq+8x
rqYLCK881Cdp9eI3aI3er/3T34BxgkfzKv7o3xB+FAL83Mf0Tdr/XLstyHJhgFdu
suW3v77stIPuIsIb7GEVuRLnPcT3ETM86pKhz+10zg9Jht9K4Q3hK0KDXFI+Kr1H
sKRMYuOKM5jh7BRrLs8Nd/ieNjXmgn21E06AKl8OZYYBO7kL8vM76wgkNkgTB16g
EgA2HHeWxnuY9Sv85NCcdjZ8qsrW6KlrR2kBWO0QfjPReXdp2gqhiSwljS9TeKEL
7F1BEr5KCAIdBHmdAor1+L1QgJ7dVDqnjnxM0mX4KSAnIrJ6RuhozgrMvTDHjA8I
0pH4kSpSxyjkJ29FA4jvwaJ8rOKp/UV1fjxycBiAPmHfSmsfbTRPJ5W58iVgojPF
wixcltS2dj+4s3WUl6mgb7H+64+InxjfAL+dKsirKlyQ+36xwYTk0RCcNk8QeYMg
utqMwQJi159nAR1wb0gsT88wEPGIXu88lUz7JzhG5OhwMWp6l4QD/aJor8M5RPKa
8GoXZol1o2JHJu5pNtJ9vX6WeOOaMSYJKH3pkhx8BTgfru6KBeNyY7nE3GTXNZ2R
LDgjWXQ/TYJkboyG54fYIuPu/9y8mVxsBIxsRzP+v2pcPt65vtoaU5dmhEizqpsu
Ecn50M4FM0/k0M0/pGOO8WPiIVfs6pMMIaYCDRX/+w01MCcOtqN2QwpFoIivoCb8
62CN4HrkwnOEe2lOVG3Z3K8wcy7R2P2PSyPrTN2eQyMkojIfcYCyAq6zXKEptk8D
zQXBCMSYLo1FtGv4rc6HrOgtUHqd9GJniYUSoiaKU1iLiV+tqylyQxBdYfzFLHw1
1186kykPAMom2zoLMMwncQDoGurIm6NdwXQ1cGbRvmudouQrcapJYHi47B4jUCz8
fW8BST6RCVC55InByS/VW1/qf9h830+ZCsYBDrEK+M/AOCmVkie/liSiq+ejYCm6
flUlKK1aaQBm4VcsJVmf8YL3EC6FTI52V/F1WwNDp2qpgR4Hff/7Zoq5dAR0Bu0t
YTjE7z5JnjXLHRqZMOGx4xifAYECAl0XBAT0PyFwHygq86weBYZfd/IxbabsU/Yd
YisX/D9sFyq1hsdgzC9V0jzS6/6tsgwv/Igzzoz/Iro4WqBLiiG6LqCWydLtWIo6
gPFzHMY8spT7uhfMiF9p7U/yUKOaEiv3q2UQGGUh48Zi5DDYOTUxwFG4IUw6hC6A
6tez9kGiQht7RG0zp7IX2LRrjV6jQK1sellgGP16LCNJ7fHZ7142ilMZFiWKKUzl
kb0GTTbwwcxofXRUzadEwrZ8XLkkB4+oqliaUuzsy2UtrzKg6S2662DDNUlasn6j
cm6HrDDOmjd2xtMF76jflyG/7/11ebMR7FbjrnPXEf30YXmgxVq4Zvyfgvx4XZiy
klzvTprud0XpJ4lp6AxKOxeZaN8rfpdGO1/9WbBJfF7hCgtKCGgXXHro2rmOHjZc
2/HnomeTLgx5+C9qa8ZB5xlkrJMJRmLF2Em2PcJJhiu4nYvdh9DO1rMIjbm8wGVL
LBDfp+1dMiVoYiO+BMWulTxBShKCsGdbFZkmYHFQSyYh6JKczMP086TtIZs+QV3X
7Jb2N030rrkdi4SvfP7RwdShAdxeg+pO8b3z2JkyBMAXEX7QrMdeHEryoTHdViw3
XCFYy70goSZ2EQy8DZ/bQJeI9M8ohs/LCQvn3RSg3e3VrHR31gXtsP+4qHDs8H5d
0HmAYn7N/DJZwFSpUyn/KQxfEK1FOT60BpkKYl4Bdywh+Dz5Qj23xFKAPAgzQzVC
76c+n180Ew7FLfQT/rULeOm4OtOWWq2+WRPZTn9XxrMlXq+hkATg7NgNIyZF+bNN
tnYOiJcVoIhG9MM2YGQ55PXfb29ZggpCtvKJ8fYnuCduR45c8E3y41ygDSViERgd
srzXzjgjwnmnXAdLpGNUR35/+Vk4tGlZezk7Biqn5DnfCBtYIyDY4q4ZFQrhPcS2
xyEdziuvDKrzpG1mteyLFXCYMOvlAOLWIsL5ZFA66R2pwLZRtXOATcXrm44I/pu6
J6fqDwl4L16bpWlKDvAe8DvuXfWHFbBTPp0JvANNk6NvsjOh9whQWUYgKkuKc8qk
KsBMVgQc9CXkiF51G3T41AcTU/XdaoleEnB8MUwlpcqgPAsB4m9fnqTcBk2nHywh
/Kw9/GMSHgZRTqXFUdVwMlYY3uJ1V7gBZVW82NbEMTJ6W74jZe6ilkYTcRCjAqcc
OGD1uVikb7PilODlmLtCjmNGKao909E+Bcf6UJ08rnHiz+yHvekIja5ztDjd2ulW
jcPT7GH2yNXtBZI+jKYajIZ5Zw0viVUAOaEHgXvtFgCW6U3auX3s+kg/OMMJE+CW
hIVWaqEpD1qztSNE+HnZHCW4zqlnx0H0JmMs9f+TcUN1ovSotMz7Ol+GNc743VS0
deW0YsvTRP5neKeXn7OkOswAlGJ0nTAklKuYpcni2sofWAYN+5Xul1jwzkgBFVjt
h9Jlbi+wYWrz+6PqmlEX+jWAA87L2NtxEqv226SXMddHI91YhxLwWSgvQ/tCSt8J
NTGeP64kjirS+yJXfsMNDtn2ARxcDxi25c0Rb01oXeLFzwnqR6fb7TV1a2g2y/IZ
9GL72xJo4PGu42LzxZdq3l3GGfkBaE9izgYJZaaJuLMHiWZr4PVEUcdbRZ/JwlpU
cuuk1gK/NiuWtcfEh47Kp8fP0oKODEmtIHFLA1TiqlEyG/dSTr0s1csGUJZo3M4A
FnPubU9y7gtRP9mP2DOUeZSytattGR23W5rJ4SDnlrqEIgT9YVFNODKo+jypyfRq
UWoz0jSa8meBOzB1hi0boRC3LdNNkjjjrdDdOFfl45k59Bu8045OO9B5UyohxXFH
ODxcQbC6TM2wxxPUtBBK8cCTr2eVfXYhdFL2WIuwBichk0kREFt35U+xkRSLK6V/
+K8B7fYj8ZSrsD9nOYrrbuqDUzao79eBHa9wt65QmjcH4/NL00NY49aNZAQ0IiAs
0P0LW84SWSV8JXzQPSTEFdGx28YbIigYj7W3E2+irKlPC9RXH3yPRwf/JMfZjAnZ
FrtAYh5bX4JPYsLrbC8jA+1045WlL0Ktd6Dtv1jE67svL4NVjFJ/CUHDLu2wAqtl
8QO6q0bG099NcwYG5CS41wPEwQ14YPJFQoD4vpNWXhSQnFSUMJOJiVeAHCMIoEC3
zUaLCXyvoR0qS+1MyqIppAlRrYcCLuukUgBIKoY8MaxWXCA6pb/a9h2Fijts+LR+
gVmB+6KvIOk83OlWT/n9JPsXqBZvL4cONQymADu1lgzC8+pIYrSMLEE40DcDKRBk
FjyMfXc2p7jr4OAAarLg1T89Jkus7AGBggGa4+/5GAk/6J5ak65EfHRcSfusRDeI
M3+CGXnW1Amk2T1GJuEJl/vfnXQveoHnmuS3orePOte2VQIXzNA2594fq+iDAihL
NCDAK8Ue8Hav5ntImngzC98rJfEG2X2su2aA1QuwCx16CPUyzwg6SAvitVpUFfNF
RtzKYXlNKqohrDioU0xTugATstrvqBDKPm6PtU/zG0a1VBdwWiPFg88nKEoV4H1F
Ik/IloFWJDNM38k2ju9cSe+PwQkxJbijoNO5RJCR2u6HuECdeKsJLDg/KQtpfZWE
a2eEALYKtbYarm9ou+bNVp9J/4QG6tr+PjlZkuxBaxkKGiiXJB1waTJU7jbVs69O
/hioajKW+V0pJKFelgoQ4nSBAavphs5LepjT4NwuMja6+FRucWUQHblgLL2AWp8u
WtULwD90KpndwF6C2zhUBxWUdx5nH453t5LeBQqFys/fb6auiqbfN0NSC7q2kccH
ZnaGC8n+iaSfVSNrkQK4Y+LybP+DDzeUPh3WK+CYlqB9Sc9wbCcdSAwP9CWsk7pJ
ZT5Y2ht6hsQC/MMCBREUNuhj5XAh+eNQT/0ekvoZEF/nu7biSRVz2a9rvmk70NnR
igfa4zenU06mKCVmK/2MgLM2OItmJehrzsBYr6f1Olg7+7se4w2u6mWsPXqTzU8o
xm+q9zhWR/uCSN7bD66ShB3z4XewNJ3oC2xcCSgm9EsW/Uud/QS5O/fzIPqd9eD+
H4bY49XR1GZJEMrCpy164/OYSLepQdkw67L4043Ithi15boPPhsZBt7Dfw9cadkP
LcjQlkCJVibeIu3jnE5MMoBdrIDS8jIPRsNN2PM1O67IqQ8ohXj2bUbHFUYBsYPh
dQWc5vBIVtyyAfVbKWTxvZN3garH+BcD+fa4H+nwpW/oaMe3A5cfXyfc/Vv5GX1L
cAqxxeo2R0zbIlDe2mgaQylnVMu94kKSF0uVDDUXWLef9DmMDJq6bec7BZ9YfcEF
Tv8nxqqIOO0DjifGQscpO+CUXooUe9WAgXlU6d6gthLSTqEnkbop5xDVqG61l0ho
2q3Ekbta3LCwyoA7q+2YZLt8ZJ2YrJTLHqA7SOM8kuSHByz1lZu5xeUR5ePtdKRh
Enkfd2IGcIIEJLtYX9vpkk86bXdekZdHC3EKmlFO6bTYaePoumsVhmFGcTMebpyU
HBlfZp3jY/PFZi6KYOWthSgRxQjKz6aS7R9eH8AWNTvZxpE5xJ/a4gJ0wTYElCkK
Gkiu73iD+duINhREGP5cgta9thQ9A/EAwvf54fjXx4GQFr2Ob8VrjhZUsEKdcoe3
/kgtHTe6bLUYKJTDlglapa0bZJi81IrePY7Huci4Z8TBRXIClgvaStACVzZFNczN
MDz+uYXLUjJ+BHFWxe3i55TsSjprnHWDv06iZyi+65R5QAM79sXJSLDqt1f6Ne0W
Rl2j4/SEi5PiI1VfLMoCFyf5VkqBHggdjqc3qPPdIUABklwNpzQTYrmiI9JkAL2J
mwKAgvvwRVJhtW8huCnr/qwPcsIOjCVZ4pC/9528blryypynZI8hpChj1f+CBhBJ
/GivL9xP5kZRW9kICF5cLn07o9VG9m4lZ0rY1q+FSCwzanWDv6xUSD+OtFRazaz9
53vI2Wdnaxd8L+bMGSn2uUT9DJOjeYfV/C8xoSx/I8w5k9Za80Z4mYaYl4gGLHwD
q8aEcZ5Kb7X6+GzUh6FMTFbslgSpN0ps0GCGQlnk4zYEKZIWkByQ9Y4Gb4RPoaOB
SgESe1XNLFqDN5p/Wi4fZM9ze6t6c9bzChRdZuZxlqKKX6NqT6KmsaUn96MjN/Ce
qBWf4aiVGlzfhuyfbP609ghuC6KKjL+iwot5HKVnujIKr9t5TzfsTYFM6Oxo4fAl
3Zc1rKLOikVjKuiLRVR0POzWKfECqCs7Q0y4penQbrXVErvbvSqnZunaNdEzfCAN
+oblig3dPMPifIzpVPcUXf33dkFvLH2lqL570Jvo6eYjfgaYLf+yCwIASscpajLv
BelXCySJdiq7AxEzDSUzyLXt3BDMbPyk5+xdIcUjavM13jglnXByON1w10/6RwOe
oiC5ukhUdwVcOAqn5rhiiKF8/iyJ/EOOluCajnyhMi4t5mlWNIChkTBs7ZpC4oL4
gTQqTS/DrIB7pjUuXKzH1kLvNX52NMHy+D1JmCpBNuWN5zIEpx11hj5rChMx0oIc
kGOLMdxmKtp0181NOVg8/f8VoJ1wT1f+b80cJaalKFbse650YFX209yEOcL0c2YY
Dxi8uFkTgbjy3LbPjhwCbML50daj8pEJcIsq7hw6e8wbaWWfA4Oo6gbew/SstgJh
EgahqqrMbuEThu61Sd8IjB/A4LN94njfdjmAYsNSGwY6pZLP/pb+jmvhYOHORcXP
6RUSdhERznRZwI8nMX7QMxwQrqmCCcato0/Gx/NBJMgLTxgvLm08L77/8Mwg8vgj
ZTB/yRr+6pLy8lQ+z/GUtSbLlL//DM1QDlkO8BJxo3JHNqINHXO6gDyvyT31UIa8
mhNZQUDh/DYoT33OCMDAiBiZAk6XtwEj8iovLz45dM4s0ANdSIP8dp9WOjx/Y1zg
hpgLGbUScQ8ZVVZfHAKzKNAkmZ3e1+zRi5QU6wR0+/0+2Inn/yEOh9ps4l6PxbDO
gYecyGV36Zz1gRnI4JA4dpuEL8R/I1OWdQ2LkEwNLDCs1LrKky1Wf5H0rMJP0xTX
rwWhKVrA41/Hyij7n9Q3tZPLi7kLWyzd+P7m0lXSPYxf+tqz2843HS+7qa2GMcwu
Jv3BOa7mSPk9xI/1DSGdCOUde+pJ52avpOC5BvOdDnD7avCSOhI3SsqTgnQircYZ
mXWj04kSH1jKjvKQJvNBn9sE1kUuMiL2yReFr9Hpf1IeziexsJRuCB2TaSPS6zgp
EmTy8PncQ7PGsWewrf1W2VWtMh16OcBTy+uD5Mso9TXpFiQ8TlcnhOdyd1N12sUE
OjcXmU0b6A07hyhQ7w5z7MBOL7vo/OyZSEfeSiIQS6ehUPY3a3mQQYawB2AQ7PzV
M9CbjEkYFFnGxUlIzOsoypEbwuXfmbNrEnYjpjPo3eWwbLK2yDwUmL9iGzdFB+kK
fcST18OQU6tGIV2G2dDVlz0HJ3rQnEswr4n+OF/os/hDH0d2taLK/gL2xrHFrmPQ
b+6uKU+lIuJ61ldVIF1TwDSL+MvoCvqbP8qm1xGqQFZ7UkbA9U3GLlmJYNvhP45z
sHAtHl/xBiqyh+Qn5R2dZaqk8Y6gOz1tagfGLv0dglIHx7HDgKqWTs1YGVXOAkL3
kpnwCiX6wy5rOU5zunK48MY/ObQTlhjXn7PzLayKg5XObHpr3BabgpkFe4J1M5dv
TWvn9i116CKYuS0dqiwaiNd46mP+K/N/5w6T0fYHo/m5lj5lhiRZSlkQrpPGZboC
BfrsR/bJi1FAPQIJzPm4QKouiW6d7LwQN1ewx9m9GQFWMMrU6bWv58R8vaPJ3/EQ
UlzknU4k1+vuTXaSjp+bZ6QXEiDHZvR9l9L50MrMPQZuRmvE13gr5/KphGn929DQ
ySu8FEti2OH/n7b7334Og2JXg8HjsZMQYD31HX1LhNmN3WOdVVQlobNJ2ztazSf9
42Ms0kz+X3H4dTLj9dNnmziwoS9iVVA6oDHoPQxqwvQ2QBB8d330r+NxZDtqIsHE
GEX+cPeN+h0tghnA8Vc7Nli/cJvMsZ0pdvNDrQoBayj+HbuAUzlNFq6lsLuHy0Td
EMSXBm4u0p5/ZKzayW382YJefazh9JK/LcmXbjPhx8uSsCZ/HHoO28q7i1p57sEA
hh6C7Qx/v4jdXbCJRw6q7lQLtXzT+fHVEiEty+Fb5H4IakZ7tFNwAH1h3uLpEKwC
F7+l1L0rwHghihFudmFSAfySCo+nVWKGUtx/Y5ONyqMIO1yVMWsHRF/MCb0wiY/g
w2cPsQ5uHmgj2B3g8jUd4teeUPdWm9khwnc9Dwup6lXAQhOSblIJdDN1nu2rEZGX
m1p4USyuTQ0DB4TgiAsej4jxqYza8uPn2I1KMAhcvdEtLhVz3VpZWRSZjBOTREqS
AMsiAQvh/x+mLGIgUcs6vToKQqmS+kEtbVvhC6aHILrz+crmTghcWVbqlTy+VfqM
mqDjR3smmn5/16O6g8YlNAt9rmI7nkUw1rfSsjJ5ga9BBKdtcpGzhWFRMKTVFaHm
7Zgf7FWUml8IvjUfyt5i33RObkeK0wKEUSv3dZY6PNUI3hiZ0BsVvwbzEOalyeSE
Eb1ly9CTcWDre7oP3lTbyhlITGQ53LDMvlYPgNf7ErqqHsK740hto7cymct+p2dD
hnImUHL5BU8cRb2bkTfJn4x4E5YB1G78iNQBnaBh1bGChqUswoXvsUGJSAeyFxcY
TTvb8X2H7V247oUoMr4NVUSnElDt2Vn5hGbnJf7/PziSF3MNwCW3RoE3aLNibG1C
sqrWBMAxtIIa78x1L2gA6y2QuibUh6KVQpVSlfy7d7z7mlcpz+IOnYXkOUP208n0
xYi2oxj6pheOhWQYt14G5CmNAo7VuxaUZD62AlMxrErdr3GWo287x9U1dR1jYj+w
ZsW6ugGKgsU/hfRzdvsCZi8TpYa2BHMjRxrt4AZvqht2L4Bp6Zi8JBJ0kUAHuo28
UupY2Ygjd+iO9husPGuv2AaxrLjUs5cxCvorOi+9aJn7/Qt77iZAHVG3M5lu/GBK
oxB9eZi131BKq3EMDOKNduKpucmn02nJLKBNpjMHLCuuDhneTVMk7+N/o6WQ6Ujm
PRFZ1a5+mBMNzLpNOj312N+eZYa49JlWaUEUEF0WGz8kIlnRPlyAVB+lrlylySJ8
j5nRMDPiAx2U8DjeVpfuMezEJyYBHy0KB2iqSrmFdHghb82O5MAx6/C/C/vYOHM2
qAsWQhr5pO0FpEJuMGhJjuj0SxbQyTK/AG3pTZWYHeyeg2vninB2FKWnjLbRpfT+
qFz0Vp8tTFoDINwtq5gFFOIZIn4EheNdpv7nfT6V2YyuAjroUws7kDYordb1/BKe
9ZYceSPsOc7ComTmDHc4RnUrQoWdlAnqO/6yOnE/7AhBkpqAWqDHoFEz9d9TP7vt
fZgDHXDO6vj+x5ALj5UMyf95JdKDpzMYlz5Ry32MHn+Kk+7EqJTTHpMDtCU803KK
Q3isqgLd6M2qmvWp6KLeja68QAealZHLKDyJf0h2quRvDojZSRGmYTLgyUZH8Q/q
wNM00yGH7hdxzSkm449KMW/Jj0Sj+ReaaqlgwpIMk8ULOEKGQhhN6EXZBhNcadbw
2TeFuTvYx0P56JxnUt4aJfynL7boAKMzxMIC6/hCNL0x1lkkTMD/i3kNJA4fucdi
uY2nHmpcQ92T59HJJE9IC9vdEiFkIWTxRlF8YLNAng0iq01uhz21LUH4qN5Za+4a
ABuTMepfWIVihQ+MPZxBrGPkcdkERkmKY9EUsnEVyk17u9btSKaa4ITDqNfz3yYS
zk4gECNJmfuVyK/WzeNfqVCVX3NhGOUpiOqaaUkDY7Abw+9ax4ZTqhZOoRBrjohZ
5xEooGcNLk9q8wiqCM7aHO92p4V7Efg4o886KvlzeVGSr7nmU1hqm+qzJa0YHnal
FL2tnxobazUl8CREarte0Phbmy+nh+kihSVeziNYCeNlwC+RwEIUKjPp/dVAZAIB
xp5Pb6pwRu0qLnz4Nj4aZIWWBMlj6RoZQ8TodQGfnQBVVTxXka4OVqDZL463jIXK
QOeacwIUf8N8n6GKCheEOlKp+q7ucKwLYiOvLl6WWh4qCNhc68ihcHno93s6zJmq
eucOiACpXhLI+TQ4+N718QA8PFXt/fMGmLhoe1Qbu2//pq7Qq9kHu1XkpP0AfcUz
T+JFbL0qkrXQwwVE1UUv8Q3YnsE8FnVUbT6dBFBfKFvK/DxWV3Nh7L0q3bMErTgQ
fJ0BEgtwiXkXzE6KdiH3dzDtGfWJtUXevtldx4SafZNshQ+WqRo2104MmyVLPQle
udnfWNaV4Xum69enZS2XPgMCzlY4D4Y67huKpoDk3k5xibba6ru6L69pekmZ3/af
+QSJltwEqt81/iGa/QxlKJJVHZocYi/GMmHY+mL+XR9jWFjiYAhjr1J/aLq9rKh+
3uWoTVEtdQz0JfxrN73WWCR6jvp7/xNk+JEMR9L6E6mi53rwl6JDDQeTl+plIT1A
sUaFgzYeG9s1ccHRpoVW45S9SOQpzA+A9epSR6AbdCDEwI7WjGwSjHglUq9eGqWo
yTljkZdOZpiDZnZ8noQ5YiODSTT/7b1B6g5L8fu2ZuGgJLhP9/WIflGVuT/eWy3p
Os6pEzYmO3aIXYqZNopB8UhxDWqAIhzcQ8qKPYmYbkBpscuu/2tjOTxGZzRSlQI/
s1YK33m0goXTV/kiIe1tKcQRs0/OB/o6q2Wae9kqitxp9XZ8+Td6eBW7fnOJ40+z
DUODruEQ4dw1nr5nony2Ut0KrJw6QZb1ILyjE+mm1EXYVTclvuhH3ZyAKfwWQiYE
tZhaDKIx9W4SUyru4be3PzTxcSAzmLNRmCU75tfCLPYjAt0V/rMYlnn7GNG/NjZL
aSwXXJTlYYwDCjSPsrr484SG84OswCJhlcfJffAt+eHpHyL51FnebIcN82gv0bZx
tpAhQs4YKx54dzqt0ME+Oa1SvxdhERDADlLuEN/Wby4/De92H1CZmpUpri26hOZk
7Tsv/vXmAwNd9CdVgpxFBXmdlfyWJqhPXFStxzTQmunEUmVeM61cIUZklJtOJEqu
1PQxIVXRtvFvb6hvWpsSSHM8B3+ThROCDzRxNoUkVgTVRghnsU7tjbN/3PIPiEUR
poxSUjGv9OdKXdMlkkYnuiXbMBNF4sJ5ehrFOQzRBesoYN10BNXFLg/DwhVkXsSm
XYU/ZOWHj26NmIFTBx5jSGVciZZLUFYL4fCm30IRokx4zY96JNoIdSkqjUSQxLR1
xMr422sBunIwirUjSjFStkqYebVBOkwfjM8X/9Jnn4Pc5DBABLDGxHNJGqKwqdtU
LWhlE3JAIo4G3G5aBB73KNCJs3nF5TeNT1C0LWAkBTAG+/DKT/KftYWU9fxVE2xs
Kqqpht3J+5Cb9x9dxgZTxqwDksZsmpQlAyPdsjaRg3xWmiecKQCCTV1HSxfdej/n
vBDOAT0i2jdKlNzC1//l9f2lM+DKpKD/W+kz3FhASAFUbH8HO5JmaIkZRK+In2M/
gDk2EIWYv/dexF0fE0RuLAq8oQm4uzN4VitEgDp1m+sEpqazVhJW3QGyzmPQMPm6
aXJH/ARzjsU94RBiDOJkVVC10zWeV3N/T3jtPoUGAOaxVT4wRNArSD4hjy/kVtzt
GoGIaccd5irN2nK4T/VsNTHyj5woeoW7cD9wixOD93DfakCdNpCPA7VrjjaalqA8
TZOTORjBks280ol8eVuIwe3u47+adqm9mgxzHtrnGgkn1kd6PAQKS2qgrCv/40Pk
eZqGCT8+8wx98rQY5HvyNnyNzcYhG8J7o9GYPPSHLesCYwfiQ4kJTV/tMf6wYZbI
DziY0XjCClga8KDwIQsYyZ/wjrPohA1bBhjqrci7IiSUxz4sxE3ePtFS8RnRMkxU
MV9L5PADviPWrSuIn3Y/6S4MhHmDLuQjDwgeRasqgzNHAe55x1WhTDSIphKONAJQ
zPiY2C2RPYlMzGxdWFQwJ9vhUVTy8wgiEbAz4W6pzNwLl/89Vv9w/sjbL/YY7wKO
xdO9wEYzkswU8H/l8ekZy/O+obpVRgl6p5UsnmsLs3J0IQbbk4rszdCEoy6HdbfZ
nBOD+HQPE8EJrxr1pxz9x5H1B4yJxmcer2aKoerUVKdT+D8qz0B/gz3wd505MdnO
kjkxtarHmPUHerU6zvXKfNl9FepU3qDbxcIMFvBmfNCRvQ7sccIaheOjczqddvFF
rCtFbFs5cBUpd+MyLSL/0TMugTZFqavEJGrZNP781kJ6SCujF8pI2XLXaQg29fYW
/trMvDzg1dLEY3Dyr8J9PCLs1pjVJwRaxgX/q3quDAd0sJmp+Y1SKWCrHPXoNuSR
aXZMr2myfUYLT8PQ3pExR7CXdrmnsonBI5NCtsku/+UDWeG9wHCvssmA0F+ck12T
XSTOh34mfoVrffA/9PvK/u64ILWoxaj4p/GE0EGUX7pNJmSHbOOgy0OpRet5WDe+
n5promC/6Zj7K8H/RkZLpKHDo0yfhLztwDBfZdi8afQpV/u/zWwABMz4Oc3fKrG1
zwHLcKNcIoqQTKLGwp3x7207QQRiR6hvT4TmyU9o/dPvFdgvS3TWJvLHDql3zue4
Yh6POFvgpZWwprhT/CmxERNWCEySxYC8gc0amxHiPNQdAvqYzh/fMTv/BmJVQ3TX
dvsilyymRps6QJuqkqWQ0DXhCPcUlzs+QcB05GOC+h2n21n1KnWfha4Wi+oVZ1cZ
5FUjf1AcTHCvyAiyhtvdLTdbYtNxnZ6cd7TkJpCFjgvLaSfScrnX0fKC9fHuF+Mz
/pnJ8hDqiEL9EAmp+eGfNXNyBOqYyDw0NvNaF0kfBFyBiubS0YWpfCAugOadmITL
y1pvZVpPhSNrLMgj+hM0TUdPpdBdfcKSFlsgO0BLpjXj/l5UBf2OS8xSL1Abwzpl
l10OiU+vL89lhhNk1bchniJZAFtrNaDa3fUBXfRqk3uTEqPt36J+Qo7lfmAV59rW
0M0UPHWjUWysIbkGifp4iTpomPw8KdEteEpH1RnXWliq7Y236gMFtz6mJt7F3mS1
aFS4mLZ1alM4MTbMmLxM0/ocXvRKTUN8X6zfxlW7UOMMJHKTjh5tuRy6ZXI4OrAB
MR92+yPGnpKauVP7fcQafh2Y8PkDKeaJnFUYEGKM2tp67p+lbAPzVSr+/ZVoR9xs
81dWmcrmQkVDkTo8Knp6ZqkxB6/kPIcjdPwXKOm0ED87erFllBEPkWk3ZxfluHve
y80TNfdiJfUUOagohK1bQZCQrtfxtuz4/h1AkAyxZZcANE9voU47VoHADGqyOPUp
napBWzQCbuBHK1qQAN65Nt9ReQPxE2ghozAIceIXJ6EULsSMZNdbZNorK2OKUb6n
vt5SrebQSM++bk7i/tXgBxKBbgX+1xMjVq3+ySvkd+0Zqe/nsH3xw6gIuujBzmC5
D0k0CoMkM3tww/11DXsLMTnPgjQAw/17XneQ0OCXABtw3sQqkVwtWc6Wnxtqflce
l0kd7Cv8emIvg+1NtIkGNQd2yK8MO20/4oxqrBbHxF1iAHpTRWZNrFtPHys4ZXZP
X1t5xkjWoCLAjqX/rAX21ssc6+05eZsUEN0pxkzmUPPAZ2I6JCNUAuAcT/hr9mGl
vyE9XQTsmdIQG0wTrvDFfXAi4arGvsuHy7Q34/24tqZKejjAp8Hg0JCfdVlhxzkM
K0gzxw19eeZUH3LSHbB3BG4nY8jLpC09Hs8WJ8C15iIDZVwys9n8jP/gPkuYpwSj
Ou8k4sPenjwsIlqor84/XJUhvupHOhaczuep0QUWqoGgNnS6Th1t38vIEgO5DoSq
PWD05vjQqwM52wGm55AJ3J8bPZV8sYaZM2A/9Rs8UD/JEPxHDAFtXrx9WVpFKJKQ
IJUXiS5xlFoTHaYjLd0UwsqCiZ6HiUT16p3QrzGGY7zSWyJ0ez4XNheBTuijyXUC
suQ2Jlrz9ZM5Oo0zBbLs+o4EnKgSUB4fzbp3W+pYSo3eGmIs42LjYbKnS4SxWivP
T2Wl3R1eOREkT6k8YZFBoHg8QJo8ixlfDVbwUGI7aio93gMrZFzjxwUhnnZmWdiB
OTkTckhxEN3LOI58ZlGTimLn7av01lNwLxwt3UWYyc6agb5ITV/aLNfKe8O3NzIW
sEzUW4Nsq3PRV3iXFWX0p0z7PLxQfdpy/pZ/n4zoOIhgzfDjCSA+5gqD8kw1/vxD
FC18eEcGR6JuxvcIB42XhqpBgWt6109TD3f79mQkSm8WIY4NGwmDWA1TCJJS/uvn
pKSQiKyYAIQqnhVvt0/jmieZ6z84mpj4Ypp6y7AmRZBrgWBZK9t2c2UgVoaZBkAp
ToNbjdGB+01SSHSsz/snF7z2eUREZsl8qdHC9UOHO1YJhG4sxudSb+M00Z4RX6YT
kKf5kBfqeiYSfMKvQoLtgrvfl6UvTq/dRMUdScds04eSw8JgXeh+AoHgWQ0sApX5
8OE9kgcqqvdB87FxXRhYZmLX9XOJ6pRi41fbcD3CaZWi3CT5yaOUVDFsPxfiJBbz
lMGNAyMSUdYhVDFBolGGKOOsOb6K+HQk6oaiZc0fuI4NV0oEkL8JBOx9PNjSnjOy
vPtq4yuLt55TSRIJ4VpCMqk5jKTuL4MGg2UVP0/kLIViFlSV+SDLUP7rNscOLCq5
ATPQO5U+eEakw1bHsrVoADVKaL6C9R9Df+EwxCdligOSD08vvgdvnli7RXZSGtCl
UH8nKyqCcoLAUUE7GhBHoLEJ9Ra5Cisli5W48tO/xKGb9tewD4IammqhM022+LD3
+g2hq+ai1EW+XLkzuTscz9jNsiDyhyOUSpI8u9sQ55XoZSobwi6ofn2cMudp8p1g
nuOAtAN7SKtTGqskihFFAo/yf0xiTt/nG0e7ZEz211CcsFGEJjTG4TpYkRvmcYtU
erTDRM2ZH5sOwCXyqIr/u91Nsd+TjHQoQl58kNQVs5xDQKNtDUK2zTeE9ZkBpQF2
R1QbtByVnrRB3DJ3c07mkhaT7IajBO2oa0W8ia1yHBIeMqwcWYp3RpMK9t1OyoVO
AhulJ4wU6Mb6AIH2SFk3RIVUOentTUUocFHPoQh9rUMQ1QzlBPU4VfRd0aU4OQ8e
DY7i3l7mUdnqVfVEXXaY1L5f6rwb7K2TQ51q0uYS3Lkibv75p0beToYevuSFnKG+
o28KlwZte1BjTSywcB/nL+mGK+oa0aMF187R+wn8N3AFd48YfOxpaxMx5tOqVZbh
I8jEPKZqboXIw9fli01o8TWBr5hY7Ma4MRi1WHhk6v+sxX/4WMcukdfuHigZZ3Am
j4rSfpyOlHUPaxk0cLVaJC9VKOalSAVSgMiOEMqSQtGMqCoOFcid5NS6MWHM/SG/
e50yWJk2oQHkGZ7eKhsrtEHQKudbX6JUDqS+0bLnnljK5jtDq84DUfDUa//n7gSK
rTt48QuuNCU16EyHncqKpSBOgFukUOsY0WWzuOdW8G/L/0l45t/OcqX9ULiQw5Px
62wUCB7gz9RDSJfsYf6I0EpSVut2FB9t3WGfI+VBAcF7LXTQd5tnhE26eci86ESr
Nw3yN9+q1ThW9H2FzyfUF7tOZq2Fnq8L6Xidq5DpAAKc/eBbBnIP1nv5aeyeuEaV
GmNSaKHRDF4bNEy3orR75oNsyxD1e0VyzEZswUVnWzqV3WQcjsYnyS6a5Fp+jwal
F9Fnk7hMivJ78febS9Z05xAku6VZXGeg+DZ8P4+FFdzCb1x+CHcpoJs6bchhTeTS
sJtHGGEK3DmvthHdXgzgyLi9axhvAeItS1B9Xc0J5ZJkAzmkVZJhgFbBvyYoatiS
ajuq5s58MtfekXqAuSRSAAad2hCKaNhoyRM0vXTw0r4k67CtFniuKd5SotQLUDQJ
MHan7BbQk1PxDZWs+vEU04RHV+nQJHMBlweI6rabvJQp6uRUWr/+eNPhT5US/XEZ
6pyUR2gTPpxBDBeSgqEYa/tamitDbA3I+p3bbHcbNH+cIcNLerxEGWqbtlYjRaXe
YZhH2v4v6IP73ckCTSXKR6RaQeg4LpAdOYYicWhgrwVgmYw81EbJS3UDI+0ppHy8
/BuMNZdYW6pdzCSoJ4SXCG8yUuKQjBBOiokbyPdc4dd3AI8JsoIXyEb+5kttP+zw
XrxAg1xGgAvx/YSCVZYk6FWvkEKIf+zH+h3rbsZo5im7XHRtorPZipUExxc3hoJA
bGGX8L2LXtkOgA5PXBG+rJ7HFdeHcm+QLXRXB5GnjrA+K0iGcVtr4HnXyDVO4uLN
CliBNeK2pyiWLFT9E40qFwDWYaMcAAZyGhykCQkBnzLIOfqmWMsNczc4DmibVKH3
nACKGjVmycSKINGQn3lWLtWqTZWVDy2WoYkHf/H7+eyv/zAAmff2mpJKOy7oDLEX
O+SUwreRGmJbZtVKYDtCeyHjbYZQHEfSyOhGt9/KzpqaQAArtK5tV1mqY5z3fJlM
qaLN/uwKZWRU6cqNz8P7Rh9G8+0Oh/WI0L0sXkQ86Li8muC70Cdo2tftDwCU4DXS
X2HAFHtCMmQa2MMrKdYFwIidM3h9Lh4yUPT0ok4kSLztl+DT4O+LtLoAFlo9Td8R
bQfpQiUek3V5emi8HrjjyygMFBJBD3QzXiSvLyBLFG1LML2CAC9coeJmXIgd+Wqj
2195pxzejQuIc6zMo/G8wjIOCpGIWaNLW1vA9A9s4cUnSQU+LoZPQtCIO/BLVdpW
qIE0EsJHaBrROb1C8EyYXbA6QCwCpuHSpJndqyE3sDZgB6ZgFsvgrFip46WSX/Q/
Eq3tO+tDRqbUjrcMuiE0MvDwUK52K+jxWLYR3iIyqhuqbBrDsa+BZ2YyP7aBFVqL
XLJKRcIVLV0wYSenrJzWGNJzwzzi77a/+8dAGwUiw8miT1qa7r+/Jv9+9z2PGXuD
cGmY36bAWW4j9YxhXqZUr3a9u/4FZVOC0Iu9Dx/drrxijwCeIcMKnsRFbXGS48ml
DnY4wz3GeKgNraUlH0bzIAr26bmtP+X1ww1IWoiccqarvq0HvLOJKAW0KWBgGooT
wJgW53dNcTlreWl1u+dtZDlZQU+0aPdafd6HFnYRir0yGtP6T3G35tmpkYc90e8u
4LjNgDHR54aZAhUP/j6rECOQ9jkOwAdM6ISrYEITzVHQ/CEUQoTDski0qka28Mra
7OrpW6B+wAxHfS4wnmyU/h+HvMqM3sgPErPjL/h5EmaX5X0U1vMRVRRvxiy8MRnP
09W5C16QJANpXkzPs0CBEvqGx2cIr3AO7OYHhM9hIiptMJxBwTVJn8g9ZiP4MuY9
TxOTYC7XrO1SzLDwgV+KyGzXr6br8rTKZ7Ib7wu6VvnrHWDpN339t80K+qLP26F7
/qhtZdwzTUhIn1XineMf560mtgxJmfQXv4Ae06r4EX6neT2k5Y/sddz9YXwwruQo
91BV9195FfaQoKl5kOnqpxSWJkuuQqZ1sCma1IpQ+QNKRYISYOhWn3kiE8ydIrQ9
VHvnUNkVjGP4m3BBdq4hVgM2n+Pg4CsTM+HGE60+nRUnV8ZwbVU9kGHRapuvS04R
eqKAlRUFtnRJjFF3rU9KjygbIg0YkS8/DBC8tNlXCg3M6x0/jrwvOaGUBpWu6cbv
AoFms5cZeuC4mvob3TdGiKwaLU7ef0420LZ2nmcn6u4VgiLx8laeDvDR95wBQ4SE
BrYIWg6m9Vr/r7JG9itG8+apfaeoAqlR8jfieiHGMTliqD354pn++25gX1n5/DHl
n6F0f1L4q74lfVPcYK5v0WLJyFGYwHOWFl0j+JW9aaPXZgqSkttNU0yYRPa073Jg
Wx5eV40FN4fsulF1pir0Ex4sUrNxjMgIYkZx0D9wr5+A2I9MBRg43HUcrM+8v818
c7FDcHsh8hvF8VN6mK5l8ldpxxXNmcF1VVaFXOPbbzD+cTdnlDCZ5+xyS9Bvh38x
btHXpdCDn6InVSdPSGwUDF19MVTVXY2uJ6sZV4pJOCNMyx/RwCm/iEp5upI5DtKL
D7B9Hb6vT8bKcgi6WddNf7visvW9ClBVx4ebvDgHmKV3pcZBn4GBLP1jO6Y9xkxe
nnZ4tY4ILBEZhGZLskxe+lX1AKjeMFomlpkRHONY8TVaNMRwUD10WIQZall6xMca
Z1ypbdbTclL2XwZUSzGPpdz8a6di6Vt2bCz+tI8ZjwCA18dJ15PEVH9/7WsleP4r
8Qt7nslv7M428bISA0cWKuqTmt1p+lyH1vK4/3ocaWrXz84Ws9fXkVws7c1Zi7Pb
dFTViORhJ8PvAdfN29NQTznfSpnIsPzANq7bcvJlIE3bX9jQiXdVkoIXfqpPOQPD
wvdqBxKBufC0eGLXubRnNYJuKoHiqUtAYNuI7XvfHav40sFDi9ytXUZM2klLEXQ+
cqzi/sdsq6LiaeC8WtkB8zLlTLM2Gl3CPW1yqTZXOoiFwDC+zhQIGsbqpee1EUlj
dcxfnmU8DFFYTRhonWqIpHsxX9sInWcApV1xsLJyHegotlLg/o/X1FjCc12k38NL
MEq2mxX3R7p0mrMIYT7qMMZ3Ehazvtr6eYMo1RVspPltdYBUU4KVwtsuMOriDGKl
YKQ6pv3sHhjkhCzm4F7vxxaElomgBMaaD3XJ6hZYIQ+QVZlsaK/igO4GA+HVM3na
hYOhtne69q41ywp1S/k9Zzmb9bGFcGAGiVO5VIM+GIA24vRYJTt3EaFXgc+mIV3K
qxwezrWlED2chcBtMTkBOgxGOJDudIFw+MDSGk1cpFnLGQMYOYipuO85dEOD/clL
hk0fPaWA/CBx5+oyMPogTWeLnTEvbkQ3ZHWF6tjEU8Pjq64QSMTlI8kTzYc+r+8X
591FoZ2HfJmEUvQ8bz3jgfgj6CZZ0q9R2gm7HEUEdnDQbDPrVCRKZaNv9TdppUle
uojCURBt45w3kQ0nRixf6bEbmI+5H4G91UbCHaJSr4/BG7Edx+g4u4rZ/IjILuN5
M/PFZs5ZWfIzh3IqsawiFb3ugI3WGcmAWsKHNALT4NkZC1XjG/eolph34czELlJE
4398z8xNKB3DY1B2otGQHUQGTjUz/WfNhWxMFgtRFDypLF+G2xHJgRi8kd+o8ir5
eO0gkwGgtx0md4k74z8J/sh/s0170LK6oX/MNIyafL8A5xtCxSPjYINFYnwcSFob
Y9DWBEOkUR7yvuenTderAtfnuLLzOCfwYop2Yk8a6D0VdkkJN+XzgdTMUmvVd/49
lUtzC/vIqOYIG8U/RqF8pvNHgQ5lm6kfsbh4GT603YTYCTRIa4vb6VuZ0KXQt0h1
kfBWXfhvI71KdAzduSWcTfRuPmFW+6HsGdPOlbmyab5qzhxJJDXHv7XKCxyds2KJ
aReqzXHyKJkCbtgiDuEfhYWLwHirE7PeonQ+IO9MqqsqHhnobSazml1B7UWG9hOf
g2ztEjk/GIQ5h/bOQGqwfGNn0lX9Qfviw3kDrLk/F6UbR0iEpUSwM3F/YSoD2bvJ
UBZDhJAX9u1S4JcqGtGE2uHQBHKz/7NDbCEASQhIJHqOGJLC35M5xXNVRCoGRvh/
eNZ6NDQhWL074km2xvKU8E/oOo7z6GPxPAR8jBUcBI4vqiiM8rDULXoQLwdMJAvU
oWXx5T0Bno4oc8bmAiUPVIs/Ghp5umACWabi4ZYAnvb3RBCNYunRFOQRebztRW3A
Yv0XfZbwOW3iRKcez+BztXSq4rtZzQ4Ghx/FSxRQhxiNTOfYF9/qBfvvfmOEvhJ/
Jb0y6Raz2ytLIOp7Zfw3pNyWyYcsH+D8wrAJWJWFRCxkmNatCjaJ4AMTVMll5ZIa
GkkkHcMj/+7HM3mkPGXE4wnNam15K/dG2/OsTPF+tru+NtBvnRidsn3G6rD/h8ag
ko7Ul0ZQwipqO+03Spse3xJAoITf8DlqYsC6uIKo1U9rfh78djhbRVuA/w57kpzs
I88IGaUPJrPXDpuKJGa9XpkCK2hlutOpg1xo8CH+Tkail4Nz4EDInuOMMDK6JUHt
yvdwxCXxXzzDwPRGS85cw6qGNc3wq43UWhpmjjEKqUarblPJng1/MtLVGGf7O87N
E+PiCdbVwqtPUUeHIF1JtES162spyPmxbysoBKMqN9n8DLPftlpuKz981ybf0YMM
FaOQpWRr9OKGNktyj0EOjj64lI0XTYJK2fKx7+xwEpi11/DNM8p/GOuwK9VKuAhy
g01xHl2VWBiZFPEueRQX79yh8zAhv6y67qKbKemaeKWSKuEKskPYrW63dSt4ulww
TsjyWj5yQmXvyw1sodl7XMWowEk/NOvlgvo6KW6T4UDvQgUxPPkiHs04x57B99Aa
/xwtdo4qPBjP1U/ZVJ6SktfKtqNSWXT4HMeIuahKfcXFjEGxBK3xTVAHfI55KDrT
x5en354qvBsgmcj2WYXNB9KP/0F2hKNKYeJSy/dtfPwxQLJe6MCHXnfxpPWmUVVP
BGRUHnENFVPxmfYjnQsxdjbzdb/3PzZSOxGxaFydBHYsqG54Kl2ZaIJa7dXEXOzJ
99FERFAQplS24rxl4utp4gdnI+DNbqmSD/8oL99uL76QlNEc4qRZGNwdrvy2sNWR
EnafDUX1d973bUmSi4QsfRxpOimYaVjvYMmdcV3jJTBPU+svWvkqIOJMyb0OJ/6y
vY8KWCxE8GexQp4flKXZ8lUadSgAEJU3yJd/xsInA8UArtdz1DOuqbN71hIoe4/Z
dhlhlS/noVokQqLiO90HVZ4H6skGZHGvekmQfqzUTpI=
`pragma protect end_protected
