// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ART8Tr1hJuDhiZ6dEuF/dzV6w3rJv0DaaDUdBUFul4HlVJiHhhUmRxJu849HQ3yp
En/r3QT+ul11YcZ6H921tp39/kifWUL7bPY89vPgPU0PFSnhzYIG98pBz30glR22
ZPXTDf85mo7x43WaaXvP3Pqt7imrg3bTCw5uLa2noVg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8576)
8/Rk0Sq3H3KkGIhlp8kk+Qwov1qcyoGDcGPYLykzyG4HwTamJs17NfS+dleun1JI
hm9r8QY1gtFhOWaKEfzZ0jAAwSZKgdlQ8MSG+aRdfhZo2EJNbZ4EKlympdpqKIDA
UeyTIviC9dx+JoNzI5rFd0P/5kJkQBB9KkOImIxrO1dVNgzzS8zymExGeDYWiDN+
P45CmXCeS+ykfn5pRNu0jDiMatTQhc/GK9r9ThaZJAAtnanTiTHhPp4c5nCeRHFS
+NPrRH5xqlDQPw8lbnoVmNmEzQDDkgkVc24zIih8zRaGCe+GFM5rdJuy0bacP7+j
tm6PtiNivn2QLE2mhHsddJHqjRcr1oadCalfgWCycA0Qt0OHkA8lRWPftfUTZIJf
DUjZxMbG9Pb4RFbd8pbAMT4aIKbZDQq9e0+D14k7ck4GlVxc6+ywDGahtUUpQ7nA
blrwffinj3R/7bfd96Yjur5/Po33hIaZ+SRI9R5g7X84hKRPDozOjdFzbSf+7Yy9
A7U57Do/TDKyHmd8R+pUjP3G2Jf5DkdjdqUJ+bSaMika/292E8dFVOuC2TGOnmlt
8ao/P+udltfRYlmPT3eGA+3i0UnNdMH2Wu2fhEm2jUKcgw0H+I6ouhbddPYCNWWA
Du3Lg67Du6sKvPn5MbFMF3ajVCdMmGgMyJf1PJPwnpshDi+ThcYRtiQR0dChVGw8
Fg+xU6aMVBbX1iH+IaBsbJE09qZKskHnwTBknJvupZrewiSkprhNZQJBvyaEN+Me
FYIgbuA4tug3yhkjKa1bxnoYeSyQY9KfimbXRX3ZcJOqcSy7desRxLVl61TI12eD
DOqhYv4oAbsBZEthD8bZ0To84ManL6Gn1bnBXdqVbacgLifB7d3qlTk0DKlkvtJB
XXEjdpdwVzAFY5O4nvwuhkeicE4jhllTBEVPkSuxnHcBugLS5Nv41fu3JRaI0rtv
eziw64u28Ay8NPL0hAq41eAuu6pD0xwZukHxssCJpmlmDC4WbJudMBOdDqKDuXqZ
/WXG/qhzE/CR7c7GUAkaDwV0iFyLi0w58m6F1M3+vePUOpueIGrZdyQD60clawjZ
jCK7gd7EILOrZlZgcADqrtRZmhVCQn2DaZstEtu6BB5VMq39jgE1wjjSM9wyVqfh
7MHZ8l7XHcrX8wps+g38/jQQtxBsLzrb0CgM01FOG3UaZLeA0KwcwAGGbyCq5n5t
MaaIBUggwrQnyfmas4wWY0u2zmn+UW1hXl9zonLmux5LlXsge8Q+jIhQPO6Y+VEq
7UEjqewgZAfbpT1Ofmt2UqXUIcy5hOQUZLW+WFTMT1KLMm41DtRVgOhRjoHfXYPE
XMeQ5ri+i7pJ7SCrU1qSZpHtc6wi04c8dU/V0XFLkp4Bquk1REeCh1uHNb2+iR/b
VerkETNCFTREKb2gtor8uwoZDOS6BSwh+mbSBVcZgs3El7e3PPzFXebrNORCtWtd
1UjvsbYlUcQ9mbL3mKSzgpkCQfnw6z86KQmgjXgvcxalhoUqjTndu4q7OCnAf7a2
z60Jst52icgTN49QZkHsGr9XjihleTpWoP0n0otmit1uuHaIvoegiWSEWyjiaPe4
NcY5gZ4PEU+9H4jZ4VmG3tcE+y10pVb3As5bOwzS3ZBu4nQ+WebCd6co2KQ9v3sg
hWbokwSJ9o7iRQHHUd9YNK+o5uKDbn0lEHzbQhFCU8LnxIIFkeIjHsq/rDjIERPq
LqkBGYn5OUpoZPtPgD4TusD2kfqbgvJr2807XrTR6b3xvWyMAMBjvv7K+0dyC6gC
quRT6MxTIXunIsMsrivhVUkn3lCo4024Ehfvkyr8TThuHneuyanr4aNEaWf+0OFc
bmVGSrZHlUzoVMmBMs8PjOIBGwToNFMamfJuWl7QbLAC0vIqPKmCvwL6QnReZBmJ
QRR/c/8P3hdgg+8iv0mN8g5Hd0hzo+ax+OtvcAmxzxakD0BofAjj7XKrBBjjqF9L
2N/L2tZAc0LbkTpZsOsgOmjvGxHcyLSq9JqEnRckbflD2yzzfgIP3IqYChFqLqDT
LrOmlDdmvVy7yXGkjfXHq8pXhhvUvUQpNOztOdK5g2EdnGFq2q82O4NZQ2vdFdfZ
sGY20rNb4Xd/feHe0VOz+mm/BMbsPPrVJ56lgl+jTtYDvfAa0Ac/gVzo5XTDCv8A
qJtm0mVkss1T/ojd+qDEFFguQ9/sZA0fEj795oDAjvGJfK38f7j1iab0W6a1QYgj
enRM3DEEJmPcOaZfJ6dYdGZI/Qg44wNjRDHQvh2YyHj6FmE9ZE7MECZYhZy0rJJA
N5X+hOkh6ShwPfWltfiIMSf11adYERXK0xsqdKFkoBQ1RQ0j15z3ae8KrCEVWt4B
6+CwciRPdHtSeSCJlL41YEx9s07zTW7QKo7jv7sqk6vjilLwQKTeR0v5clkClFPg
Xb8nCgkjImKz+cJdNDHHzD9wj5kK4iZjG56X+uPZEQwlTyezmQVFt1+D4O+ifwUU
fUQCt8CI85ZxgbVx2aZ7BlXazM0X5o7N1yq8iL086P52vGMPYZ+lZ/ZqDBwfFwI2
5kxXupdR8fXjtb6XoSceUJSeQDzNb+sXLytxj33MblPe/Emw3onZKi/rLCnyUjD5
E+MGJgYuF1KhltvqpR9oWFdJdz1rpr8qB2mS4H8z1Iam4SROF6T99uGryS3iLxwM
gUWkLQU21RZbtlsBO2SUho0lFuQBchGJ73GQrNZtY86II55AbVQODK/88Ak9f89K
wNkXk+s2v8iHfPZWRVtPC3Y48m1ZhpWegdoWRcI6PG7mJgMj6ka+N+ugSthRagAF
508lbqEPDMBfXBY9Dm8MAx2PqKt9+2kBah2oi53vX15ecKPNXadDgelSnH0JQVSN
LUk/zdDyD36jtabC+Qd6H6nE89jiZOvKA4AXYxTTgeQ5l9sk404CfJ7omXKpD+C/
OE6yCd26ZQqwvZw22rFW0NO+B6Cecgo+a9ZsKVR22VheC1e0gouDPA/NpUpSuDIe
PZi8SHlyA1jBwf9Yv6HBBhReytgNh3ijqUlP/vdN280go7eMJH6afFaNqd+FOS9E
AuM9NP5Rz3BFbSIzl35eVUEsdW3D3cC5l05AK9oJHOLzpiQdY25s905EthH0wAmi
jfQsVcC4o/Jka2mYjLi3K/2OtltKF7KJRxZPKRy2Ohw5o00T0XwAUqwz6tApP9Lv
dNOabtMLMMvr4HAYHTb4PBiwEddCYztexONk4lPZi9oNsIXbF6U2OyACWFNfNfqb
5FW9IO+FNRljPJLFmLXUCSxiInQuRwe40PmxCJqX9Rh3UIFeMaUbPFR0XEKm3KVO
/8BM7iBKjb2tp7x4tu/sdkuOyqqhfo2hgqlxykjYm3CWqjWJXCYCwx/UZk2QdFxN
34+hgZ+HzMiyTQR1+PR4K4aViGajdy1sTr+uqLGBq6LDGPgjjKICEgRG1tB5FxKI
kM7k+zn7K4VZMRXC3fCD0zTwBlB7DVuFE54oEtVAXZVHh0Eac/0Ne6j8cd6PcKJC
wQosgx32oCoNGgI+OIFas1MSIkQ3re1/ftX6OiceeapS/v0gHKlvqjfj7hejmr9u
tefsqBstDgAXqYlLxyJYjiuSwM6yMo2MXbRLffutCtRj1OBv/gFVZgyRBwLjQGVq
JdjVrGu2cQb4n5TlBLBLq4oJoTiA9oAvEZE9nQ97DXA3b7l8ywv2pGQWcko1OEYv
MaSIHiKUi/4BrjfjC002TD4jP1U1U3ZqXcL+wSJgIUMtLq4rKxYqxGaEVB9az0xN
P8ZWWW+vgqaKpURvl6ex4GSaxDBtgUjsg+4u3VoHxu1uy0cBrrdqMzYZg9bOYKNY
OetPhdBs4kgyYCCced0f4SznQWxnXabqMEhjL+QSCjCkQQ84ZQoZypIj/1LKX+fQ
3JPihHwrWHfo+/ZgaO5TZg7ws7eepw8ODrOMpL6IUeGo/FwF906Pd2vIZ49izr8J
ml9EwnxWNmlezEBkm7/QSgcHc8dw1nuZrzFZyzxbUgrjgLkW1XFTbE14T6dGnkck
lh8JQkR6u5slhNo0r2tBzV6O+iww4Iwr/5wp73eicarTE+6NyINL+HEZ51yrIYxz
UlP+IP31ilBdIIeDakEYBCtR91BOoJ+U/evKRC6bZ/WhkvzGmbXh8eF8wZa/aCOn
bWh6lNfIZYLy7a2LPTN1EeevfISx1vBQwb1g3wXXKz3G0WsS0hCuQDZPkjJPMJnR
/Quenlnxx6Zj3eCNTJoprUKOl7cRBl9QbsRnChXkGT0RSHTElIDIF9dHUib5U5kT
RdPg9UpyRArIjxlp3itIX320nC/ZWwE+MFvCtxko3cpWlYdALRAolT0nahFAJtm3
UOIdWeN+TuW9whUaTPHU1yfkbGaxtfZZ/N/XYrx2GNXINHXUt5qlMpa4wOMThDTR
3GKGoOEKRu1tF+ThiBnVrn1nFwedhXU0TeuIRr4EfbC1kIq4rkjB7VdllkOgt9+h
X9Nt67Z06y2NEsUzXaZfukUKeodo5hCkfksgtjz0LRNKceTc9yZtuoAkxyxrCCkl
vZZGd1ZHjEnOxwePNNGj44MKnXBE5Q1gyP3G9qrMO9Aw1ajL+bEC8nUxgZZAGgdW
SpryktNCdy5qXDDA2gz9Mdk7qgC4rIKKj61W8Cnlys+fbQMpjG/DbhAcBZ4pER+0
EhAaMSAZ/MF9YVrvg5NJMsa48zDFJ4g52NWGZWNp1dZW80WeJ5Y48NX2VTibvsfV
0YyxB8yC9JL6gx4dBfdTcdIP17h7nPAnWt2JKyANkGds0OnWv0F6PZ8APO89+v8V
APgWBqB/xbCY0UADXbXIHY127DURGyBNDOA1Dt331xMHD0zGssXNACK7egVI+xi2
ySG0xuwW+Chnqqa5QPXvZ4bOe0cii06ekHmvxGRo7ryUv8hL+2Inxia0z15kJ37X
p2mfMD8SR+3kEh47BS/nbyZeRfvFpqkRLg0JwDVMxcLf8mHpSibWLPfxELIIfGy7
xNg9lcqibAlugGnP0FTy95QjDhlKHI7cbQtFKIFEo4rNM3qFc3JBbhuCpBzqp0jJ
WOWt0cy4T+QN0MdmVlmRmbs9BCkVa2gwqEJ9iQzm83v2sGuOYWttVerecMC0ov+h
mS6PZEAMBVs8IFqyUpOx6ICAFvu5nFHnDDi1t0Tl6HBgcE5YMojYc/lJc32+QEGL
bAjphT/ZnE0Med2mmsxP8XnXSK3YQm+sIXZdUFAZM7XvqYRbVfVRJ3kJMgpsizkw
0/4Jm/2ZcEevHG1ju70U/Mli6XxY2GtOf5cdShqHxRyjDClNS+mFhqHxtxPTApL9
c+hdvJhVsm312BEE/PIMuL0DxQxq667Fd/l0/sdtHi7AN2z6wV/bDVjXGDf1TF8t
iDcYKPehepWwfMYygHd8kHl28x97jfsIq3IUfu2iPtz9uPPR4ywwBLqxaCJWT7lF
332ZA7OXhOHSiBfhLEHYvab6jsBD/fxpaWX1fa3Bs8kIfhZ+1JGYH73SaSr4ZDd0
j5cwYaOR3zqG94Ej5c64b1cG5pRuYcyWTnjZn9KQu/jd/fi9wm7FweuAZsx33iym
zW9djUa+az0IkoV6QsQxpNOW2HbdRTJWuNLkgYEwk0VRaYSrVlm/KPbfW+3RI2/T
Iag0ZS26Qr2pFEx45nmeun8QQDvKS1RC5aRtZ1QEY0dTC+hOOKjgVOdFVnqqauX6
fGdGlK7YddDhO/t7DrccGrCItp0GBy49Fm/RjQKJJAVk3pVBxkdgd4W+pvJBwhci
ocG58SCvVtiiiWeea4tggmGabrfkMgMv+fu35VQ6pob5xj6SfaytZPU89Pr2Qkye
ANHRdozK8QRlCNE7Km36QOObBBsMoRaYxxNzUnHA9mTTohlqyKh1BZr4bA3s8c+G
cpQgaI1TSDJHqfhpYrXNbbz4O1a+6Me3EELlYcLZygTxtmFVrtHTWQ3FLnR9hn/F
B++2xk4b2yY4dHxeH8kCniD6xdWzutsTOmVyRwZXWdTz4atIyQ9mMjloEfEry/a/
bgjwSfGr+CF3VZfRSBu9UxJk0+G7dAMc35tJUc0f9I8z+DkrtctMTjCGoWqEywFY
un3Kt0g3koqImzTydt4/mQ/zF2oEbwtMsZ+7HGP0OLV5Z8qeszEpLncJp7DCcIXQ
jE0d+W2oPbAkmfAPF5or43yvy6KPf+iqm5mdZ4OsL2ttqxv8T7OfjVSbWRgDsLz9
qywA5boJKimWF5OucwpB806+GOaHFlHDGG3PYTXI3PLcTQ+yIqfdBRguukuNyocv
YVQ8gHqPzwdWQmUp07K2aCjBNjU0c1o14P3H1FoHri6XrjpQHhtbIsAQguFswmpA
fezSAu9BsMb/WNd45ADt8f4V8hY2KVkBfK6OH8QdwDQl41HALvDPhVUb4UjL/Sv/
ojisAe9HjKY37WPCp6et9Zd3x2NggNWZ8nLjeCPYZGzjispTEHhOLV5nBFwxedVu
SYnVQsNIlrTxeTQ1ZQL2qTeDkso5vrJuc3YOU9YJDbnEWJf/syA5QlrIJqtn9hXZ
dRfu1uWaWj7sXeA3awSYO6bePnSTx4BODwPuRoAx7zeN+s71CNA61co4fbgSgKkF
fZCIKifd1zFgweOjTia8I7XyGZv2fBeCCkfrlp5rbrthdqP2ccPDdjc6GeH9180m
+koIBI3NJO4gVLbbKsB0LTkaa/kyKx2bVs9WLyzgiSuB5EHdAia4wQUgw904tuuP
5wqFxasQaZCowiWoynqkViKkNoU9eeTlUuE2smls1GwqsF8DFo7kmtMdIrWLTVc4
S5Sn++Cz9wK2oNBq71n5cFnifaoLHRDCl4f9Gw2bf6inrC8zjPO7yt2fItFEsSO1
lFEqBK9Ozyeu3AfZU2/QFA0A6sdUQBXs1Ys36vsHddebp5tbEaFdiiaZCs9kHmAI
DdQX+NpiVc+oPTQJlUoRnrIVkZjLtDiwUYohGqMHYbBiZAgbON7oxroA+59Jz7cu
+XAFsVaBuc3nNsGewYFVGMVgkB9Y95bvu4V/X5G1G23Sl0pchW7X9ryqzlj6qq1R
2WRg7r2eXOZae/wJmoeXmWtPG/QdkZNxA7ompcodW7RT9a+hBgfwNXhoOSF7yQJM
QocvbdOQkUv+K9NrH1uM6QEjdncXiQX1781CTqdCx3RkNi7UZDTcaX/YWIl19qBo
yUErQbp+JBukLkdTgKIcFVIJ2SA6nRj21Jq5Uc5hJ4ZdmcPPcg++0LGY3nKOH2RG
dlVIv4RGsOUTizLsowx64tXAr0BJrnzSrrrSBYSw1ZcMTyF9giTPOHwac40X7xre
GHBAgVSFutRujXdoVe+Hh9YDKfEQ1zOffkpmfMreZQ8LbiIazbZRIqtgAsBgALYd
rU/EBzpqGIdoLd9ir2oB8oMPLt7yVOxRZmrK2gNFmoHt3eIFyvGOsBzBIlMU028H
eOiDaE/jf3x5Vb2aF/hOgqQnFmxO6qjW+HIxkonQGFq+HH9ojWrV/ojvjv1WvwTC
W0Ph4DpQzKWlx7/v64X9RxAqsUuF807RoWsl/+t6F9Omw1cuFCvnaDinTJszjzyh
a9Lxv/mAgDHDPLqU8ka68U9S5lsLNRxf5zf3ctEtduKZO3vgMezIV3vuHL1nsWkP
SWYBhQ2l2sMM+kO7KlqsJpjJYNUo4xljX3v8TfkWbxJFsY6VET5n0kug0iUqYFou
N2OETOQbNY9qL4v5/Pe5YgByw81iMCw6Du/pepHBz8bgk7MyS6LjxyoZhIyAbIwk
DrO3Xm7gibf42ZfAJRpgDtb0vjAMgCRuabejWHwFVX5NUwo3SlEECMSBznF6XzLv
5hDCZAg88gTZQwcikpp7Nkojm1w1GSsVduYI7atofOL+KLVCb4YFJVQJ4P/ZCZ8E
viIT/NPmnQIsTrZEI/yfzZ0bZinvrQH8lFnWprOdNsay8RFRakqnbB9I8+PDEJME
2To1Rs49c9RBllgVgmmGtYSFlqVwtXmdORUupn1AC+o5Xapv9j0xwHmFmzby4VcI
OpwZtIH8cc/brcA6Ca6KW6B14WHGlE8R+T/kUhY/v9UxIsCjoxWvPP8m7iZ6X+BK
gEGnCuMYovJpRLWcrdra+ef5N41knYV3GSxH9y4GJrC9oIEZXdVdGARkw1WK5cef
RZRDAShk4aLt6CPGTmOcve2iIztrJx2aduJXF2pLNQ1jjnX2UHsm2ELLmlca5Ufu
vpk3s2vWjQELNGSS7yb16oh4mDEU7bt6cVYFFkeNyirkccNvqwDMTIZvGJ5QROba
zbXhu1zN6MteKSZg/f+BXWnm7U8SG8MnGDeK1rsAaOtXbb4pZQyj41rn3J1YNXMZ
Zbkt2stXMeZgyxRspYsgo/4g9KWczImZ0TkLwYCiK301QQUj6fm1tL+lqJhYBclf
ybtIfkejbgbRZv/VfIQJQP82JZuZ6qHqSzH9Qb02SlZOCY7OZiBoAfLG/E0b/xxG
iA/y6V0MkTvqaFljNWewNS2H5FyJXt7ypH91No7Q5dcHlppuxvs6qh316lPb3E3Y
CPpUcjW2JZggAPujftYy0NC+osUYDw/DG3LMlgq1HUEq7yVOh0sZfL+Bf79d4Low
YNKZuq6g+RKLedGGE5ZCP16HDJg2cybDdfGmMmFldAwFanc2akseT6OEcLeJGma2
gju8YYGeF07MTyAS7e4/emW9sRBJuadJiaH2NYN/vb+hf5YVsYFv/z2fTGI01aO9
aD/+Wwi2WqQRpxYkQy3UDTLJliYx2hvTIWQLsMRfjDeErLaGUCxbfVs2DIvW8LEW
SrFsTgW+ZtZkoZyDxjwQgV6QRmI3aRkrVhzIdtENsRb6ZWZNgwfW6XUvVsfkLcIi
RMXN7FL1VFdF9vQWrZdF2bhrKFCQb0RJDAVnfXMdHAB1hEMfvJ31gwLKXGqy4msp
39/vLHxeHF62XEbc+iFKo91jg3TcAYW+WWsPJ6D2p76IDHJwbtKhUvxq1i4u3+IF
gHX0B4uaxo4c5pgo3ZALB/G7yP+vGLSqlnj9DBdCNiUJFLGQ+twHMdudQDOld4//
j3Z5P2zYWCk5xOhVu6M/muV9y0UU1ni3Ss3Gq8IKclib+XexS9HLfTUJHONmJVQ0
HaiNYz6IfYSPf2AIRak5gel/nBLeDxVah90GkIz933AIHqMv4bPyKEu2cSUe71/z
nA/Zi7oVY1lsOx6jk71HRg6aBOBT+t/+pJDmpOXStC8cZP0qpYk3pCn8ea3mwz/d
WQ5D6Xh7cuC6B6kuxEWv+RiWubpM4ptDbbDBKTzKJnb6iloRC6jFg2Kj54IzIlmZ
9nFURBMStvDcVWgNE+MhENGtkRNYlYZ8N41Yd08+nNwue3MybkgIpajpuIpYxotP
dwvmEN65DFMpWax1rukkiA+hQ4K1aDJDbVbe4H1c1IC/BZKkvLYCr2UENuMlGSCH
UYp5T/bu2uRRJllPMInYiRw8RnYt2d3khvFjDw9L5YTjvqAVFTdP1xQv/qM5OZ0w
ohSC7GdxW8VyDPipjgM1AtIvN4kwj9JedN6mgGTnRhzNhQbtUW/w+Fa2zFp9sGnN
/Tt3ifWXxdWg4TF24kvvYVlBE4V2w2t+pGiYlgm85DKrzUVGLiUqWBvxsb2w3g8X
qj+I92yiWttUNjqkVSPPAu3J0jU1EIy7nQgWxNCZ4faWFyFH/0N+OA7Yro+hbik8
MyBLqdAT+u5wBkxeeJ5jal7axVeCHmNPhzWdqobxLhoLzOr4VRl1yDS1Q4p0vcPl
3mCDGmdao6Tjc1YRDpAZTZ4+6plENzQMMdCLXXkz6AtEY2SiitFgS7ehHF002zud
7YVzOOxyUtoUOibumAw5ap1oppLbUkMuOQqUrTq56JqlW0kamwRZdSfc+CdzRjrQ
vqYdMr8P+qBkMSOAGfTZ6w7eStv3cQE9a3r39zbsYcc2fLepdH9Er0VHtiFc19jS
eS/mZdilNTkVxeRI4WX2Tio8OasqbrfFNYQx/2j07gbu/HL20yiXeDHtzwfu9I6X
GqlQje7dT2r+FgoBg0g9yx/Fi2C/UIkLHFB2Yjlc3Y9KZwpYrMSj9JfaZPGj2zx+
lLpw9YntX8Bl7dt0n5rI1MiOjeD4266E1eswxSIsqTWezlX46m5kEO/0AqI9oUxq
CmCxLSZjaf8rhJDTlKBW42j0R+kcfcbVzz/5H8LGH4DtuyK5MqiOsHlGj431vqfQ
Iqy4XjHi3KsQ4Fix+D2LT33iw7QLLuWqGk24QpJu4FwoO4sNXI3ZD3sD3MYOwQtK
HWDfaJuOKZchZbOUtxeIA+p+kPrrhQScWb4SOrSPurze67vSFV/mKxvA7doiTEuh
2zy7ppfXnzBwFRo7SnKrmBloJTWwMIso/6gsL2zU224uLvFeK7iMab1vom1X0hOW
cBOehts5jxmMdB+S3v/Ed3cwUD98Yiya/cR4nL40OKq+jaCK0NfHpTMUT5XukI1T
X6E5tpR875JshzLYzd5h65ID6K8h2BZiFZBrlaJdxikIvJqdBPKYhOI8tQvFeS1f
Shxopqy5xpV5LRxXb8aj8gbNq0maxrw+6aJg7YQBs9N6YNolMvk2/4x0mrodziJp
0mX1WN6lVaIaAvl3aj8RwgOPfhqlMKguL7N0CT0UGgHLOhf9twE7s6QTcraLBWvr
cOwabtO/zezVB5zRf+tMi4okOsrx4AtGuAZLFJbDAPOPM8yCxhmy3cR/Cpe4ra4S
YMR3rbIt+htyF9K8sDRgUh3koc+LpSH4XNN2KW1s/KcgpO9q1Qq+11JQUgvZ+Zje
MHijU05svgCP0557ktttiRLI26M8BuaT4qHYJrBLB7iODeTeF/++qHzoJklktac8
3p0j0UI9v0nBk2gJxNtxdBlnTb70WuYfXkYIhfzddXfSt2lPXFttLoOfG7DI447E
uMqyy1+Xgu0NO8btSVJpnzWD45dlkqrTmGYmL5NU6SeZYKfYNiCwwGI6lGJhg02l
yATGEXTHmhDQF08Xt/4KUBqQM/VsRJzGqpSpI6gbmZ9J8bmfLialh/drY+lyMl4j
cHFdpi6E8WMdijBuNbEjbxoho+iqVhxEgmHgbbqnx7N6JPn8F7FuunZ0yY6t9EyP
XoaO9tC3WnGgjLlU0PPOCYwgMreDt554+SnRithphSDfjBSJp/Z3sUs4XjIsCNYk
N7BVxtPpKrKEUIP/yyzAJe0IlLB/5GxieKNmPibs3Bw3yBtyFrGSBLkYK0qq8333
EGsifneL81BnHZF5KOqvSLcjoYBNV28FlV05w7IeC0W0CbnidhPZSHE79BcpmeTE
JescMEEpkbSSrmEFDeyYJTg17DJC264akkfmgSbAv59dSoyHCImwHt5F+Zr/RzNz
Iujsfj689ncfd1Hi1/Kvg1vPFY6j1jRO+/CYudusKOHWCKF1jfN0yTbawJs0QFW3
1zH8K0KFsBQ9+7KbVPvyip0xBuA04vmJmKRh5Mw996U=
`pragma protect end_protected
