// Data and address widths
`define REGFILEIF_DATA_W 32
`define REGFILEIF_ADDR_W 2
