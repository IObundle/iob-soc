// megafunction wizard: %Low Latency PHY v16.1%
// GENERATION: XML
// xcvr_10g_dummy.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module xcvr_10g_dummy (
		input  wire         phy_mgmt_clk,         //       phy_mgmt_clk.clk
		input  wire         phy_mgmt_clk_reset,   // phy_mgmt_clk_reset.reset
		input  wire [8:0]   phy_mgmt_address,     //           phy_mgmt.address
		input  wire         phy_mgmt_read,        //                   .read
		output wire [31:0]  phy_mgmt_readdata,    //                   .readdata
		output wire         phy_mgmt_waitrequest, //                   .waitrequest
		input  wire         phy_mgmt_write,       //                   .write
		input  wire [31:0]  phy_mgmt_writedata,   //                   .writedata
		output wire         tx_ready,             //           tx_ready.export
		output wire         rx_ready,             //           rx_ready.export
		input  wire [0:0]   pll_ref_clk,          //        pll_ref_clk.clk
		output wire [0:0]   pll_locked,           //         pll_locked.export
		output wire [0:0]   tx_serial_data,       //     tx_serial_data.export
		input  wire [0:0]   rx_serial_data,       //     rx_serial_data.export
		output wire [0:0]   rx_is_lockedtoref,    //  rx_is_lockedtoref.export
		output wire [0:0]   rx_is_lockedtodata,   // rx_is_lockedtodata.export
		output wire [0:0]   tx_clkout,            //          tx_clkout.export
		output wire [0:0]   rx_clkout,            //          rx_clkout.export
		input  wire [39:0]  tx_parallel_data,     //   tx_parallel_data.export
		output wire [39:0]  rx_parallel_data,     //   rx_parallel_data.export
		output wire [91:0]  reconfig_from_xcvr,   // reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [139:0] reconfig_to_xcvr      //   reconfig_to_xcvr.reconfig_to_xcvr
	);

	altera_xcvr_low_latency_phy #(
		.device_family               ("Stratix V"),
		.intended_device_variant     ("ANY"),
		.data_path_type              ("10G"),
		.operation_mode              ("DUPLEX"),
		.lanes                       (1),
		.bonded_mode                 ("xN"),
		.serialization_factor        (40),
		.pma_width                   (40),
		.data_rate                   ("10312.5 Mbps"),
		.base_data_rate              ("10312.5 Mbps"),
		.pll_refclk_freq             ("644.53125 MHz"),
		.bonded_group_size           (1),
		.select_10g_pcs              (1),
		.tx_use_coreclk              (0),
		.rx_use_coreclk              (0),
		.tx_bitslip_enable           (0),
		.tx_bitslip_width            (7),
		.rx_bitslip_enable           (0),
		.ppm_det_threshold           ("100"),
		.phase_comp_fifo_mode        ("NONE"),
		.loopback_mode               ("NONE"),
		.gxb_analog_power            ("AUTO"),
		.pll_lock_speed              ("AUTO"),
		.tx_analog_power             ("AUTO"),
		.tx_slew_rate                ("OFF"),
		.tx_termination              ("OCT_100_OHMS"),
		.tx_use_external_termination ("false"),
		.tx_preemp_pretap            (0),
		.tx_preemp_pretap_inv        ("false"),
		.tx_preemp_tap_1             (0),
		.tx_preemp_tap_2             (0),
		.tx_preemp_tap_2_inv         ("false"),
		.tx_vod_selection            (2),
		.tx_common_mode              ("0.65V"),
		.rx_pll_lock_speed           ("AUTO"),
		.rx_common_mode              ("0.82V"),
		.rx_termination              ("OCT_100_OHMS"),
		.rx_use_external_termination ("false"),
		.rx_eq_dc_gain               (1),
		.rx_eq_ctrl                  (16),
		.starting_channel_number     (0),
		.pll_refclk_cnt              (1),
		.en_synce_support            (0),
		.plls                        (1),
		.pll_refclk_select           ("0"),
		.cdr_refclk_select           (0),
		.pll_type                    ("ATX"),
		.pll_select                  (0),
		.pll_reconfig                (0),
		.channel_interface           (0),
		.pll_feedback_path           ("no_compensation"),
		.enable_fpll_clkdiv33        (1),
		.mgmt_clk_in_mhz             (150),
		.embedded_reset              (1)
	) xcvr_10g_dummy_inst (
		.phy_mgmt_clk         (phy_mgmt_clk),         //       phy_mgmt_clk.clk
		.phy_mgmt_clk_reset   (phy_mgmt_clk_reset),   // phy_mgmt_clk_reset.reset
		.phy_mgmt_address     (phy_mgmt_address),     //           phy_mgmt.address
		.phy_mgmt_read        (phy_mgmt_read),        //                   .read
		.phy_mgmt_readdata    (phy_mgmt_readdata),    //                   .readdata
		.phy_mgmt_waitrequest (phy_mgmt_waitrequest), //                   .waitrequest
		.phy_mgmt_write       (phy_mgmt_write),       //                   .write
		.phy_mgmt_writedata   (phy_mgmt_writedata),   //                   .writedata
		.tx_ready             (tx_ready),             //           tx_ready.export
		.rx_ready             (rx_ready),             //           rx_ready.export
		.pll_ref_clk          (pll_ref_clk),          //        pll_ref_clk.clk
		.pll_locked           (pll_locked),           //         pll_locked.export
		.tx_serial_data       (tx_serial_data),       //     tx_serial_data.export
		.rx_serial_data       (rx_serial_data),       //     rx_serial_data.export
		.rx_is_lockedtoref    (rx_is_lockedtoref),    //  rx_is_lockedtoref.export
		.rx_is_lockedtodata   (rx_is_lockedtodata),   // rx_is_lockedtodata.export
		.tx_clkout            (tx_clkout),            //          tx_clkout.export
		.rx_clkout            (rx_clkout),            //          rx_clkout.export
		.tx_parallel_data     (tx_parallel_data),     //   tx_parallel_data.export
		.rx_parallel_data     (rx_parallel_data),     //   rx_parallel_data.export
		.reconfig_from_xcvr   (reconfig_from_xcvr),   // reconfig_from_xcvr.reconfig_from_xcvr
		.reconfig_to_xcvr     (reconfig_to_xcvr),     //   reconfig_to_xcvr.reconfig_to_xcvr
		.tx_bitslip           (7'b0000000),           //        (terminated)
		.rx_bitslip           (1'b0),                 //        (terminated)
		.tx_coreclkin         (1'b0),                 //        (terminated)
		.rx_coreclkin         (1'b0),                 //        (terminated)
		.cdr_ref_clk          (1'b0),                 //        (terminated)
		.pll_powerdown        (1'b0),                 //        (terminated)
		.tx_digitalreset      (1'b0),                 //        (terminated)
		.tx_analogreset       (1'b0),                 //        (terminated)
		.tx_cal_busy          (),                     //        (terminated)
		.rx_digitalreset      (1'b0),                 //        (terminated)
		.rx_analogreset       (1'b0),                 //        (terminated)
		.rx_cal_busy          (),                     //        (terminated)
		.rx_cdr_reset_disable (1'b0)                  //        (terminated)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2017 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_xcvr_low_latency_phy" version="16.1" >
// Retrieval info: 	<generic name="device_family" value="Stratix V" />
// Retrieval info: 	<generic name="intended_device_variant" value="ANY" />
// Retrieval info: 	<generic name="gui_data_path_type" value="10G" />
// Retrieval info: 	<generic name="operation_mode" value="DUPLEX" />
// Retrieval info: 	<generic name="lanes" value="1" />
// Retrieval info: 	<generic name="gui_bonding_enable" value="0" />
// Retrieval info: 	<generic name="gui_bonded_mode" value="xN" />
// Retrieval info: 	<generic name="gui_serialization_factor" value="40" />
// Retrieval info: 	<generic name="gui_pma_width" value="PARAM_DEFAULT" />
// Retrieval info: 	<generic name="gui_pll_type" value="ATX" />
// Retrieval info: 	<generic name="data_rate" value="10312.5 Mbps" />
// Retrieval info: 	<generic name="gui_base_data_rate" value="1250 Mbps" />
// Retrieval info: 	<generic name="gui_pll_refclk_freq" value="644.53125 MHz" />
// Retrieval info: 	<generic name="gui_select_10g_pcs" value="DEPRECATED" />
// Retrieval info: 	<generic name="gui_tx_use_coreclk" value="0" />
// Retrieval info: 	<generic name="gui_rx_use_coreclk" value="0" />
// Retrieval info: 	<generic name="tx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="rx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="gui_ppm_det_threshold" value="100" />
// Retrieval info: 	<generic name="gui_enable_att_reset_gate" value="0" />
// Retrieval info: 	<generic name="phase_comp_fifo_mode" value="NONE" />
// Retrieval info: 	<generic name="loopback_mode" value="NONE" />
// Retrieval info: 	<generic name="use_double_data_mode" value="DEPRECATED" />
// Retrieval info: 	<generic name="gxb_analog_power" value="AUTO" />
// Retrieval info: 	<generic name="pll_lock_speed" value="AUTO" />
// Retrieval info: 	<generic name="tx_analog_power" value="AUTO" />
// Retrieval info: 	<generic name="tx_slew_rate" value="OFF" />
// Retrieval info: 	<generic name="tx_termination" value="OCT_100_OHMS" />
// Retrieval info: 	<generic name="tx_use_external_termination" value="false" />
// Retrieval info: 	<generic name="tx_preemp_pretap" value="0" />
// Retrieval info: 	<generic name="gui_tx_preemp_pretap_inv" value="false" />
// Retrieval info: 	<generic name="tx_preemp_tap_1" value="0" />
// Retrieval info: 	<generic name="tx_preemp_tap_2" value="0" />
// Retrieval info: 	<generic name="gui_tx_preemp_tap_2_inv" value="false" />
// Retrieval info: 	<generic name="tx_vod_selection" value="2" />
// Retrieval info: 	<generic name="tx_common_mode" value="0.65V" />
// Retrieval info: 	<generic name="rx_pll_lock_speed" value="AUTO" />
// Retrieval info: 	<generic name="rx_common_mode" value="0.82V" />
// Retrieval info: 	<generic name="rx_termination" value="OCT_100_OHMS" />
// Retrieval info: 	<generic name="rx_use_external_termination" value="false" />
// Retrieval info: 	<generic name="rx_eq_dc_gain" value="1" />
// Retrieval info: 	<generic name="rx_eq_ctrl" value="16" />
// Retrieval info: 	<generic name="starting_channel_number" value="0" />
// Retrieval info: 	<generic name="en_synce_support" value="0" />
// Retrieval info: 	<generic name="channel_interface" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_enable_pll_reconfig" value="false" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll_count" value="1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_refclk_count" value="1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_main_pll_index" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_cdr_pll_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="0 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="0 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="x1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="0 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="x1" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="0 Mbps" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="0 MHz" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
// Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="x1" />
// Retrieval info: 	<generic name="gui_mgmt_clk_in_hz" value="150000000" />
// Retrieval info: 	<generic name="gui_embedded_reset" value="1" />
// Retrieval info: 	<generic name="gui_split_interfaces" value="0" />
// Retrieval info: 	<generic name="gui_avalon_symbol_size" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : xcvr_10g_dummy.vo
// RELATED_FILES: xcvr_10g_dummy.v, altera_xcvr_functions.sv, altera_xcvr_low_latency_phy.sv, alt_pma_controller_tgx.v, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, sv_xcvr_low_latency_phy_nr.sv, sv_xcvr_10g_custom_native.sv, sv_xcvr_custom_native.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv
