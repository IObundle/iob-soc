// SPDX-FileCopyrightText: 2024 IObundle
//
// SPDX-License-Identifier: MIT


//empty file for now
