// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VabeGcDK9X9jMmGOA7aZma8uLXsu1hXsFD1l2bMPl3foRQKB7pw3JrWGl3e7ROaz
9izsPAL5yTtwKuODD96Pb1hVXtOcoV3cmyRIokk5pwaDzfngmF2RMmpvbK5xul9s
zuICe0mDSllXBEzMCOiv9uorRA2J8js8useuvmkUPek=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8896)
RIxFZCvhlCxidlqCJEu6+8I/8Vp8Aosa9dAIuuk2xMj0nKsK0Tuuk0+6kvAm1Xuu
XnK0jaooeHNA1W/c3EJIXhkgC5yoI6aMt96brE0IwwRwuZWY6n0krGxwc85aT4b7
XAOdvovnb9FlhMvTaGtPweMFuRtqUhhrotzR3iJDS5X2tug0U0Z5YTIe8HV23n3s
/Ovex20dTF5S84+rz36vsL52wx1IdehoxgyXmVD0YZ915ohgjuLnaAKrKmanIoYU
egFkMqV2p/KZWL2kpXDHwIRh5OVmieH5hzsLpAgzEwEa1h6PQ7HLQvldfFEdsdT4
oOhp2Vr74fdNf6AZZDPuOFH1FC+nEcqDNvmJtbjmiSc1GqX5KjA0P0sd1GoTWtCq
2GMv7eiQ/OQMSqfKc7kexWB54tGUEfA418b43pjm6N1gUr7MU81P92Y7xsCjMbuq
b+WVflYtZSL8h2S3c4O8LcX4EiI+EzPBJy4eHWiL/aOnFyMcNlOglrwrI8BHj0aU
1OvVF4Mh2Nc38/RlNrGwnUHI88+iKEPjl68p81+Xfi1ejsJwmIDVfgCDd70VwkNy
Wgq4vZormm5xS9q5g1oS8AwPH79Q9Mo7pVummk48SaTpnSrPgrgO1WlMeLcNQl/y
cajZAqmtd/nGvZtUFpPZaIciu4CarmIoR9kau4ebchdZmaEJkMVtLkez76PgbpHy
1+8jQVb1Fz3Zq2oj5X2H6HhWrbIvVPON4CQ7apvWmhJZFe4IqI7HUW5TyKxCZcLR
yohRruskYC35lSaREmzh0OJs7+grCvhufTnAe+CoVj9YI4U9TsNB/ERw+HreJVyy
MGdEwRKBNNx4gm4m9RD50r9cqxDONJn1vhGHfXxfPfz+tB4ylaOfvk5hBGu5oM5N
Q5IE5IkJuubCWakZoFKYKjI+3eddQF6hDCTFS1C698jrgwUAvnV4Qm6D4YnPsspu
R1f+C55UfPKIVlQuqOMPNtknQNkJe3JZdFMjhkRTb3rQGyJZRFYJpOk4HFkH/kkw
LNJMTXOumrKqaofTmfxnolV3shaXYK+vJ81K15ke1ddaQEq2v0ntmsUm3IQti1sz
YZuQMB/8bCW7NXWIoFm4dGI6zDSXf53EMN59kxfu2qy0hvnyzIXiSQJROxAX+UWa
Hdj7Rh5W+p5e2x8GbApS/YAAJrzLoDGm5I7gl4Hep7j5RhGSSNs1lbS/f0UvYRPS
ncLmREIChVIL2E28u9K0OHDLLkjeFOlgYO/7n29EwL1lMtZMu7uw/5fB9wj6qP/j
otKhZA0MgEOPZbC/l+TWV6eCJF8BPAgieoIots6LMLyEybi+/otCUBfBooqFfsqp
qiqwLZzv4NgJjGbaxaXNVKcJU2Rhb0Af9uSqytCkStsm6+w/n2mVhhhhoHASHwTM
95SmrYiitqvEN+yHoBQqct9h66by5nVsS9yX2YACpdsUT9huHks8+7C9zDtgEgSO
NMfGSPtL2awczuXhtXiqrbHY1ApfVvZGzwoGepsGcLmJxV7IiJaVv0ER97gyF1CC
bYXjQpIr+PtPUnP9/P22KAHvFZvLgbxXtON2f5bafC1hsR6QGG7jZ03YTftkey7w
YIEQSyCG/iZv5fW1vJplt5wHLMIXJtPtcpipQqXJi2X3BqRVXfDz9iV+3ixIHEDl
JgsBbbwVNnSFGx8QdtodOKDZcJqQe3QBN66bnCnVRBGcmAApgJucIoRr7cMYgjBu
o+/sOfQFo+YtnNqtgy1pnluR68QEZdC2nWqAHvtJOlVUGJ7CXX1eJZnIrU3g9OMn
dJG6Oh+L5szMoLP6pix5g8cgVahOE5eF/opcrpTzViAtIDktOArYAWlkzJ6GGfC0
4UAUH46bU5vKSjoxheQqfguC5eFmSCLdeJnUiRvke9dPQbH1NGovYAPBZhbXpja3
PTSahXYNn4BHdjEOoxNHHxykaCb3rur7SrSsrUlco8BpUjqfwFlq+im0TWuwb7I3
qGwN8rasVdpO+M7J5h7y4FcOdG8tptn0zpvb6uD3Np2N26vR8PfVCWmUOKMbVl1v
3ewERsLiNFBWLE1FSoRiz+WJT/meO4XLmqm9cR1akSQEYk1+sZJ5PcHFgt25XuUu
t7B1Ays7TjMNPvG5/XbOVgLg2uh+UuZzJ3p99URZvv3hvqYqH0QFe7wjgtXJhW1o
wTkD/5VYZ64Y3tNz3CAXdAADnfnSDE9vbTP+7qBQaNlqxp93Fx3M6UZhB/K7G1xI
VB+s+s5eJuGdukeWBis6PoIpEzgtADwl13e5OUsQqqFqyvs6dY7l8taHXeQAG53V
CbskungodwNs0/jsNYSJW1aUvz1Q0xchccoEaEIAecaOdrVAklnX3VV2oJewSfmv
YuUEp2QBr5MIGtyxigkdX6DEJi6o62grGc4Aqc9T71jXH8ZyzUq3B02AF9vUPkxK
K0hcEf9t1G5PmNW1CyWKw6WLeDitYCjn/JOPS33RzXP/CqrGS+6C46Qkgawggder
3WC9LsXA49QqOOGw/z9ph/Yq/69oQxuQqaQ+d9Eb3zkR/yfENc7H1BSg1xToRMmx
atGq4jn54AYSfkZvi//3V3ViKC6F4in0yw43fsweATCAJ+1UOB6khQWB3vqGT+9d
BNjdDv+U4rJyVmRyPUfSkgdpcr/QIZyNvWG/bi5qtW+vMfitmKO6kOUNGCKVtIcL
5gWe4s6Olhy33pgGpGgc3I7gmppW86OQiHimEOrWUjyjc4+Xp87PZfY+poiRjJ2U
YNW6PpHhCAziKbe5jaOv1k0Sgwa8+2fsAb8OPFNA0kX3TIWHm95/vQyF01KMWNtM
Iso6rIMkYlTOd6ukMA4TwNjgQKf+a2Yf2etiOZV12Up+vSd/q0QEP1a8DD1KDVIM
eeAP1jqKZgTT3q7a92VR0pO9/mJLa4RjA7tFF9iSuowF3gAN42EHL/o1KTvkwla7
w0VGgnWn77d3LvJT/PI5de/mtsSh4VWOqyZIB3mzNTaPgErcLInRYRITFfvCrk3m
REbNMXIf814sEqZli1h1ITE8eN0VydPwW17+pE+7tU4ygQT5QMWnSieUWTNAmos8
cDSMMrUK7WpdV7izlqKIk6os4hLcXK4+nb/7oBWF7V/YJXtLjfG3uu0ffiZrrW2W
fIyP5xcRza5v05SEsKSZQrYMbK7pnoyYaci4owPj9uAmyyGWhrwmLudL2A3+3UJk
I5h7Qn7wWedqcrm1di0dq0ZIrCTSRYayDn9ERrVsyoFaztUrkBEN6ZPrnvPKBxxe
SO5GqEzRlpABfTuc0LMGRs5cu8Wf6Nq0JMNW7aiF1GglR5uSAle//EyYJa+M+nlr
leSXrY9apuOjfQCxv+yEW+OzO+qLXOYat22W7bICzqYqiRGQBhTWKE0zSoHUb9Im
1FivezqT8baX7sdaKN+lMZq1Z8i/mVF7jwWVrMJLu7dPHDk87iUsUy3r4H0U1WQz
2ceGs8zliP9dIVgKrsgLQkPCcMUB8i46Q0JdUiapSstz/72WtJ9ijxXSj9YFwj2b
B5ZpGPzJ8Ln7uY+seBaBGN6KTv6HCRHcPCnBqAdxvt44HuAQO+cJ0Fqh8bM7NHuO
XMo2RS5XBVcUBMN/ME58oeklDVpHxWi2Sqz4F5GQq9NGEHUp2GiZjXPfaYO6/IHK
NJyJyrVCdxiUaOBRLw6MbXJ1EnIiSSf8wz5C0SCsXQ9UT13r3PMNg8p9C+66oE9v
Mu1TTxZVIaYj3Atf9hCtcR7Kea4Vg7DUXoJAk7yRUZc0le3PQrwFIpuZ+CaBOyW+
b16YKDdbBP7mMHdS/PTQrkK/qX2vyl9v4mZ6IM3TaDycBazr6d1pOhnSxfZa7DWZ
/hgTucV9NDmCVmrW1j2SzRw8NtKHSrsK77DRGaC9B8KKySH5iLxTskrzkWVFhDGM
YzKYumiOIFzWn+s/o6QM3bENgBpPKgACPptiJBN7bpVBJxdFS9pgRfh3O12AiAh8
Wcta77/GUaKhkmsHAxlV+4Oo41o8Y7UVaI+1F4hRL42610g3nhJQaEWpQj6uugLX
X+ufzDIb1GRMAwVdWebs4fsPuO/dLfA1C9rBZ53xtgFC9pGBzD63BX78VbQsWohM
fxST1c2ZaK5UiXt8LxmatGg3B3VAouPVmRCt4ZmXGFzZDmZsmZoEarwDAYF117h6
6krjTmA0ESX6bWsTke5EdDOWX0p0VRXFzZxwouRdc0U9humqYcLI3Rx4buFM1nxC
iFK2/trAZ/Vxsfgtbte62blkDOxWhmsFiZEPFG9h2sY1gWJTXcazhmQFYj6kFpim
jj3Rm/fgGyy1grFqZY/GHs6bQjod4xULk7Rc7EjZdIu3ljckXAnQ/WVUsRSxW7GC
B5XxQarSsJL+XZolmTUklr7rUFgmQUAwjr/5mTi0N490sEhSc/pYmPSI92tag+8K
4Qqg9ifUWaSOZ1Us9izLwgk8eQEh7alIblxFh8dL2izjuO2jQtIUaHu2CojeyUs/
iSGm0eLCRy4M5T1DR31Xnr8qgevYlFohVkSQsT8eEKMrMVFnix+cK4la/01VGcxT
qKVGukAjyH/PpIiGe5nCM8melHjhslt1FI1fD6FJ9JezhaRDBG01iasCzPCaYjFc
ILnUoJWmRZdAE6CONqus5nR9dLIf+YiERqxJiu0Y0dgp8xvCuWkTTxvCuTqgv7CW
b62wPuuAEHuQb1SarmRuc/3SKOWfpvgd7EJkeihImBdbSu3teaxwXzQ0zU5rWYQe
uFTjeT+KX2JULzblPq8V7Al6Qy7k+y3qTeX9innVONgzI6oTrvivFT6RRTXi4ucF
sCScOgzLbnIh8UnFXrKtjwcgfx7Gq6MzkFzIE/cgZ3N8CKoGXW/101P6Ph/KQx85
gIyMlnHtWuFXOVLDTARRVM3xVCn2/ifsgS6jgVTXrV1C95EqJSyXCE1bWQNum4oK
kBHHEydWYNTHyzokJwMUT6XLP9ulQgfHAxdXoe3XqluDCAVMtVHPqT/bNOfkpKzO
ACMqR93FzSAmg40QgyL6h+/0g7kaUFGiauF8lDMEQrO979lyqU7FHvroDFwOmokY
/jmEEC2KC5TIsa8PIQfuopvrbq0H+K+Lm5caY2R7AufhzfghNBIGaYAMZtjiDYkw
SDCbhEQ2EokANb58SK1EQo73IejUYAn0aA99YIdEMUFxl1C9CoQPcoqLjYbJgkmu
uyjL2fW499WAjAqvx2u22Q1bx1em37yC56lm+s7pbl8yYRt7R4L4o4Owdws/mfZB
/VagU//TKiN6ITTVoJWJ3J0ap12pnkfGyfrFw8T8IN4u2x+aWINFUbeJaa/1qk/G
wLrc7dSPgQYCNLb5qy+LviQ4Eg8hjTHdA00PiADdhh8GF+Lshjj5s0db+Dw01qYr
F5hxPl+XYnWAeHVyz/o5KZbK2e9dDly/RdsoX0nHqLgAy9yTgBDW4JXoG9vPkWNk
Oj4JmNNaF9FK1bhhikOD/FAFtjbw5RevIcVIDOXSecdrrOknQRasYFhPBnUysmOP
9D0TpNKDob3jwBhrhJrtDpezY8LmPpOP/RbgIC9a2u7+iLOMaBQc+MhAHuM7EF7w
F3P4xZKrv8odSHmKXVWDhp01xf63NMMnF9KYGDF7DTY/9TLJ18Idcllx0dnXIwRn
H5uKC6Ci2J3Qfbu6lM2memEmB9wnE8H3SamJzQR1pZaLwB8aHj7s8fkvDsUFZz/i
196dvYHgCaoD9nmdHZEQuHuweAznR240u9UIEY38c3p3R+I7mDU7qRIf6/Qm9LOt
dIL/FuO5kJ8SrpbFrjxoJfC4RQf2uXc17RMElLI/yUW6VMSG9dTXJKKMZlFP1Xnn
DQ/KMymDO3rNjjZdHfEtUVhVOVGNXLp1IyYK804LX/skv8XX6l6yefbTmmQitwHF
A9r41umtmixNyipM5jWVFcydt0esgC+VMDPuFbj5Uz8MLHGiFF/sbE4JpihMawC1
MYNcc4Hef1klNsv3vTt0nFFFFT/+YWMVXPjkItSdX7hALlJjYaULQ38OWnnw+7ra
Zp/iV5K+4NNpNGxyglRE+g5Oeo7znb+qln+ZGQrANdM1KU/E6mJ+NmgCqYNMSsf3
OnSHv4wch9GQcdDggB8cRC4MYRISUKVIxTPS7hCn4XVmtCwt0Qn43+F9qhy3Rdgz
dcAlhY4+lieR8+6SOZ/P3qGi0lFVmNa5zFjmBd4zt1dl/fbJ+0WHF7oL7WfE7zNT
5oO8VQIHDY52Ro0q+DdqeQ4tr8RrBI8keS2PyEbU98V9bvWYvkMIYnvrgh9KpSWB
IHL9M4A67vfUL69VCHGX7QIHgfE9KS/1E25YMCF5pcA7/RVoeVZu9k4u2B5uxjUn
oafFYcKYb8tVHImtgwkdw6Y6JnCnCj/riDwBaNMKdn1gH5qQkNnx3blYvY5sSlpK
Q38ejNlY26vnDJ9pSB65PZ7SajNJzVFAsCuG6FqfA90NvPQ6HxvwqNy12Ja5NXve
DDdFyhwPFuAmsyEA0O2fsRFgMisXrAPKX+9IzvjQFQIeUgLkF7AwLp4/H+X9YDGH
9EXMu9YUwFJx4F6m6pvUFYY1gWMiB7qE4531+JykcxNG7mQIkznpD1pcpFDxPzOP
tiXwYWwY41OzTqmJMlGEfugXPxmjsWgZs+me6O9xbivIMRtCX0eNlZtQOY/5Tbtb
HvoS7CRJezOPD3zWKo2iK9IQzhDQgED1ToIOT/ZueX6xewRwu454Hhv9A+2J5T64
8lDHFs6/+Qp8tzSdKc7xNI4PZ8snSWVQKBOUtjHqcDHcVsPLaRPbhNAR0YUzoti/
iIQcvdBvGzD8uembFf95/GBUTBwxxZIhTcefo3SrYQZcZAQj2QaDG/SZ+yUDwasi
Z7wxyqCPD9dYseyhUYJ6hwW12saIJPvTAve/O5a4AsWVfWcpMKusUA4eeBs16V/r
AyBKRy9/SW1eDIojMhu20v7Cgsm9M1iD6gcAOJSV1HguQPu3TpHEora/2btzuN9O
+cbkbSiLF2B35oJWD4NgIaOcdOSgXtxQorJPICf36V54Y8iLczLlTECrrdG8BP+i
n3ZjGiUcZHX9z9dGJo5RZG4bdqmdarZjzq7fI9y515BDQwxl4Kj0i6YlHSGfqd+y
gFPcwXKoiJ7WlM+HjOgNn7p9dS2r4FalxFb7rQrxgs401WIBbXtKYUYIRA/A5eo9
uyR0uY5LbsexqAK4PW25PjskXi/8Zr0t1zY2xf6a3Gt43g2p1NXQai9ThyPuzJia
Oniw8x+K3aYKmqRvxpKM7nDuihfGJV3FnxfDcQWGGBHA/woNfRGM6a8xqbaXGtyE
qL8OaQw6VsBnfYJ3aKDCQz94Z5bdFfcPNqFHeYus85FMyx2tqZUnhmgc95uKLuhJ
g+t63MSetDsZl15xJr/uJqfHyWrkYV3GaKo3A10iIF616o7mq3CcU+16/R1Zby6z
t3HEp+NqyQEzuDN/kSLrWYvyLf5zSmUJMGak0mz0QC4K3jYIfMGNvtIQRlam+yuJ
CSKjf2DX1bwKZ/kuHEgU2zEaswBjpj2u1S/SIddLiXRlcpxuSA/LFWQxfdO+S54A
vxHY1lLXtLhDqT408RD3rbSgoI+RuZPg3PnCLF3qpE1pF5A3cDUJTM3bC8GCuK5g
DKvycwbeGqSh2O4Q8ii8YpgDKskx88vmfCrLo57QDedAgVInDjYTSOrzQmoyEYuY
XOsgAdSz5kgBZBkgpr3OP6Dr7lpwmYfFFYkquY/G1/fremxsa+VYlqsnY29umfCx
xqaYMl9pZ1RyDCvDvXfIPclgUNUX/GOYKzTdRqbsP27JwbjUo2OtnZFmETAOh4sW
VyXokoG0YMKQZP/U+41j00D7Nu0/YeZVziILkIW9PYe/9uYmafwkiZy0MyUTHwkI
ITLPmtlNScneAZPhXixRbD0QitaPELw0UNxvfjXyLvXbTvYsxSfIVecK2bBHSLcA
lOpesVv2pbGJaPSntLcWwZj7seVkvFFDwQ7mY6DnqIin05z1zyvc4WRsPPKCWOZy
OBOnrorsaGT2xeY4lNIsOAnbszER+xJb4IRrDA6uoRRNpBvJ2DdZw6IyGF3xFSU0
EiTjBW4ppKhOcgSSm7iQVhi0rBf42ljLyqDNGgdYNrl0ntTw6HnbOlpGBbeS9GqF
Oy7dFIA8KdQScSVY88Ndqfivplpw2hmkutWOp3edJrKfBcIYtqn/Dbw3+DAhrt4A
tQ2AETdK2AJ02X44Dwj0gznuU4zoCi0rjJKKLSrfL8plOUsWSJh0PXM8oNjOini3
gqRIq9ocvQXfTICNYpWSIRpdMQLcQ+uEHANT3QM0gHiBhTd5couxSHhQb1KH3Xm8
GPMoBKCgWp0iopQXIxazYXNSndXX7mpRfduMBoRQ1PTOLgH/TdkMyxKNhvE0kKt9
krNWGopFwb7ELxZqMCjrpgg8ThQMYL4tr7hIFdOkpmA6myPLxTBa6MleWU9PFrqu
lScgMCpok4GYbQPUCVrDlAvIJAuZaLXGid/PCkb5myIbZcgLwJQJqBXi9qKaZI95
tVx6C0Nu16MGw/DCnkCIQoUZ0430EML9AbQSLZWemxhExa599WsLuwQvusmCON4l
0wDJgSHPBCNTsYa5xa5zwTYb0+idaR+QshvkmGk36pKMKg48hOI406EPUPzkcbt3
4aLVO+BfarAMehkkA89ksz2edgIkX92k3Wwr7cevT8KAsempMV3RP2+RuNJpvQ3r
LxLKd8s7h5t8DX35Le5bmnrmnNEcPCvovNyGtyFOvlcX6ZRR0LMCJuaPFVUXLzJ5
Db3QAFVovr61mSQCxPnOPwG/Ba0LPo1SD45kUE2sw3H80jvohpPgYX4iAN/EknuL
3dfom+bpDg247t/CIMhxk6Hk0Nb47oN6dNO+4edVFNPgWs+Kcxmy2fwCc9Se+7MF
39E9CBnPQACw8fZQq8BhAqEjJzQEPnnz+NOT6DkYvrj7hKXmnvGv5M2g6pof2qVN
wOCJMU7YNfS+Q/l8bXMKo6Re3+I8pp9LqTgnNxxvWvVvHZP64Yb4m6RaVqrWby8M
E+4c4Rp4lmlFRWq7nhrzvCcbKJ6rCxtDq2qLi7h9oWMDTXx/l/RTSPXtJmrDgB3r
gwHD2PQMavv0FxPAzkkU6hitT42eQJ2iqx09uLRsVv7k68kOkG6mWlBhYc/SQphX
S4zDERXXWeDEXsBHnGmS0DJv+mnpDbS3xHeCQ8/cYS7Qd580EDNiN2xlP+MhUw9k
bj1kzETtVgsYMpFbABjOkiD4wX7ZcPQbmhAAimmouJ+9LCOcO0KR+2s6NnfGcWEM
ViSESIfHWdV0EwwMdsCltbKQoQpCvEXZvdEGxaCoCe0VFlD8mDIyuGz/uaSyHGcI
b2yuTcVhtwOMUwzg77RDLWUuzQ3fdlL5TzionPxg09/fzeV5UFJYVC6xcR0S/t6x
pu+rs6B4oCxLlqqvYbjwXAH4B2LKH+DDUhlJ6fJG2EcjPJnBZm2mnflis9hd7syr
gMlyDvnfaAfyIhluQIEKbnWHT0minPNoC80FOn3jUQ5z7JWKU6N23UewhmVDAMYS
koF8LCheEuMDLMERRqhGjcOjTCAO6ZWXaNZfku3Yq01HJkhu5NMuXk3wAQ80LA/e
V8vLIBFxl20S5rksaCUFnuthCzXup2D43dqmrEfeyTe1WbapNjG3pQ061LOiBgxX
R+AyHzp0rJ1l7T/XIE2zvFmp1IovrkQqZyM2zU7xson02U+6VSpIGPUUvBWkwEUe
+ORBI0EpxBgWKXbsXGWpnW04I3z1ga99KJFDFsViylFytgy85mhpNK3drmYx/f1s
7jLfW3jMpcb/Rbi/eqCWogQIAuyeywdBMMhq2NUKUIwztTOI/ERxE7BMRkgon3Yy
CALuJfLeltRMfiEmjv1+b/EsVwf5vAYyH0019m1oUoBbah/Fln+36YI/LDGzxiRF
nWeYtIvpdwIvJ3bIBupqhQRzAtQFEwnMlIFxD4/CE3OoaqUMd51tw7O7kD2q9zsp
RssJyRhkyzaLZcFbJQVfIm27UKgwS2F3W0k2n8kJ4z5HLq9n7/ZHVHYAPXntJ5ZY
0Ww6/aiQbyeuqBS1xwL3GXCyWoQ1QJ2y5YjARO+yrjsgJbdmnH7BUislCK+iF2vK
N/xR1yxfPiidKocW94tAZIcYRNKUOpa8vP8ZUDTi9yPEmk3QHrDXONeLsHPHOAPp
uZhrFJ8bs6jktaO2tmCM3WrjRm3LT/xa49KvYl5aqx0R2Lh3xRhlrd/O+DFIu8MQ
HVK22/u9CR6vyboMTI+5gkrvm87+DgJuDjUojS2n2W5us/MYBwKZEPVGpFnBUrG4
wqoDKB7CcKz6Z+YUV26aVPXPJAJ+2vSq3oE9MOI8GUlEhz96WOSyW7DfRj8Fhahb
j3X5YdInvWMSIh5o+yO2WL+Hjx6MOimbLM2amXgphmzccO14WoI8hEe3TZVHYxqS
tVqDr2t76zrmb7/oV2aPyT/VdYxwOhArGYXbqDHQvYy0InBfatX/fOActMXChYKQ
SP//kzfKnhWuFRSNX2gVE6QLfane6gyiB3cdaCfuKJcqBWSKK3RyWsFf/GNZChuj
HMep51CJdYNiYGuFv7PVypgXa8z/zr3AOMjUZrq3zDRougl41KczuIhpi0kDA8fl
ZBdH8F83qt0XadDpPkvQZIRKdUTIVvS8CZ8k35LHjv0EYNiBzqeNHrllAU4UKWnA
O5Ov6yYWLVdqgk+bxsysIwGJVI87LHFN1AAdZT+0AFzR5xeQH/pDiNG04h5cnVyz
iGxrSlks6hdFrpkC70NZlIWv3UXCmjM7c/SyRu2p3PCN0kfhwR9EoPARWSSlbOtm
XetpCp7CSqReT6sMj28xSUgaH1t8/IIMwbKbQk+1y3y/k2H7/QcfiA9I/Qt+qets
UqsIeaQw13tFdb1A32kFED2LCVjsc032tS6kkNsnEoep2FHMxSn0bNvLV7H1u781
QlP8LS8uTqWT2qhLW0W4pJY6a3SFqP4wAoKHUYd8HCmzcuIaoyITxYSmkHS7952E
F3w3HuaXDbofzIbq9OSwfZ1XPbaZZOTi6Wk2wdKlHwZtb/6NnnGZ0XfdIWxjKgJh
VFT4LW3/Ip0iooC4OrKzIZc+NKU6MUk/EoAGlMCgfh7Is7PfucmSSOM25zjSp254
rScxsT4FEA1fVTGlFDq9VCkL2dp84aQVNqBUOB+UUfL6uMkfL6BqziFAvt6CYnny
EtACCdP9gkBrQ+R5ZAXjNQ5Ku/mJD9HMWcGWZlGPntxamT3yZm3okZtoswRK85DY
4os87I6ukQhgd+1gXdtuasmD9bpINzzidqejcDhuEtWhhs3FGNZWnVWNYElRR4WO
lclMXfcmVtIvFGwEX4T66syB28HdCcL8p353b1O+++jlQ06CK293MbMnHEc0freZ
TEegmUDwrbC1ZGlPVFAh+ZNqjrko0y89eLm0L2+qTM9JleTJG/EUQuOZPemsCkxP
KEV3JVkx84lOBlTca/3UVTC/k009a6W7id2R8hd7zOh3noiCPsNA+Jb+tALxdgKh
7VNSsX6r1mft5c0f5fxs1Oftc98t1dyvD5tzHRYRyzLeyPiLDjbC1zEhxC1A0w4o
4pdOs4khtRSNY0nVLq4Ks8xEE/cdEFXVpRv9ZNtePGAM23oXE5ic5HbI+jyG2V9J
jDyGbzYozwvo8bfi7qtNL7tPGuFoRLmzTQ5sxAZe0aWMHeyhg+q5lDwxW0qUk29P
fqI2QWjDsjJTvhFpPvIqbZvN9wh/G0GpsEJVTh03x8YAc2UwViBE449wjsH8g7cC
PZ5ZVWRvyzADnWtPMLMef9B/n5GwMWw6/nQlMXZfKTdeNNMRWMmcHnH10KQygCWi
5aGuuIcog1vyL6KWFNmETg==
`pragma protect end_protected
