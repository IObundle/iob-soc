`timescale 1ns / 1ps

`include "system.vh"
`include "axi.vh"

module top_system
  (
   input         c0_sys_clk_clk_p,
   input         c0_sys_clk_clk_n,
   input         reset,

   // uart
   output        uart_txd,
   input         uart_rxd,

`ifdef USE_DDR
   output        c0_ddr4_act_n,
   output [16:0] c0_ddr4_adr,
   output [1:0]  c0_ddr4_ba,
   output [0:0]  c0_ddr4_bg,
   output [0:0]  c0_ddr4_cke,
   output [0:0]  c0_ddr4_odt,
   output [0:0]  c0_ddr4_cs_n,
   output [0:0]  c0_ddr4_ck_t,
   output [0:0]  c0_ddr4_ck_c,
   output        c0_ddr4_reset_n,
   inout [3:0]   c0_ddr4_dm_dbi_n,
   inout [31:0]  c0_ddr4_dq,
   inout [3:0]   c0_ddr4_dqs_c,
   inout [3:0]   c0_ddr4_dqs_t,
`endif

   // ethernet
   output        ENET_RESETN,
   input         ENET_RX_CLK,

   output        ENET_GTX_CLK,
   input         ENET_RX_D0,
   input         ENET_RX_D1,
   input         ENET_RX_D2,
   input         ENET_RX_D3,
   input         ENET_RX_DV,
   output        ENET_TX_D0,
   output        ENET_TX_D1,
   output        ENET_TX_D2,
   output        ENET_TX_D3,
   output        ENET_TX_EN,

   output        trap
   );

   //
   // UARTs mux
   //
   wire          uart_txd_int;
   wire          uart_rxd_int = uart_rxd;
   assign uart_txd = uart_txd_int;

   wire          tester_uart_txd, soc_uart_txd;
   wire          tester_uart_rxd, soc_uart_rxd;

   wire          soc_uart_sel;

   // Output
   assign uart_txd_int = (soc_uart_sel)? soc_uart_txd: tester_uart_txd;

   // Inputs

   // UART tester
   assign tester_uart_rxd = (soc_uart_sel)? 1'b0: uart_rxd_int;

   // UART SoC
   assign soc_uart_rxd = (soc_uart_sel)? uart_rxd_int: 1'b0;

   // buffered eth clock
   wire          ETH_CLK;

   // PLL
   wire          locked;

   // MII
   wire [3:0]    TX_DATA;
   wire [3:0]    RX_DATA;

   assign {ENET_TX_D3, ENET_TX_D2, ENET_TX_D1, ENET_TX_D0} = TX_DATA;
   assign RX_DATA = {ENET_RX_D3, ENET_RX_D2, ENET_RX_D1, ENET_RX_D0};

   // eth clock
   IBUFG rxclk_buf
     (
      .I (ENET_RX_CLK),
      .O (ETH_CLK)
      );

   ODDRE1 ODDRE1_inst
     (
      .Q  (ENET_GTX_CLK),
      .C  (ETH_CLK),
      .D1 (1'b1),
      .D2 (1'b0),
      .SR (~ENET_RESETN)
      );

   assign locked = 1'b1;

`ifdef USE_DDR
   localparam AXI_ADDR_W=`DDR_ADDR_W;
   localparam AXI_DATA_W=`DATA_W;

   //
   // AXI INTERCONNECT
   //
                         
   // SYSTEM/SLAVE SIDE
   `AXI4_IF_WIRE(sys_);

   // DDR/MASTER SIDE
   `AXI4_IF_WIRE(ddr_);
`endif


   //
   // CLOCK MANAGEMENT
   //

   //system clock
   wire          sys_clk;
   
`ifdef USE_DDR
   wire          ddr_aclk;
`else 
   clock_wizard
     #(
       .OUTPUT_PER(10),
       .INPUT_PER(4)
       )
   clk_250_to_100_MHz
     (
      .clk_in1_p(c0_sys_clk_clk_p),
      .clk_in1_n(c0_sys_clk_clk_n),
      .clk_out1(sys_clk)
      );
`endif
   
   //ddr clock output from ddr ctrl 
 


   //   
   // RESET MANAGEMENT
   //

   //system reset
 
   wire          sys_rst;

`ifdef USE_DDR
   wire          init_calib_complete;
   wire          sys_rstn;

   assign sys_rst  = ~sys_rstn;
`else
   reg [15:0]    rst_cnt;
   reg           sys_rst_int;
   
   always @(posedge sys_clk, posedge reset)
     if(reset) begin
        sys_rst_int <= 1'b0;
        rst_cnt <= 16'hFFFF;
     end else begin 
        if(rst_cnt != 16'h0)
          rst_cnt <= rst_cnt - 1'b1;
        sys_rst_int <= (rst_cnt != 16'h0);
     end

   assign sys_rst = sys_rst_int;
   
`endif

`ifdef USE_DDR
   //AXI DDR side reset (ddr_arst) : generated by MIG itself
   wire          ddr_arstn;
   wire          ddr_ui_clk;
`endif
   

   //
   // DDR CONTROLLER
   //
                 
`ifdef USE_DDR   
   ddr4_0 ddr4_ram 
     (
      .sys_rst                (reset),
      .c0_sys_clk_p           (c0_sys_clk_clk_p),
      .c0_sys_clk_n           (c0_sys_clk_clk_n),

      .dbg_clk                (),
      .dbg_bus                (),
      
      //EXTERNAL SIDE
      .c0_ddr4_act_n          (c0_ddr4_act_n),
      .c0_ddr4_adr            (c0_ddr4_adr),
      .c0_ddr4_ba             (c0_ddr4_ba),
      .c0_ddr4_bg             (c0_ddr4_bg),
      .c0_ddr4_cke            (c0_ddr4_cke),
      .c0_ddr4_odt            (c0_ddr4_odt),
      .c0_ddr4_cs_n           (c0_ddr4_cs_n),
      .c0_ddr4_ck_t           (c0_ddr4_ck_t),
      .c0_ddr4_ck_c           (c0_ddr4_ck_c),
      .c0_ddr4_reset_n        (c0_ddr4_reset_n),
      .c0_ddr4_dm_dbi_n       (c0_ddr4_dm_dbi_n),
      .c0_ddr4_dq             (c0_ddr4_dq),
      .c0_ddr4_dqs_c          (c0_ddr4_dqs_c),
      .c0_ddr4_dqs_t          (c0_ddr4_dqs_t),
      .c0_init_calib_complete (init_calib_complete),
      
      //generated clocks and resets
      .c0_ddr4_ui_clk         (ddr_ui_clk),
      .c0_ddr4_ui_clk_sync_rst(ddr_ui_rst),
      .addn_ui_clkout1        (sys_clk),

      //USER AXI INTERFACE
      //address write 
      .c0_ddr4_aresetn        (ddr_arstn),
      `AXI4_IF_PORTMAP(c0_ddr4_s_, ddr_)
      );


   axi_interconnect_0 cache2ddr
     (
      .INTERCONNECT_ACLK     (ddr_ui_clk),
      .INTERCONNECT_ARESETN  (~(ddr_ui_rst | ~init_calib_complete)),
      
      //
      // SYSTEM SIDE
      //
      .S00_AXI_ARESET_OUT_N (sys_rstn),
      .S00_AXI_ACLK         (sys_clk),
      
      //Write address
      .S00_AXI_AWID         (sys_axi_awid),
      .S00_AXI_AWADDR       (sys_axi_awaddr),
      .S00_AXI_AWLEN        (sys_axi_awlen),
      .S00_AXI_AWSIZE       (sys_axi_awsize),
      .S00_AXI_AWBURST      (sys_axi_awburst),
      .S00_AXI_AWLOCK       (sys_axi_awlock),
      .S00_AXI_AWCACHE      (sys_axi_awcache),
      .S00_AXI_AWPROT       (sys_axi_awprot),
      .S00_AXI_AWQOS        (sys_axi_awqos),
      .S00_AXI_AWVALID      (sys_axi_awvalid),
      .S00_AXI_AWREADY      (sys_axi_awready),

      //Write data
      .S00_AXI_WDATA        (sys_axi_wdata),
      .S00_AXI_WSTRB        (sys_axi_wstrb),
      .S00_AXI_WLAST        (sys_axi_wlast),
      .S00_AXI_WVALID       (sys_axi_wvalid),
      .S00_AXI_WREADY       (sys_axi_wready),
      
      //Write response
      .S00_AXI_BID           (sys_axi_bid),
      .S00_AXI_BRESP         (sys_axi_bresp),
      .S00_AXI_BVALID        (sys_axi_bvalid),
      .S00_AXI_BREADY        (sys_axi_bready),
      
      //Read address
      .S00_AXI_ARID         (sys_axi_arid),
      .S00_AXI_ARADDR       (sys_axi_araddr),
      .S00_AXI_ARLEN        (sys_axi_arlen),
      .S00_AXI_ARSIZE       (sys_axi_arsize),
      .S00_AXI_ARBURST      (sys_axi_arburst),
      .S00_AXI_ARLOCK       (sys_axi_arlock),
      .S00_AXI_ARCACHE      (sys_axi_arcache),
      .S00_AXI_ARPROT       (sys_axi_arprot),
      .S00_AXI_ARQOS        (sys_axi_arqos),
      .S00_AXI_ARVALID      (sys_axi_arvalid),
      .S00_AXI_ARREADY      (sys_axi_arready),
      
      //Read data
      .S00_AXI_RID          (sys_axi_rid),
      .S00_AXI_RDATA        (sys_axi_rdata),
      .S00_AXI_RRESP        (sys_axi_rresp),
      .S00_AXI_RLAST        (sys_axi_rlast),
      .S00_AXI_RVALID       (sys_axi_rvalid),
      .S00_AXI_RREADY       (sys_axi_rready),
      //
      // DDR SIDE
      //

      .M00_AXI_ARESET_OUT_N  (ddr_arstn),
      .M00_AXI_ACLK          (ddr_ui_clk),
      
      //Write address
      .M00_AXI_AWID          (ddr_axi_awid),
      .M00_AXI_AWADDR        (ddr_axi_awaddr),
      .M00_AXI_AWLEN         (ddr_axi_awlen),
      .M00_AXI_AWSIZE        (ddr_axi_awsize),
      .M00_AXI_AWBURST       (ddr_axi_awburst),
      .M00_AXI_AWLOCK        (ddr_axi_awlock),
      .M00_AXI_AWCACHE       (ddr_axi_awcache),
      .M00_AXI_AWPROT        (ddr_axi_awprot),
      .M00_AXI_AWQOS         (ddr_axi_awqos),
      .M00_AXI_AWVALID       (ddr_axi_awvalid),
      .M00_AXI_AWREADY       (ddr_axi_awready),
      
      //Write data
      .M00_AXI_WDATA         (ddr_axi_wdata),
      .M00_AXI_WSTRB         (ddr_axi_wstrb),
      .M00_AXI_WLAST         (ddr_axi_wlast),
      .M00_AXI_WVALID        (ddr_axi_wvalid),
      .M00_AXI_WREADY        (ddr_axi_wready),
      
      //Write response
      .M00_AXI_BID           (ddr_axi_bid),
      .M00_AXI_BRESP         (ddr_axi_bresp),
      .M00_AXI_BVALID        (ddr_axi_bvalid),
      .M00_AXI_BREADY        (ddr_axi_bready),
      
      //Read address
      .M00_AXI_ARID         (ddr_axi_arid),
      .M00_AXI_ARADDR       (ddr_axi_araddr),
      .M00_AXI_ARLEN        (ddr_axi_arlen),
      .M00_AXI_ARSIZE       (ddr_axi_arsize),
      .M00_AXI_ARBURST      (ddr_axi_arburst),
      .M00_AXI_ARLOCK       (ddr_axi_arlock),
      .M00_AXI_ARCACHE      (ddr_axi_arcache),
      .M00_AXI_ARPROT       (ddr_axi_arprot),
      .M00_AXI_ARQOS        (ddr_axi_arqos),
      .M00_AXI_ARVALID      (ddr_axi_arvalid),
      .M00_AXI_ARREADY      (ddr_axi_arready),
      
      //Read data
      .M00_AXI_RID          (ddr_axi_rid),
      .M00_AXI_RDATA        (ddr_axi_rdata),
      .M00_AXI_RRESP        (ddr_axi_rresp),
      .M00_AXI_RLAST        (ddr_axi_rlast),
      .M00_AXI_RVALID       (ddr_axi_rvalid),
      .M00_AXI_RREADY       (ddr_axi_rready)
      );
`endif

   //
   // SYSTEM
   //
   system system 
     (
      .clk           (sys_clk),
      .reset         (sys_rst),
      .trap          (trap),

`ifdef USE_DDR
      `AXI4_IF_PORTMAP(, sys_),
      `AXI4_IF_PORTMAP(soc_, soc_),
`endif

      // UART
      .uart_txd      (tester_uart_txd),
      .uart_rxd      (tester_uart_rxd),
      .uart_rts      (),
      .uart_cts      (1'b1),

      // SoC UART
      .soc_uart_txd  (soc_uart_txd),
      .soc_uart_rxd  (soc_uart_rxd),
      .soc_uart_rts  (),
      .soc_uart_cts  (1'b1),

      // GPIO
      .gpio_r0       (),
      .gpio_r1       (),
      .gpio_r2       (),
      .gpio_r3       (soc_uart_sel),

      // ETHERNET
      // PHY
      .ETH_PHY_RESETN(ENET_RESETN),

      // PLL
      .PLL_LOCKED    (locked),

      // MII
      .RX_CLK        (ETH_CLK),
      .RX_DATA       (RX_DATA),
      .RX_DV         (ENET_RX_DV),
      .TX_CLK        (ETH_CLK),
      .TX_DATA       (TX_DATA),
      .TX_EN         (ENET_TX_EN)
      );

endmodule
