//empty file for now
