// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s13z1taFptYlLtp5GoMeV/BBipXUyHaXqSnnNt8amR6q0bM3/9USSeRV7HhYdcx2
w62E1RtlhN4dVBrnlPhukLLQABk33/Hw8WH609S6e1EhOmbF5aNaLsYForu6Fmlz
dvMZgvKjH9Vhs3j2WAwNbRck2BbXzirRpps1UffIgqw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 180736)
YRJGZMrDq7t5cUl/4GIYrl6U6+c0yaa1E+rOzFBF3TPRjaHD6lzX/3GsBhcY3uqN
B4GEJzJPD/FD7Yfg3ohNTyfMMTSfmJuA1o9aRVpKSetMNXu6uIDoRNiDOO31E7xt
ppOJOmQeAT9Uswql9tJhREp+g17BF6ZlzjjN+FECsrnHazB1s1brkhXHPBS6Za6/
kkkQQCQAhDWFmyFn4vGbxQ2Jc3YFeRVcSauw3KaEbkiJqCwjABkpK3/qRcptBIgM
DDr+RSCgYMYciJQ0miUGgpNSXpfkVCF//BzdUHkAcbCFKtdP/ARperNwew4uROii
fxJMnlbS484w3kz6BWB/+uHTd5KEEhoKXIB0N1KKJw59q/cL9omY+GDHuhudyHEk
0m8BpaJQ9hh8wNggwh+FHraLk1DDtLyUXW4GqA3kFaMVtIj6Do8b75dNB0l4iKPI
SJj+7/pzB+DCZMhaJt2R30nVuGwWfeMtrg0+XIJ9eI6suGvU46xiWLkBo1V5vg9Y
Gt7ZogAWi9reFG1pzEWNgR6ffsQ2bVD2H1MbsV4OWplgTTjKPI+wkjXHNjl/6EHo
TxhliRB0J0v21a6AqZgJ1Iln9rusWn+jnYKvwYTNAyWC9DswvjhzF3UcNYDl31EG
XbeDQY5SEHzJFxNC83aWA/cj/bs3jJ3xg7LWeBAyhv/M16sbEVrzNlkzQcaOo9MH
DspIFr6pJyi9E+X9P829vB2CyUXvybC6dV5GisVmC+x/a0oWF8LD/cfWCJa0+viq
vhVKJPEcTnHJGeA6xMJZI1cCsMW7Bh1gQO/UsXtfxZaM3lmp3yvM0Pgf92EsPl/+
HgnmveWMBuoLRcbDGLRu/IWDAlSbDs3m4fIRwXV2at25muqlGAcZG43z+qoKD4nB
A9g2d+IKInxkcsgkV4pPwo6ZrbLy2mHC9uWCtJ8I4kGzbPmVOZsV6xbzjBK6NwJY
NR5dxBV3eutB3p3+CcnidVNPOfuotNjzM/4Ihm4wVZ2zb3Nkm9D3G8659v1uwrVC
5YJG95smKcnemC/Mfamlm40z74qBa8/P7biJmnxQzzSziI47pK5/t202N3OzkNkO
hAUICDQmrCWMbz6w61ow9tSh2tpuaiCcnu/2pokoFIy0A2pG4arwv1MdN813nI49
uN6C+l8YqxS2E39rqLO/+lWFKKwW+jSLH4YSavQRosxsglEePk2TcYQcSS+KBWoz
3W1axp/zbcCjBwdxGl2hW84cXbjqpXvShNcvs7VXRbBohXECaIkYC7flzViHAKQj
8G9QFH+Ov6cMxWUBmLZSJ9XCnzed0Ro1Nlt97OeItjNG0g/z7J6WdkheQ/UEAH8Y
DjOeONFkaztA6IuxrGsG9iY38Ev0fbsdVLS7ZfiJSNmxFejIo+b9VJXBF+1d8MvV
QDoJNgA6hctrQH3DbfAqkM+MSPa1KNO3V8Nh6W/2YoFkw+76tuNMWLGCohx5w+7z
r/sN/dyyj7Ru6Hc/sDc+xDfaLDvsZhhkWX8uAN0C2xWNXfGdmvzpBwEo33BT8UMP
pief6KpFQNltj8v8XP5KGi99Dvjd92k/NBAOdtTNdvhFX9P0bNk/FpKmCB1+dY25
632GwXB/Q5pYFsu6eQHPkEDkgiiSSyP10Zpcs3Hc5XhFLOEDOD57D/t3ot7WEZr+
YCY9rm3rLxijp21l5BT5mOY+XmV515K+Pj+sHgQUGezdMpCkx+9Ir+6bbSfcs8xv
PC7LuU9CO+eI8gQ3AOlGocGREGvoVkSW2vqJnPXLxo2R1tU+d+5YdmR9ZbURV+E9
ScjMOYdKVsmUz89goYF4PzqedTjsFXYZ3AvNkds18iuxMMR13b9sklFH4thUpRID
55TIkl7ok3amqUYdmpiKeqvk2Ydirytsy00wzGky33rnJx1Ol3zVODbXenKX8vtV
ZRgrGyG6yGzXZgGpKpFe5PEBhYtAcYAqR399EneMn9p9L+7hCVPvOosB8aFeTjtn
uHpvpImKFEYp0m4+chGODFJ08BdXHghHa27BA/Zc+aV54j7fCQ4IjGaMvfzopEoa
R15qTHfl2n0pRV3llhE1H5jEqWM+KVooFfuKsCUlr2eBDQxyvtXhx7wnHk/1lzcN
H/Ptigs3yz3aLBZQn/KZoNNIr4rsVPP/MoZNXDiGAlKiGoHsxeU+zNmOnK0cGaAq
xMfmayrj3m/qnbD1y9DNO+cJ23LLtO5xAIWOqGRkjdkxtEkiXnLUvj7krZBUie0j
TJrXjuhP/DU2rt7QYIiEQUX2pD2FB2QVQJlW1z1roqJF9gf/4PJriypqGeLBmgbz
zt+Rqp4Y90py7PiMDWAxkYOf4Dz+a4oPcrlnDZ9D7SOlIFHiWrux/RWHE5ULBLmR
SogUgnZLociturVJMZdrIITpqPPpZLatPYnaCQDNA3KD2tu073UxwesIb4kXOasG
rGOdeVjyP1HCuoOgPYe3V2/7s5ER5PEyIBPk/+LYOHtnK4CIoRMWpMFKixl8r3D2
0BGxUosDFZRF1sVsByA7NhfhDNo8ZFxsNuoF9OV8qod30UEYt+eA62muixnjPZdW
wooRmB+sWlFs8yx5qY3j5XDm85boV8HPQ34xYD/wNaTVLRcOBtSEZTKiMEUNqbOa
dWt5XPJghQwIvQon+09x3M1xEOPrsOhrUUohA8ldXPSIBoPiBlJBiXZPtag2/koS
ytMer/nvr36KcWTQY76j9cMeSBCCkdi+X8U3eWYNREuDBPxmwYImScMlDcHvFyGA
H1Tea6fIcAXdQxavI3lJaSi4EDj+jlaQag/UqlG1QV3I3gGBROgUAb/GcgjrKtGU
RvLJ77BVR3aQiRtZ8ChVekgmQRn74+n8D47vZztvnDtSuPg7d+5FIOVGeFdWD1gz
csjOtNOMIjjshrhxtYsWUv91kDT40T+A0NV56tN7VXcLoTzuoRFt3Y7q7rwNKA8a
XFIxMdpE+uwn18IToqqRXEKBbHrNDr9T1R+m8xaciXyh28YYNo7SSQnHM3dWdQEU
WrPHbzWeeeDeTPmYp5x94b+yY7jkTVcAnvwCIYVR8FXyTSGGGtl7NYQ/6jfDzhSG
R2BaEu2ncGZf3J6KxTjs81EymCi0BmS2f2+Cmt0LHV7a8eIMZO8A7V9sRprdm1qv
iNa8QwlncDBKcwh0kxwGoPJN/CzUfQD4dzT5+y5M3zmE7dw20I4/Qj/jl0tMZPWQ
+soYmdp8wJ8QUJs5+ikDEQhRKctqWxwkM11ocyRl+qqWnYus8ebmLSoSMrTiNb4P
XwSYigyrhsu0I57d7WpZAQiIIUPLvF28HLZYR09VDGO8SwEEKBSGwJRFRIANVQER
SsZnDg37Mb0cViHbCLuRixR8saw/3nF+mGpeV4PAS2nQnKIgdYnjGAt6seeimXoY
waFsdQTiCFdVfRBsdnozew8sQkScl8z52GmtImlGfIScV3En6lhIQdlgtrRy62cr
OrL6IT9O4umdK8gBtRLh1kGUsR9Cv6wWrh40svLErp5Fiq3XKS0bGoD1bo/VokL5
I7U0v2xqYmV+RaggYjcYhLRzL4GCcdaE5FUlCKMZiqSDGfhyK5LsLtrvgs9E84hz
PBK0lQh3uwcdZgA67JgXA3QicCAXzOHRJNi/p2K+lFsVdhZ0PfFuLFQClpHHkJoY
b63JqUNz53R9J3ctz+ZaWqkbApmNYli1srsE00Dqk6mlhxK6CjIknkl76QUNjdSI
3VVQrU8f646ET+9vKZ22L/v2zstB8S2Ak4Ng9Zk3GsgFrrT9GWq79fZFvzjMl6/l
oNOGTXGu4gQ2msUXhDUVsMClCE2WVFJFR2hxQKppV2rQfz6mLPv3rwmhzq4+N2sC
a9/I1TngEQx+SScGohD6V69f52xog+TTx3mGvIIBToAeFXEKm7TP2KXP2VGYcLBl
Urybl5GNJ/2VWrdsAIfsExKZWkm+qity4g5SPP1pU0GFmBo5fVhbhnv+LSeD5c8O
W8O/2dKUPgF8QV9DJe+85ehJVQeA3uPa+OaMxKirhci8Ab6UEGma0S43LenEqDr6
nGlncOjHoMn/UJrJ6TDIZpRFCMvXHbbRnpw0JFFUxnbZRCfyXyKh12hX06xgWdGS
gvFDvTMO9d7Qu5lO4/Kpt+1UaJlEdadSIdQAW5R3b5Je4+iOqgN4Rser+evA4CWX
9hjou+43I1vc4KmbTyKeo8tZjK6c3oHb8DNEgffjTI3cLk+qOZtCjshsz6hrq81J
5eEgU9qqZQXyZ2oxpeBGXf5LquFWjF0cpj7FXiFJG6D+S56rnu3B7bQysHBvlRSR
vYqkYFgFNQUQ35qUbrlYiC508HsqUoGkNsQIoQNm1L8UfcSgHdiWW1ZKVUETM4AW
reS/eWd8CsV1Luai1erVozhL3klqfDkdHD2pEyPXOYRdUav4exrZbCDM8s2AG90g
/pwJnlgJartdxtAqGXVJG0o+KcKcIvRpam6Z5tGB1K9nkwy5dyTvwIdHNjVk1kQV
VAiPSYoY+LlbzmUlsdie+KNqIpD0z2kqSjXB2T+VZnD4zG2MvEoRaZsfUjHWQteg
S+3m+2RVm8tmqL7UefySaIZfEiHWuSLsEVPrT996ULoCLkoaqT4oXaNtvuiKphLb
t29WJ8zflE9cGF+zjB1l3n65qBjMOybroWsnDmYYoAdApWXzulSvU3i7DD0Q3wUV
q94m3XCtT/H/Kv+JJ2KCqS3LATfssXFDr9kIcjh+p5vJY3EidF0YDfqgsY+/p08E
2d9LB57/fY79K/IJbY2ccIq77YhglkSaBmWaUlgAD4ChfpoTcYcOuUIurTU2GfnG
7lg6TJCXq0LNpsfK4dyrYucxdkWmk1EQChAQJSd9SJ1bCt8shAgDTLjCXYYccNpt
e//cjD+R7Hd1+U9TDwWisUKAIx9pzMj8Rz0T14TNzI6WXIgAQWkVq4voq3Fa1XCe
6rVSzCwBxBFF3GE6HqBVsfVRmqKmUq0qTWztoYZejEsNIeOzeuxGE+cWri34hQmI
54T94wX1WrP1NY8lWGKenJ9yTdO7DBG8zgMYmPPpLz14dzKfvVnfFRiqT67zAG0x
dRSFcp1VFVrKsCw2fCVDoMtPeLQNruzJxlUK3t+xMXurCuVWoYXM627cq7mt7aYz
/BBaR/ChBFuvoHcaGstMDGMyCVUXiTfqVJa8kYEd/riwJYyEwV8W0QWhGWE4gm6W
VyIwAnK3w6SwNnS6nseOLa5g/NIRjVD1WmsCx2CbONMiAlZs9PXX+acXWTo0hsKk
OCFZgDxMIC15lHn9HHyf2gsqjlyeh8ena8X/dryBMe4MP1yZgphHnkbEUTkMA7ol
e8vwbPqEQjgGiNn/EVV/VoXmNn1rwTLdXzhD/hcB8ZzFprPpWDqN06HhS3JukALm
nt92htIhZK3jXDPrlcF5WlBME/vcJ7zEokxokiOkoyZywJBHScskVF+LiOGzmQ0c
u1RHcmCXPLSO/9lyYrrqEh8WpsEpPjI7dbJYSzCBVzdxgtk1oFhlY6aa2MKtt1/o
qBZFlg1M9+VUxf9DjHerulb0cQxtcHE6+Z8YP1BgQmDCnQGwHvs1ARjcG4BOyP6U
z7WoCp0hyj4zYBqz0EfrA4itnYQzr+kUGUFmDmBf8BT60lTKE3eh0rJKHAh09G+4
76XKn+CwMKo+Tb6tiYqtTA7c9Egu1/mlpFIfngKMhG0kZke2OzkuR/qosq0K8niV
7szJf38okTm1xxaUt4DXky+1wci3s/R5dt/V1JqPpuJ9T0RSEe7V6GJDHk7rtIwv
pCGrBpJzqusukI7sfROHQCs6MBYcBC9Y4ncmvQ80QUy3ArvPqt7u2WUD+nGyiXBK
Zfex1d3wRWB1vd71TcZOxfqS8w6B7PWGOZ3KN1vBhECGrjUa5FzdX/SJ9nad/xio
08smUQHIE6Ts6+8RSNwXi5wcFIc5XuX/9H850cRhA35DEYNo2f4aVx3bSWrmACf2
gV/EeR3f9syO98Ttj+qC/cYEjxvzX8w4zp9gzYF8A6PMORN0zlgHnhhd+ZIn2Kv1
JCDpVNH0foj/91npatCwHmfslIl1pvPXRC5+7VgRlIgvRG4zz7haPmTS5ZALNmqH
K/+9tU4BVYybshQo9R6LRVtaHahlD+Tlx5GRlMsvl8HIH/AE0RxE6hQQbs67+WC4
aErSFVkDGnbuUYWDsYVExtU9cimhRIpkmnpTw0LiZaqVfdmXv9nSB2qtUTsHaf3T
ARgrgEZOqBAYQ6j3E7+IKSCum0O2/MGHkTyaRuvax2FwolybPukvk2dfyrGSoG6U
uCEfoguZJ/4xlKPumVfcAbkbqujmmvcO8PKmtGzJjV5EKAolURqDiAN7uNh8WTLM
R0mUaHDuiJtOtkgRig8Beu6TR4T/u0ifp5jMJRVYX8w4w14FK7oGBh4urBYJA/6C
Htn5KO8MFCtfQ/V46Bw3m5pW9jIVnGsc0sYwlPubUoE2XqL0Hi1n2JTb5Oxn4799
+9FexAynHwevZ5CIKiyx2IPyrF5UVVPRttUbWna2aJoAm8W37q91SASGehfudv6v
Y7pG3Be4/ki+jxqs7HLqQme+w/hMivgqByz7HJ0qQn+gBQwSEIIbHD4o50SQiuw4
eGJy+bxm+Pb+DWk8fcyGpGifnf3eSaMSIZ7coqDRjPSGH2H2I2xsLpsE/p7Dow2g
Ymbr31/CaV0j1kClOfZm1U/O1K8BdbH3hLbFDvc+rbTZnQZp/60Yo0iZmoxXTr5t
BuMNOhAIsg80HPBhSfzjKkif/6KBEks9+enHizG9dujEtcygVWmL1VMuEG55XxvL
VR/8VI69yMsfI2UtPV7YGkuSLvhviuK6KIOc3jRzMuY3iNJR5gwr7WPICoOv2WXN
JeT/ESHM0b9w+hdFAl4ScGWxrEJU88bjHhbU4mRISX0aYBw+ad3yBMlJRw6vhGIL
+vOFqB3JOPEwerZPirRqhuATapx4VZ0RuTxzcWLzmq1k6ZBJQOP1z54e0GP5JLmU
KODwgNWLUuHN7C0zcG4Q4eQuIJu5wp2YaGT+vbHoleuY/TkNpVV2kK99HCELYBIZ
W12UpAViZ+O8mEobhQQHXuEMfYHIVMORWEQbs6yFIvCTIYKt78ojJMkYbBbw1daV
XxrpUcWucraXr7jkDRys3xHQxvUG5aAaxum93DP9enP8bBTVGLUKwx1e8MP6MqBM
5OTTwil2kEYrHdGla55nh3XjKH07r8jZjaGAeDnnW11ABmHKaftCniI8rOZJ7pLq
wjeKLTBnuO7X+yQzJtKjTXEodj5mpzfCYsWIdB3nIkX1S05AzVi0AYQa8AE9J8QA
kDA5HlBXOBOX8CTvDCe9z0UIMKJC+vm8MRCZZYyhHlT4lCeBW6M+G8h9qVEp7gor
SclQD7D4aidTn6Fl/SsP7rYhK2/wAb5eW6QW0Rai7pevMq71/Y1ch+2gysMbE37q
Cbtu72nvMEJ9zqy+YILRJ8f5yi3ftmXrPlfliKSjLJushU27yltT4tqd+dA1g+kL
Mxql0fOtnjU2lhjcLplHJSrYU3MOy/sIH/77b/2w/cHx8H/nNPbkIakWM6LfJzQ1
HEYQrfIvEaehBHuVlB1VDA5rfy9WW4lVC5bxb/XPnWLYWUI/UFiYdRL6trdWY/tc
3G7tvVD2UVyjF9nZdZEY+AH8VXvXQmfk86K5VT56vAci2Pj/RUUnsN7/K2H9a2Jz
DdbZK70NKuYM0q0J+y4sJjJKk+xciF91xHHEfQp8ZeGfvw5DhBRvjx39TsLh98w1
1kT6qqPTOa+CDid/3pvDQshVHAfT9aGU2u4G4H3hI+2ggJcSqJOeKD0FSEoKmLAq
UQtyDN8XmStWKTsPVD9pK5SzQ5GMNdsnwTkfFQiSuTk0EcVdEMzJ8Rz+ht7c+SJB
vO+mAVk8lM6yZAlb0nczkIrEm/DCpuFjFNT27fzzBjL+0thic80ktASdy+9pBdk3
3/DXn3JdcjHN7ea3rDf2mEf4RvH7UGyaVE9aCTldHjvUyoy1ou3WA/jrd+JRlXLu
tKwFa/ckiiO5IWDuh8WnoAKzi5NWnoouINNA1PxzBiviUksIJZrB8PbTnZEm2PtU
aF6jTUeTDLqop/cC/BbQVcIrMD31sLcgdwIOgh1imQEDHURIxB7unybLdMT+v815
R4LzgcBbjQVNC3bmY1w+uRej4EU0nm1a4zAgv8615+ajDAzwmGCzltKeY5Qsfi5f
tgrX1qe3mC+EapYuDBRHP33rQH9zylKlko0VncOgjiqb7qPJb4UjgxzQh1oEtZWo
0+sA85BsHFQ2R4is580Azik6G2/uZ8aX8JbqeHlQtAKxJCC8/IVepCT545UizpK1
lLBL0RgRPMLwIZTdQlWWVWOWOY3HKsDcrmXvpxMGxyCOkoUKFKK0DZv1YHDLbHVV
VNeV8Bd4zZALXEAnfxQRu2Fwckk5ekV+IWJvfA+XZbI/8gJk5ayb42GEdnTfcngK
w8vdn6rlLv3ukazYGRJMBpz1bG9r3rK5CTNF3qsGZnc1TbfmWsfjb6ERKKbd0gR1
37NFHtX5mkgNwSYNfiuLWYoM4s2iQl02QgfZzRDsS06pJp3dwTt6dhWl1gStI5PQ
NEaY/j0VcHeonykGOGS0Zpw0EkvD5d2IGP8yellsWWIVbWa7ijKCZ+yRkc5+q0NT
6XnVq0XZ9oGhSn0l8vzoKNd1hdekYXw+0+R9tKOkQlH/wFapRRiTKnAJ8Zgvt4z7
2cjKw04+qvuu4+fyYJMP3O6RaU0HqIUBpUXZxIsd0XgnnzRRqN+7bRLmJkE2i9fb
LODaMnLFS8b8BDkTS6gOGPmnlfKi35USclCpQt3I5wJEt1SDuifjdNeMiCzs5Eo1
R3Han84rjMuqZ0YNI6GqYKP7LhV8HX9+3ALVCDKkyeaDnxujyRoag1U2C13Jj04s
lB8yuvH4iDLB5br+J+5WRUMxqnEfryrrk5NrUk3Lz6WhfEjzsTPjNz4BaAFysVe1
SB91HPNgcTgfNTOfVVKBph0hf/hgABMIEQaW44nQR82cH2/Lsav81Ks7pGIqaBLX
bzkPez2zieziSd6R0ZRPJskpyGhhx/7DqI2XEI8GdWRTC3uOvqi0qmnsokgPNOZn
vBtGqAK4X+4ljo7nE0G7iV6vswel1NO79rYsziYFQX4ST7bUgF6u1Tsegl5eJdoC
XbCbIaeAC6p4pmkELETlVY62cR/NuFzctEe4wp7N8Hd0XPLCtGltKuXqbL2GPNA0
jliUqLIkjbDO5Xygke78Rcr5oBCdwYafqDVx/7ZyF8n4uY+LIdnzdgEqghz3DXPe
rApp0w3SQT5DJc3oQgdWpHAg8IP4wMrFfko1scElc2P2MJNQc4RiaSIQRNSo1Sgq
nrNylvqyWMY1VxN6V4Qy3P7tGImj0H1Vo1JiQDjAnvhKUqdn75Vj9gm52FnGvGkR
+9tW/UsS9PX/qHH9S5ShCnV+T57YpaPb8JJwJGsarf+3x4EUYBDKLPNVnoGbwhuj
iixnXoSCMNj4lFk1Oy1kLwcl3C4Gp4eLbZbCZn9P3+ATSWNyYqd18ZpGdgKpJXEX
q84Dx1i+wJYE0Wq07aoENINVjFTFiSoCt3/ukTgTborcm+SC8nNJo6xaf2y3xp9V
e9D3USypnX1uzW5gduWtRycOHdEgENDDPv5RQYH197ZKvWCQzmm1tBrC5NsGnxMB
RHyRK2jrHLwJkllde6nOPVtrT1uatlI7MttizwcDhhoYMkfd0PC9v9cz4ArP9M5Q
GmDoSXeH661i8guKlnPeBe0mQ0Myce5DeqEp7Sks4xXNpK1WTRQi2AHCeAb0TERt
jnuoIOvCV6CHxqar7Qr2pa1lcPIAHER/QSEXtqtDHsfPgdgzBhJRADqAyL7Xr5Ma
S1Pi2zDS8ZcD9uIeq651xEPuBJnaqqEd4GQpkj6uYK5/RbQnWRPwWZ5XBmv6QJ+p
8fPgtG8DQCwejQxmIXUVnkOqtQuzk8AQeMK4DSzKO40yQ2fpzDaR6ZgyuPVVfRCl
PLspFZoMXOHEDj6t0rKkvXkMj0hS3gaLqGS9sgdaLaii+VW/QXS1dHiGDHynLQOu
6tmIpol2ulySIe8aC76w+NQvYM+03nWg97UeBaAsGdazyuhfMtqJbcMnBCscaaNX
r4Ct6F5lHeorOtSl13PTMo8Hr1Dov8iXgkphGLRzmtU2Jqpd9a5pfKa+8jydahA1
HkPcH5jgMKFiKCbKHQoeGMxZAlPsp2Ihn68zaqu9fcBl4mSYB8c6MCmTUQLc5/J0
3YsdQu3DZpzEbEejG82P6eO5MVtjs57I8xpa0n1AMha04VLK9Ys75jrjgqlmVDzv
9y2uB3CguIfwadLaEXe1+S4ZFP71BRRsMqN7duve2adkiHZUC6iChQYvREsfdL5i
HcADCR7dCb81vTt+c1F96lLt5hOk9LtgbMwVdj1Gr3mZdbikwMeGf4JBeW6A+W0n
Jp+ulR13bBlwSG9Foa2eTBzdvjn735JPP9LZu/9lfwDMMhsgtGqCO1XRGMDhmIOb
Uxqp4YZu+AmSWgKza2TnCgAKeRe485t0J4wymARC08Eq264OVH+5NgBHUtJkEovG
N+sBxyceuKarZyB8XM1KB1FbElX7G0UohEx6+WvOKxjAlLeS4TKouvO45E/AKMdc
YWik3P3Q29TkiOqI4fnX68b/d2+trtdViNKu6IjAUcJI0CGdsnpqHFHZRt1pOxC6
ppleEb4e8LiVtYujNSzK8CfYAmc/43bLHqTonGJ1expZlisXB40t2O8zhn9tc9v5
nvMP1rroK3WmMxTwmOpo4lGwExUYlEWaSWlxoo8a+kvf5baaOsSnmlmv2RR4fvYU
RJQKIQrY8WvjdRUdfAt+RWAQp1uAxKL9ktdf8M9cLo+lOvbAq4Pp0NqJDMEDv+4H
L1C15idYG7d9l4BLsDLPkN6XVOTNMJ8C13JznWJsL56NaYGqZhIA4vHNJpkHCp99
iUOR0CPKwmhpxg2xNI9NP5tilQYX4Xbu6TA8dvxtZhJaMDCtpLGZCsY4BVohq5ja
Fa04vXgX67/5GeoExvKtNpFwMRJiVTjnfYORzIhKWBsndFKZBVVbH3PoXxJQKFBW
Da3OoFZdXOwj7Y1r4RURnayyaZQqE3rqu9Bs8cNYU3jl0OJW44aZEE9qUL0VrfZj
AkO5gacLP/JG5jt1hbYj9VbW6mPanECltizNydGLeQrRe3JsHuFYdF4ZTQBJtPpY
7T/CoKG1sBTjt/j/0f/I89rI2UeVUbM9Gc0qz3b/ZoiWYVufD1lofizI1BEX17Sz
SQCKzSzWqvT+7cF7SwOIm58/6D/yMwXtnBnNo8wDDsZXkR8jY3yfksAbvtcb9NYO
EIAyxLC4g7NGnz25xPLeRntoR72WgJJpBuc5jd+88wnCkx2sKgXlL4Uf71QZkb8B
ydsw26xDkF4xU3L+nxL1OXS1Vow9H/T33RS+E9oDlLNmR7TFvTSiWfdVEatAiwlo
tOfaWQ29Eh+nvLqWhq/wu3XuXAH3bQiS2Al0EYCL3/+aa8i/Dzy/04glQG2Dpc2n
uq0EEF4P0QJPdO1S5Qv9LKPyPdON+GdHh/ISkJbO/unVgp3JxpCXN4j2ebRefClE
Fijptw3tBjmUsmnHFROk5vxgLfIioaMDCjs00ZGXtpH1+WanwE0HMMFpSrxb1zjP
G953tyeE4Fxi/gLVnzc6Pt8whvcMKtMSrQcdwDYMMJ2EMcqhBjrswfqZ+OaTdDpP
sKatLQdQgeBgYwVORZZGOy4dwvR04ybv3ffIvx+HjBYRzmjc6m0DcnJ9T9KP3NqG
vx4lIH755xif6dck7Rv4ia2aydJMmZCJkMm8tyhE5v6GyrDNOc0uJVJM3Fom5Tdp
irXAx+r+pRFuC/C2iO9EXTWTeF4wEMOB4eaCwm5xzvToO8kFSihdP708SjRo/sUf
LC4TbFPmo/f2gqTRcmyV7c3nxCpBi+IKrdcnYPrPBYNbMyCv0uluR8fJlWMu58hf
31nZbB6E5n4QoS9wdj5JYc4eRk+BhP98lh3HtycW3C9OVyGcehAbMhGvq2SM9yqt
GqOi1LRnyMZG/dlrwwrmE+KrgiTCEhO/4YWnN8Mo0fYUXH8rOGSU4uH47U4fRCl9
G3NH7oHPm2rX0hmo0G/IyBJc0cqDHPP6RB9esu1XjBuf+bZyH/MDl17Qh4uA7xCq
qZy22axn0HSOFzz+5Yi+MUWeVzm6mZQjtprWPA7O2dzrz3fzue2xbATzS0waQ9me
/MeCVksDGjOvOgUvgUF3aGZAvGSvxtNYCKoFS22Y+wopuPwlv2TvUjarcvc1ZhFo
SZnX6dvHf3cwend4dvDoTOwF0Bs4TY6ax5I4gykhhaCrnkdEDTD+4lQy+c2km2Hc
ekodKHqIClyvzBLRE+5fLSccYDKTlODcbU0uUV2pfAw+iEiEU0RoPRbSKgBieoBJ
YbloXQK8fED0BV8RrNBCt9TwmvqLrqFdAmNyli3eIookyQnV6kMDGWgIiGv4nNKD
evdORcqnkrQK765WY4eDcXWnVi1U8GwHOz4vN94Htk2W4jL/tXTgfdTNzgdBJjKV
IzFc0o4sFHlSkp0MkfAmcRLQtxMmti1Jvn0PEEbcrLLm7yHjcad+PrjCihVVcRUp
yWBuDTmkHNhy5oB0FMcMvSi44I8IG3mII0hD4otljYBDWZgkqPXoSs6aNULvraO3
8EyiPLnJ/RiURorJxi+SXcXR0SqSNF8oUa0IEQQgakuyKzEXGhXySf05PG1hdKOr
8JWOrEYTr2ps7VDJaKgqYCpH+3yCJo/o3lmnTNUyE68DCuy7ESNxDg+EQTqbxmuv
lit8K5m+gz/NG5/gDtjd9kmh8R9/9lEAY9OjzJsxUcnkhBPy/6Ow4gDJ3J5UM/IT
Dsbi9otvl9prU5egIl2QiS5RbYSdumjsfqMpZ31eKoH3dGFTeezuW6UI4NzsvHQ+
kmDLeZOFc4O94HqPWbysXS8254DelA1J4Zi6oFZNnxiYXoP5/rokq3yZF/NqB+YS
v3XF/EtlrhzL+112pos7Hnu1QVC+GKqTAnAJcUvOLGWtHNOrpEzdMy8FxyprTwz4
W955RvleEc7ZdGLIpPiDuaM4ZwSEJ28shB07sNyl3TWdz4RycJGEv6LcjTeL2IX+
d/lIK8icJym4DvWk1td1+aATsOj0E0ZYy6gKWL1ce/YwguvdZXGycrUOnZ1jlG2E
6GCnvVEYhCyjavN1br+YjwPpvNnGu5JnjrpnDmLyxYg4YL1Uv3U6Jsq/gvgHKOhH
GJut25Vldn3COxMqQbVg5n4QE9pDY9ftBlMJps8spXywZVJGa2fuWQ+Iw7cXzFse
rfzRv710b8GcosYASEDTOMkyoh8MuxYJoT/DY9p/VoJYpGJCgDEeF0oXMZ3ZcLKa
+Q/bNRWaFoDaYhDu8VbeoCk7YlnPGjtzZ0xMiKmpTSeRJsjWIQ0TNl0tpL2eZcaV
zI+EBBe1L3URkaDnVdgfmvAO1s7sV4hZBq5UKxNhxir5gW+HwLD3YTc4DooVeXi4
M7Duq/OgQLVmqfnuS64xEgFogaMmJHCstcb1UDHm0yyXkhdMdrdS7qM8+U+s1lBH
h/H7LP5QxMwOtPlxOg0QAqLNh8j9htc1cqV0bSk0vd/4otF+/SFuj1+SPMQ/Kb4w
8voF5+UBWlqjC13fkUqPQh+IprlV4wtJbZoSV4o1XBEAoXEYYYthtd9rDwxaiyXR
YHCYLBS7sRp03Vjl1U3IoiWIqD02aL68iUBOHom8+UT7Es3ZbGlJNg3hkE5ezgmK
f8cHLQbx0QwODqRAhivKMFWFB1Mg4Fwxkmt2gnXGJnRhyi2fLLDbxm+zeaD9BWrC
xzVm8/45HQywV4/OQrmjKjG6EGbPGzro/SD4VgVV0+gh17JS4PqkUrbVl1yXCSqs
KSsByGuw/jmUpx/kQG3K0JtvIxW39nqBrtQVRJUjl5GWZJuKiP5QnBKtqs5mQ5YW
b9O9zjzXBlI0fg7rKZllHhM6kxM82ZiX3tRTSCdH1ngZC3tQ5P3l1JvWOa4eBr6E
FmDDzP4sg8wDFGEOixIwKASZTswLG/jcA3TD9k8DGrM7mkrdRpMNAXaIglIUB7IZ
LIJEos6tTB2AcvjR5boqUVNsC/VrvHVZdsdjHzPMn2e1I7cEQfDdZWpWJVcU+1SR
tJ95uv51p5Fv5TcpDu7Ooz//bQpHupVd//AavzVZWDTl7c6yi/M7F3JlDxM9pTil
nO08cLW//3uxz8/spYsWewQx1+hm/e8NbDyVo4voCkLt/594rl5KzwfMJ+GwH8cc
WgynYy/PzFhem3hp44PqVA1VXvu9RpXSrKoUhuylNGAgJDW+8TLL0mPT+qBnxFmr
0+mv84te7Cj1Vnymz51b3RprG6B+G4Wa4SEtFIqu6VtzGxd9Cb2rdH2i3opREn58
7VO+8wUW0uOAw/W4asRkC6Mejjx8UW4LYqbbiuCVNjtW4ZNaJxNc+PDIAuQU5yvy
NdJrIlJP/i2o13YktNNyzD5IoDGZzdpt3S/zXlHrjrYWTWTnkrKNhxql30LnScju
+aioWPY1mHYUG0z/rMoX3+XeXGQG4LUFLw/VsfFCNK1woMqiGpix96nfdxKSFGKj
dUVTV6piCTXKjq5F4QOOT9cArvguBGQQkuDLRD5O+0sJYz90Hlwj6KFMCjRhuv7F
GXpo45Zp9susLkaWr9q5y4zBt19shpYGTy325RA7exG0gSAzDdcjp95+W/mARoh6
xckCTLS0j/dS9g8YZ2B7ouK+VWr5lTpEB37egxWDwvzJ99D/AwVrr+FfUNpvw+2t
A4A2rOw8wLiL9gVcUunsT+/fDB/naCbQJq/4w/LCsIrtXGwaRkPZGUB/18VdetLt
ZamtghjRtOnTd7PqQE8aNL9bGEFsJDmjQHTZ+jCPODTSr1pyt0Qlx+AIiQ4kggEs
8LKYGLuKI5CxzolVOBJbdVbQ4tXu5uacn2g4OB7txPEEdkMGMN09vvttQY897Uw5
N6TQTmn8me55gdaEUorE90QcQj2qfY/cu/saQYFf3wbG5+GRbSF06RDVSS/uQINw
qwnNaitJPhSBYFoVQLYu4arIzdE64TdMpIf8FXK4Q7GPrdOA1fjHRCvzVrPkrBhq
Yk4hHy40t4WRlmTd/oL3IT+mrdJ25pPyedrQsGdFojycWzFPAILTrBnndoxRSd5N
W9q5HHUvoJ1r+s6OxR2Qgsg783RPF6KbhChlXkWV+Y5bUh8Up5DdAx6EihWknhdz
N1bCKtxH4SmINY9Ye7XE1NWyIdpcNFksysKhGgq5/4+xljpbcRyWMC7Ke+1AtPkW
Ui0H0vFUNeq7TsnUQf8zJ5aj/4IvcVQaujl1vvtAQVseOlq3LWv2x1/q9AlUYTLI
RZMzqO+FhQV+3Ub06cvXlWMFOnq/ETn704lzTlqcUAP9RVGXDJkbe6QtVg4wOs1k
FqbLg4r2lJ6g+TigTUETE97wYgba3dd8AGenF0r4rFExWAXQdXYThEhXXcxSj/42
D7EmPyV6DwpNJyOFVH919iWFbi/1D8VRpE8lBZnfofZ5PFWbkKlRw+ALF40S9E1+
BxGCQFVqL83MPNXML+oMFi6MNkHDyFiYGFaNkcyMkOvlrhLDiZUi8WM5ADWwsq98
aMXI/cxwBPiSfHRVJQSpENA9NqvOAaSqSqMU87Qi6a0xrl41UkCvi2WG4/mG59Gz
1hxRmfEcdV526T0/jr2N8BFY5OSl3vXKJIdbJgjsUKr2y4dqiUi4IHGmn1VfazKg
895bB9AAZ6DqLhdHKSN7aVjzNrVdtYyCcHHjUnPMr31Zuiyo3QEoLcnMV26VSc3o
blA3zOHLRelsmcS5P2fIoPtjCXn5VTg1m+hpzK3sS2OLYYeYIlIYnR6vc45k7Kfq
tKvem4qnZkmn+LEpkwK0GFWsDCQCVhoNtXKJx+JEwPLK+1TXAPmvnvOwc8E9K/jI
8FKlmewNCSafanWS/Nsstd1uyB3B9Ui24jX+mCbL4TaE5CcibQAR0Ac47wjw5ViV
vFpfZ4F8mlAVgoWDFFatmvcWt7zM4R8DkHpZyagkQsR+EzP5wJwKdy+HYskBP58A
tAgcWhmh+qm1olUSUh/sonKycFEDinKQImFPW5IIxPyUttMVTCAf3R9PzwyOUs/Y
NYZwvT9Uu2W0+l6aclW+/an2eMSPKARCRcvAuGrqd3mxzDUHKbo81/tyIu0oCLgZ
eOSiXKPeRQrdlJVQxFfHpsTPWz2pP/u7p1r7h0LGY4sHhMTFj+aYxV43IU61H4NL
4he+8f4usUHqAj/l14RzT2oCAv5tLLkHnjRJy5g20//ckgW8b3ZMf1lpjjSMUc0s
X/wURg6gGsea2zljU+9QL/V/Lz2UQNjgoFw1lvs/PsIjTpLjGqAdeswiUa6iqWKv
iRdmhyfxw9grDgXrmBfanz0xSICTqXEQprPYMZpWqTet7XuAb9vTMbOwq0H8FoWe
RjeyVXQ7OMeWqHwep3HhZP7UJOU2ZjjzeW/O3BigVH5+3B8da0lgDDi8ZWMTZK6J
lPvs806+qc+VMgSf9algyna57YR+FcOlB9mTYJJooXJM56/eYIlP/Czy8nl71N47
s/vI0HPsgVMvRYCoyZJt3nbrqYuLh8fQaTU+4QHo0wrgveXEgn3dO1FReEwP3A/U
OlXbTy1lQZyjzG3ZHDa5OVhdk52XwIiB+kn1DtLqlJZEAlfZ1+PTGzT8hQX10yu2
JEY03z1+KDRi40s/GSPPldh6SrwuU1UYnbSNdBjBOOjnMwAOdVRZShsZSiAdZ9wq
dMZSG1VcgJ1DnA8xZXBC7vvK+IfiEseXCZwZPzFoO27A0tn1RQ5yWUtgF0OnnmKU
zwy2hVyhhgjKhqqJN8Yq32DpChoJY/IAFZE3/e5x9+9ofAtAOtsWQx2+c86WDJgw
94JaohXO6ilPVkk2vXACFWmecznzr3PfVhLkad8ESNQ0StR41IFcCiumzh4zXIbT
/oJs1dgohLfHTG1uXwwB9E1m6SCWM2jXGH9Ct96UF8np+vgauiRS4qO25CnE6DOr
wl9I3u30V61J7bOXMNgrV5nhnGe1rvu9GwsyVFXIxrDcU0wu2aiZWDXeQRwAvGYn
wQ+L6UrpJ/MSfn56M2N0T1UmFD6+egm465cfUF6ZPKMgoAJ4d0LFetnlykjN8gHl
8gO2jsIS2nDjCJdabYgjm9FmAr9RnzB+EJEwGLZlEiB62cDIEsgGeFJghMf3V0vb
iFCZCOd++u1iCXqfJQOC2kB3U5rrojrXDFpZoDI9XZtMpP7U7on4R+83c+tm0XhD
FzGrn+xfICvp6sPDlume/4r4e/L3JjOOmy/w8WtoIZu/pwl549Yx49Ya36JeSF3R
8/W/J6DxUx5FbICdHKkK2eFbduiLxgBTDNfJ15iP7ML6q3m854Z5RE92+2vM0mIO
uY6syJSMuV7klV1rds8YoJYhRwtwjdyqL4dqrGD6Hltysz57XPsho5oAlA5AykUD
TM58OKg4F4Sublqb4nTNDioG1Ljl1EBSVNAJAeuXC12Q+6jHbHl5LWIPfjENv6OU
8nsMBoI5B7to6pSMd9j7pRFjxIqYYPSXkk9Rf+6TDUBU+o2Novkrbg92aQoKov2r
G23tJQBOMuWUN0VJ52xUtXhhMYZTFIoyHLDw7NqJkuHbuDGYLllTa3M+rfIrTKi8
6+hMIIMqp76xB4KWu56665mQZotoD2OanjgA4Hb55cOaSpCGDvnPtNffnCxpiURI
/QaWUzO2FvVAD30NCUr4crjVPJVn6wpA0cEEqszWQQRpNaSm9LWVanXmx0R8YqjT
Yr/LhS/EMPIuzi7pFsy7Sh/z1WUUF4k8/wT1S8yC1cF9sX5JJT8l9/qfZxDcaSR/
3rQIXMqa1YWrJThSqf05BfFh/o4LxQGlYXH2fdkaT3gTOtxReYm7aXBLaXtuXZ03
SAGEF8PQl43sGPNMHho2eUaeqb6rLBstfq78MCOAfqDthaRY910mhf4G5v17FZqD
S3YOlBhA0kQrzGwun3LqevbuW8druar6hEbCdHvrxwF++Vf0Qkwb34cFp8wyRq+p
iozEnaVNWp9zYoSKa5ZqqbA57BLglxuUn4PfL93GVhKThlzvbJkEI9iuBzEhSBBh
47I7l+lYkUHuaEZYhfBlqqKW46Q1iAFGNvxv+cgv+94mCY5f1/yV22pEhan6g9a9
rK3LQubNanV1np5DUOnH18HehSfTffOo9kIeBUy+LA5159HYD66n/BcPdJgEbA99
3hoHbpgHjSxa/h0CM7fpEfNJNXO6tHqCY0FN+8VyJQ1vH+tproIxuHxCXlhYQYSJ
yY05pbgTIAXKdBPmpyB534yME/uDDrviAP5PItHAlI6TJj0nxQZurppnbGvibdnq
V/9lCqpcjx6sZlx2kvKUzviEQz0BBAQRg/PKkuK4KkcadOrDbXiQfVM5kqpS/7Ds
VL3uQdVBWAXRx6VtXiyfpU+cd3fUrZxNLr0R3/YwMKLJGbfXu/osZ3xHrUNCNARX
jzXBh+HahcLohB+ksB+YBnOJ/7cUUwlnXUdZHj+NHobQP+kqTiE+Y5brutPy9CVA
Y+9/FRk0/z9R/lwk7OpDUD8OPWrvkwHiDVHN5I1lr22qGylhpi0DxXOp1GKMjvG4
JI/DC0n1qh0PJ2bJjbfgQNzIDqYD+Qh582u0mbQl2qErlfMQaUudt5DjXyoQSTy4
H3ceNU2k/V5eo4IUGwkrO5Q/+k/Y0hqQnDJPt4k7v97NrOgzHY3tU+HNTYknIodt
9+cvHtzq1MxL2XnWeMIpFu44eJsXqx0rxhPZq9lZdEqUldDd8lZKrtSAC7lNmuP7
+v0QK2WgPxowLatPF+B5Er30kBZF2rEJ5H19DjIFqvmOnXbkI8Dc3m+Es5IYWQL0
is7bk3rjNGKVycfZttiiPPC8ioyRAvvOHW8K/ohDxyRTcDCsMvGt3UGTPRzJPlG9
aV0deDNJu3MXhrGl20QkRDoIxlXCUm/ZceWrCEIeLoPGsLdhRuOV3AVCINEsIddX
uohH7xDm2tDXzzuNBzd3Lr2WKpzXPSP6mHEk2b+TE9pEPIiFcNdmx5wgIeQGwNK4
m89LQPic/1R6vh3ReIVAiwr6i0elLn5HTCkFSMwThRTG4sCEunbxUYVRHb/hrHPO
vS0Wge8R/TydMTmL3jA2nJ3BHng0sy8aSR9WD+nxYJhUf12JWrO6AJjKPKmYqnli
vGnWzJeCZ/jz+1fo1z34Un/ODSvrr5UiqQDjjXsUjiQSAXKmn3PZoyMEVNzCzdW/
OCpMbx+ljDe/s6tgUTyjWPRqZj2og9bckNMvDl/jZjVsMeGlRAyNLf53G61YZuiA
/Pf1rI87kyBFzzNnYeNwDQHD/xbnfpURsfUP/T0+89ucfzJfZ6KzQbMdb7YlhXqd
2dG51IR30OF2pBQbtzk7hO8mIlBjMG9PwYtvVZVbCziLkJ/JV3RoxuvPDYGzwUdB
Cdqf+Iy5c51oqN9rt39bARW3+h+ejV0yqu4173bV/KbohWeuU22qyJfHGNmzgrB/
Perh+HOA07JTdhc/AbNuNLU3PYLp98NakiHEq9opDmC6JJXP/7EqZzAPurQzw5Xa
ukCfFt0XzJVXE79YdTp6pRlW0Ukikb6kVWGkDr6Xa4um13FE9diOQ3gLW1XbknxM
qeF1cDDTmNHIakWdrl6n1k0gpnrUeoptunOjETyc+z+xfIqOcQZbbXCjXycSN7kR
T+UsY98KtgGPBL4ySsuld6wUnGvEViqs3BwrK7pXrmqEbnBBFwjXNgkT3s08N8hW
TcSyJ9b3NnOuBOD15pWRznpwziNlDVdwT1HrkCYNdfz0+17RExgATS9TtqvpF1m2
CTJ58H38Czs4TezLr0KJPdes5ZqDNzbK8NP8vwN8jzK27ryiOpKPUn55fVo93+py
phGcR8GPpmyDNCZYYvAmxJdYT6Pb1KC8++F2lpINsi4Teo1aXBUkLDh2tRnybCyY
Ma8E1zBRI1OxbwybKOklO3R64UwaIBIaHEs7mp9Zu7e05rPsloXZXx8/EpYm0JBi
b4o1p9/csXRAtCj5DMchb/5qQMWhftETSdY+kVTUBntNSD2Fysrva5Q6Qf6P9qTl
6nkg2tfDhQ3aLOOnTTIKwqsQT6PV7iEN0WmtNeLpanq1TdowLS/+E8TvVWVKKpec
n0VFCkgeWjp4FDxpGEtJsTycHvfsr5nvnrU49Urh/HMMeZhmJdYiw/vGqvWCpY6N
4ehUpX/Lr+EurRJA4Xi2SJEAMffV7CRLyNDknM2C8KC+lT5wZRpu5Ad+zSUgpaW4
/4MA3d5badYE4rKmPBxIyOSVgGsIlvC7sHrsg0nQUGch95R8HHp2pnWfe+LIOAuJ
kFNCex+lzBCZyemtWU8uJqKmcm5M/YgFZFfFQo93smayIpzVMWE/qAdKapIvFHN9
Z8HeCbV9TwTsFIbVYSevVO7wSwXpQEAvYiJp1ojs1NZlo3R0YTe3hPDSRffwFuj6
qMZbdSOF2gp9AC6+79S17arBG9khYQZagvM6Z36j0b7r2NA6AaDcP+98Pl33tPMx
g8HeH80bLE04SPk+AdXqS5O8gxhm9IpSGJy73H/6ip5UCFFj5usJ0jEAxT8uDvLN
4eP2Djq6meyH2ZwW57haIEixG4MQrPxUpgTmKiTJhz0volzm+4l8XcZ6NkUSNx1z
McUB6EUuwPsWufOJySTyjf9dgKlIFQUMzUvEV9UpxB8AYwb4pFmf/+SVuHM0PoB8
2XF/smJe+9Is46Hc0PyJnN4WqLwxRlvsZAK+tB/FtO+xr00c/x/DTnI2nGDBAuOB
PBpFmp3nmrtXzhv+MQuebcszSIP/oZgKEB/K9VODtmx6sXAEZouJ2MSlypC9DcpJ
+892i2AKWh510du1arwDM2EhNMXohZ6C1EwAIXzVAM5lrPPgGi/h6Qq4RZB+Y9ek
ZQu80y58a4izTnLmKz7l14m6pl0vC65+0lspEikGnmmryXuwKfzhs+dsX2HUi40p
G59iIOdSCGMEJBWyftc1iMIkgikyuK3+vt95wQEaZFSZBFF06dQAz5SBriRJrJbY
vO0my/VrRlosHFPcBwX6yV7p/IAsZBP9yLkvSyvZAGTY0JHjp6txdpWDenIpagmD
H4eMXd4tkmhNjd0s+D5Yug0ywkBRdMKxL+LuSP27DMUkmpUzEzBH10gNm47Q/obU
v6WlQqapq2fGy4MciWuCYNJsnO6tmPwNotMhWFFM/8yWbhz5XhZKhHKQfxX2ynBJ
sKky6fzWLjJW2WuXkigQpA7To8+xqdpvSs8MAcRRVlwVr5bAy/qqo+oCTr5ceYNa
IeZ0Sv5s830Arbo2wgBWfQM5rQa1MsOv6URk87pnhfTqSIN1WxEBAQXIG7ZtNKHn
TCz2zDQxoRT57gtFSHwwBdzioWvDuCeNMGDZpGnxZqx5e8iNd/GjLlv8n2aPsnMO
ZTZajC1VBEu+xeL++TIsbThGFPgioUzP1pXwiWnfBNLQaotc0bcQwfLKODDXYzPc
xNnrflxeyeRsaZo08Xp6+FjnfCxiC31U2aSnX3BAcZZncqLVm12iaJD+Wn3VHoQf
77+YuDJyln5ZZyBSX4ZxiwLVs9wxZrsI2GeaWfGn1NmaouzXwqqzgc8/xEL1+Yj5
1uwYdVIjBZGBZNf7jPEqPSgFNGsWcdKVxinySslwpPskch10YMKGOquqBR7kXcsv
jTrM9HBY+vHfr4Fs1/dJMTDWR9917d9PcuPx3DSiBXWNCTDbsanlywYkKeYhx9W6
B5jEiXY0Hx6H9vFBzRnsQISqE1wWKmqBIK/VoH+P9zBta/iBExrM5NnCrXVeEMKu
fw1FzzPyDTkQ0GWIT2T7/nanbktC4NArJcdWqenarpYXA5hrdUvFMJT6aHRxSHD7
ECqi8FH6I5IZnzDN9jhVwho4T6EUFEWeuYmvEURtv6BkVrmFqceI4FwnzCsaudgj
JQDgSsU47yjsCcxRqbea2AOg81QbQngrK9DhoFXAs8kaQCqXXyLg0G5/2+Pf1u0c
Hiu3xLtnNdRoQe0UGkSmCFmkaNBOh+JoqrmY68oK96aW8e1jAQAUUPPHbCBnfY3Y
YEyWJVODLmAnDXECufovmS9FLsFSWy0O/6Y5uMQHZzrI2yisBtMyoORZZYZ9KXyc
P7x5a4CoV3F+TyVn2NdLowDG7TntYAwwCDoIiYFTXigIgAGu98AE6AMRyW5EHKLf
W/PMZhKpYstzVnHNtdazCuDFWbEONWQ/6BT2lHH/Q5J1Fu8/np/kPu09+P//ALYx
GbrqoKdcC8EapO69xQ9TVFunDVLkZtcFSN40wVcBzFEBg9zSF8gGBrJVrzckO+dw
mboJcCR4D9kEpVNFq8iNuCK96U6dFR6Qm3fom+cbTTB6WMilSbgwy97RohlS7wRd
RyBSpSMrxr7/DhyJYTbZAmbD7NyU1Thffkw2x6ALJDVQRRIL9HG/OBoUpAEKigQt
JyuDFGzxoRkIDOF1nebpRcwWcspSr6TMFK8DlHGyianxeSc21auFPsdrSRzKGCSl
NAvyxCTiNbk/Y5kckKbiJP04Wb6I+i4Rw08QQnzKAitSq6q6yYJydC+GlSmprXku
7bg8EiXQ45j8ry8vcodno8Do80Tj9bbvmPmAnhGnqVIn81za4eubdw5BF2Ud6iX5
HPrnMEm3NefgitU9nd36WQab9GFYx8T6RZ4RURkV2X83i9RXbPKLhDW9bjx7JTgI
IJOSLxWkfJI0iPu85jIqTjoMmrYek/sL+a/Ync1UXtgzowNF46Dl/4LVjJ1h32VR
KQUT3ukZ3dzy1U0/qFQxUp6BSejQofT5BW7e9yK/7tZpJpDCr51hZ7iSVM4Gw5vv
4pZl0dEVClx6PLRpAvuW0o9idMcbUr1qz1Qp57TASB6qm4CrAkdkGTECzZz5/Smo
3ZZdrReGA18kXHmGRpIUdIcTO84JM8kBvJP/hsT+DdSLHs3Y11XX9lGPS3AO51cB
wMTRc+4jAN+e6tKk/OlPhANE8/QnctKe6tZX4D0LCXrvbTCEQYsm3+0L2IcG3H1/
Ha8ur6ftU4SBQdK0PtB3JYK8Tw5ZVzAN9sCvTj/jCuIUTkQ+ZB/aYR/isaBe+EMk
7o2p7uR7BZ6sxY6hbpQLRD3tz5TfWqF8KLSYJIhW8cK1okYT16kYmih3wX0S2cMy
9yU62HLllFHDM5kktyxfaLJy9YsjRR8995WJ/XTIcPm2mP/KGoPDsegC95QuFQM/
ImK3QAGn5lgAm42mTiOW2mMAKgZjddo9QHiMhrCQA5rLADw9drR8qacNu/W3Djbr
Zgj6mpbK1exYgEkwDjdZi+4XeqEQX3k936pjXNIBlvDfKHSOYZabkFgjdXmK/vA0
CKWwUeAxIrx3XoCOhb4dTYN9UsT8cdU1BLqM4T16GUKQy2MtlTCWdh/bKZiKxQZP
4soPpd/IqZBBUTsz2uhD2kTLjh+iMgd2tvJWoyjmkWxT/NgyMPEw2E89KMkUhC/m
2rvIMnuVht4ZQv2mOiaqccqU1SkzZPnxkh0+FG8FDeH/zgRMOlMcU0yVKLT5ZPB1
OjvO+9DQqJLi//hOArWuqpSpFWNLEyvZgL0/Bl0xFMXRYs2wd819eWr9oAJkNKhe
jbtyIxsftED7vkmBcLD6gXlCW5w1OBW/0oz0cP42XjpUrh7xPL6AezRynt8HbUIW
gkm3yzI6hAv06tibrPAM7dukCTtNLgdLy/Xh9Qf96xk1fZiLqFlQVtzf/u7Znx8v
4EIOceFqNfHnKgAtQMNLJl1TifEP1ynsy9fUrYfiYuG8qxdepC/tpW8CI8q0nIzH
/f71PJKI6bX6214095oySmtZJSaR+iSuqbBEf2iWKg4/yZF1n1AMyMSZIOrkwCR7
pWslh2GosBDae9p3r8KPcD085NsvcRvYHwmGVD/0y3U3HouZP+ekh6fmnYNz5VKj
/q0XMxELfENb6QSVt/VL6xGQbsPFlPWCcpE+ey47EyU++qk55LZkgc7FJ5wtjG21
jznF3BXdmO6+K4JBeo4kqMJsoRJCuCcEBgK/uC5P370snZaiHe3hW9K4Q24QFGh9
v0shRe7+nztt5vV0Yji6L4LN81sM+wDUor3+NCVRwoMEalpVvX6ZfizE0eDUT25+
+ZJvNgPSmN4SygPeaqy87tDsBYvmVrrMgnXnSco/f9hvFDmewx3iCL7eGKDRhMaq
YBUdIeigdDW2QSoPASPQH65yAevZJvbFcP5EG3tz42H2kEuQEkCkrZFLvFALA+i7
QkQrxrgFJD8Hu7xaRvjinOWeKJw9LddKlS1nBqD5MosXHt9J7RQe9D2lTawCzABA
3P4NzOfawTmxkz3oRJmmNliU2xqubU70al3m7EHbgd8sxYsunumzjKL101Jxztl0
/sRlTuCx87mmLl1Uo6f0jwCA1e4CeQdX1NyV+c5e6VmcNNvZyh8HnVjanDasdtjc
egkVsGArzu8aCB88c2+lfvAtmzSFSuBxKgVke2DYQNrTn8SH4Q37E1afamJE1yl6
MR2Tvu3S0x1djrQLIgoAB/oI0FdsOPjaa8UEARAQJ45s6Dotc/JO4ikQYuk8wZjx
rnsYjH4a0+XfWYnlGJoI9LnCbCvVDq98rv4Yz6lyDL7WlvpnqRbdzrMJ+Wt+gaW1
46nRv2lYu0TTGgyPBOE6esSWYAqRrbZNfwq6WwEst0gUFmr00eGMlKvbTkYRneCj
OavlM7OTMX4zE7TdQkkohAUS0izi9QP+jz0yTxWT81hNQPrwQnkzA8WZB93omRtX
RdgxsWtQOcfiXi5c5/+thPCypzTycJmR5F/xk1tWURVtVaw4dPq1GITQVo2c1Lqu
EdDZzA9Z/ApzT4Pki65OucKd9POKZjq5BolSMMsAhIiV+La6NYoTViMh70eLWCE/
xSvZhXrd5pbjVCHCfBJOTqoDDbEIkhjM9aNTulfUdionQHAMvFv4ziPWGE+AwAI0
G+iVdHw4Jq4CZVq6r213kIWJ5XE3X8tq0RlEp5dRxMd2iIfWCIzSz/khGHNRW63q
hBlTw9fu1usJtOVgHk6NXT62uNPdk2Xx7lQBTnEpig6HX+ALBkHs13eEGbJfWFKs
X99BbXBUjR2AW+Nz1JBy2h56allmxM21qtwWMuT79QZliH/u2rn2KM3CWaoFk//l
l3IBDgZU2/C3RmhjROjBFO0SmVTIh51RE+s3k5AAtN5+5+LlozUtozFr43BpTyGu
PDXy/0VpFpelorwAWA+zhaNi4l4Vj5vMpRomWWXIl0vaxyDADAEosKmJ/YuZbw6c
eNUQo9CX3hxr3qkb+2Xn/sgLQFbdwjtivryQu7A6z2gP7Ooxr/MdJJKTdDxuyCKe
ishACiSw5wd84hlmkaEzi6tlFxpvjrgol60CYw9Z/i76KF5e4VirrI8Fq8B+Fo5b
y5QIykBWIsPQFS8bSMSf2sauDzI6NU7Yac+v815sbr+KeyuIE27b/2xPj7VbQmz2
f9TG8rV2fG3H38boRvsDkuyHxw2FGAReM8dM/C10j2uYEPnRYqsPvNqrj8yLEq8I
M3L3dyuffPSNBn4rIZGtykpHGZWxI+vKzffWdsPGv6F9IKbEOfemhZ50AVWC6fYe
+ut7mk1yRikg/31IZN0OwkdPpMUPCV5asW27kAS/EXYojFKJRJczD8wWZkPz/MKA
oz4/nqPPVZRn8lLYwWsA6UESSsOZ3v5s9ESdFDTXJ3LxbjrjZka5Ebs2w3KYm3lO
+ZZHHqgXtCXgaAUuDBCZ7OadThbiLqX8915NZj/RsQjsVoTZKXfMM6MVBTIR9jUJ
sfaspoenx6jLZPSycuRVLsBCfCJJHfB+N7Rf+9xMPyW9YBDcv/ySPfVrueNVNwTC
R/t2XqioxG5kBkn5qEGojfT06PwfiWEcb+oRlON1NOG/WziI9SdomjN981US8Nti
lGYrCtQxxQqCemb+hdwfJnvlBvXtPTsjbl3kN2ZLF16RvIGe5iebMfD2hA4jUv5y
h0niFI/ZRzucmQ6s4Ck+e//LhXvUtZ8+3zBEAC3zlAkxdNs5/9K+dErGsju7AeKV
f7LNkwMaySEewE/N+AVWzPPnXENjYApxpQzztDlDf7YbAvbPEO77OU859Goqjn5c
6nWwkKeAemeIM5iXivH5vjrLBN3kuoD5BS2raAA6IgLc04vuAQ2LlInUzc8vnoco
ViqSU4cwMLZOqWlCKiS0f/AYy9K3ZkFE4k4T2e8RRHyhsF4/BVJ3tjPNssELrtSx
SyBzbY7qCei0hh/OVehOw7rSpmsPCd+n/BCDmx+I7ITj2ROVIxo8tCXgW9DB+HHp
ltbHk0gjvwrzWlOX85fmYZ7HVx09icVsvSU4cOACSQ/JAWnsU84QLQ/eYnJlsgHX
vqQ6ynpoTSpUV9IcZShHu5dDYszJXmXKb9Y4UsIzOaJdTCZ9XUPYGeBOmyLzW3pi
qSIP/sMQz9VnFwFmW3fHveMhwztg6MdTLTq59I8FcTcDmFn4jl7AXRSkfJdAoRXi
LBjtNRlZtJf2DUBm1sREnMbvuiBfDHj0wUBGDgiwZsb6zUjkB+YXQlqUyENnrRIK
Ocd6oW3Ef7CzS+nqXFQeqyyBgh6bWa18hq8GwLrv0kzqLhf3Fb+YRYVI3TmQo62A
88Ue3lNRH6Wygk0Gm6Jc/gsxvXGgRaugBNAAUeMUmh0I7ONHjUbVeeRfp4ud2nI7
lBydggGkDIKpzNMnvjibTccvpBkPKKlo0BSsBvuRWDhLbJhxY4FG/UnHldDxh1hg
BkSnkCOcSlAulEah/4h0B2XaEN8mqMUTXBnulmIqL9NfIiLgh9C4HO+xd9OcM0jS
aExYHAEfCNw9itsj9qGHrSS6YUS/ptkcDBuksn4+hvflTnBIRddT40LnlgKA4F3Y
xwS+gCnKsdF5nCL7u+infpP9igTdtQzruikoiZXLGI/l6TFSlegGaVbkiwOgb8dD
mzSRsKcHN24cZzM9LrXCujFaAdAhFXBPKWu3XXkraD3J4sBJ2sq/183/hDdBZfh+
gsxWJQNBuwlNpzvSJ+g2B6V1PiPNVCwK//Q23ZFpF0v6MS10RUJvC4DvG0ly0O4i
ZlpAdzeHNW0JgFnhRtunDvD+UHmPxnslEk+Tkip83zxq9zTVWgCYiYm0Tl6ogvV8
QC5gEVMa+UlmMY8OoLmmm8tZ4MVMGQJhkHrunST1+eGJHnHz082zsyNjjPIJk1ya
dlQq2uK5IJ8MFrJ1lZx7KskXs407+ZYymmbV4nILDsErWAg2frO0KSPacwTDy39Z
bQg5fYTzrHQ5SkCTMSHTW9uXIjXrqSve4iVwKbcEYzVGI9KVYCclt294/xZdhL43
9kTnzsnAs31mKT+LkFt7EdjpAoqLX0swx2kL/OcfuQUqYp7iNd5KchbFQl+upRmP
iGHiMTBrt9ZV8xp8FjQqdoIOECTA8ieHw+Zme8SmE89z0a3mD5X/AS7ibTkjCnud
Im62m7OBi3alZhG5xp/UQi3M8W6Ua7nwHZFbmvFS+/OUzv7V4WAWLV+nGkn3XtVx
T5oY09diEm2ImAG9JthNRFFbHVckiYbX/iuRDmIKj+lBE/eGXjUyk3sxnIheAePr
+Zg1KtyQNgKbWYsEyPYqj3M445+TRmqD3WLXkPICHJiZ2NzRhz8hUK68Uh/jG/Qt
YhU+6yJrmoyb0KMbHio07lnyUlmDMawCVbpfBRlH1jZwHoSdO/AaeF2E1tcp2zao
6rCzVRLZfO1IlHjDXbbXAJ1adAZwNF0clVfPdIUHYJhep0ayT9wca0so/3GA/UHk
o5jOyjDTJdEgFuHUsoXK8+ZqI/yIZhrDwIhwwR8MV2BNek7x5BN/xB72FPSB53YH
XNjUGcka+snSw/QRlho5ZwRz7Z2YahG+PkO1tMBeBHkyulbG9oYws/IP4A22fY7E
IlnMJ1dk0ROHP23bniZYND6eQ24OXqLuukwJ3SsoFZM7EznLmU/fYcYkss6rzesJ
NTJ1Pux5wxxHCzvZn6BAajSyJq//EWzo45oQWrmi05WLPh6cV9zMd9ieclmOH3ap
MH/ymk3Ok67VhBvDPeClH9V+vP2RI6GmfJAq10FSR6HlxLfgDRq+i4FGVztKXstv
g88A/JTv2z0Tci2ZLEJ4zPn6aLm2w0GzFVTvPqma0X4Ja+53oSNdCsxUNI94DvP1
PN731svZaxoDHyl88s3fYZOGAiMkG5ity8l7t12HsGC0l9A83zHh3hxJZGHJJxB2
KecR4S1TjJ/dJX0PbESLXHptCiyWO3LcmXlxrPWXXDq8swL/vtXb2dFf+ddmMBRP
aFsOF+Nv2CkhIknAxqtexX81YD0al9Vl9UdXPy8Kc5iF3XWH0bGDhg1rnqfiNZoP
YVtsoXRsRM+euoy0vSKukXOUtNKme4TDq6iOZe9W+Q2knZj0xvYZCZxbDkEjDZHO
6zw/m5esTjgqbFbAVVdhrl9DiLcKJkYo4v25pkqkrKIVDGwfQuupT+vJhRypthOE
EFaKh77slgl3OoH89v15vlJsVjVJo1DJEqpH4khD1Qu0D/WcYAmqgx8gk5CUxxxI
FggxYRzDKFDKRQaTJCjgRRUZ+8wwtwQouVa8FjDqdyOLUvgkNL5HFdrwvPlNGfFk
X4GVggSrH5PvLZmdbK95Lt6hEyoRVB7o0fgEiJVOwdRAi5Tz+MPI/cpkKxi/o0dx
ytuk+8D/FCaDy0XPrsntD+L77z4LCOWCOQDyCqmJzDQEdpJE4/Taw99+W4vgN16h
eQ8uy+3CAxKMcTNisAsi8BnBec/t1snQ1fEnaZWw5zA0DRCFeAC2ZGTQkuMSHbog
0LoMGBqhWAMF6IL3gOzIiQGwHvQ8+NG6F8TZUDBtUGAc0Lf+ZgtMDPuajXX7GnJg
DmwcTzY2JznNlS6wDUuX6lfWZhhMDm6d6/+LP3zhO6CBuexgEflt+JSTIKaF/2Y9
S60Q109HqwhhrYdEUVGvfsF8stPhOMfsoVjoA2zJCHuv/DbKaCeKeJrO72VrV3V5
t2zTYvzeMtR+dxvzdv8q0PjWyTgP9zRuaU9n/JaA8US47ViJhzlqudTvSu78Ak0a
24O1aMPmrzd1kl6FWDUnB4jxHebRKuMXdr/S5RRi5A93n/RG0/oeZ8p7jLqK786o
0syAmNcDoW9UT0EDZnzV71EPTDhU68pRTEJUWaHpXso01NAw4LJV2FtrEyTdX+yW
px0JSD8NrEYAVsrRGZslFE5JeSL5Y0/EXUxUU3LOccou3rAcyurVcdJTnGQNzqLL
KXYotu15TgMyOtgahaC8Sr27I/CnZDJXP00rK3diQgOn5HfONNahmtQ87g4FgKf4
vAuRlYVn2HuKYa2hU+hlXNZ19/QzJOeS+RB/KeyEnMsXttOhsx5ntQv6NQnN2OsW
JXTfql+TK9QuyTVRwzyzKhnkiKt980ACjeriJWpu8Ds7Gtcot0Dok1kRAD1+Zw10
RgvUVauzuN1NuQKYWZzJFzYCmOoz6iBFGklZ02Ebp2dnCTHk6sVVaWoEo5BON67Y
uaESIozPKo5xru3nb3IPtqwlXfnVmoVe6t4kftfV/RB+vpFKO252N6GwqqL6HbAa
90S+q/7Dk2278sRN4vj57p61yFe5UHmaFq57dtJrkwTpkh4ZIQdHZg6KmUBTpoUi
C28LYuMuejV+isTLPZZlPtH/EMWyJovp1/CWLrhLj8PNHT5Vb1UN7bmGcMr6O1G3
74t3dcUPNdOWZeUyPPQy+LZhyqg0cC9yOcS1fW+FmecJThzmsKZeF1fidMvsWGgu
r4tE4i8KmsK5+Nmim8iiqm4TLKGUt60RFyFmSwHFqSfhFYPupwGvblvl2DFgqbdr
J9CyF14LHDzOO1cCmmDnQsJGvZTm6jMVczTZ8DkGndAzATZ9iG4wTiHv0nq/e+lL
BHaNjfnW8X9M4YyOpESkDEQZ0lUXDNfkG/j48/ydwqhTCXAlYguY4CpotHg1iDQh
Kg35e+kPOzSn3i9xFptDgdKaBSzYDmtVSYZdvIaLVwn6Up2jw5UBvzvgPvmmnsvn
sYVOmuyyUW6N0wdkj+3CwsLVJnRQ7l+6uz0Wy1tgGxhdreiB0FN4csfncJtt3Kne
Jps5fpm/Er/v2HWS4p08C/gqcT8sUxTOlhgELL/ZjB8BY0bGBybD1pgbSO6mfXlr
y0RwbZJe4XWrynRy0qyumENhv9Del/oa476J2rzFEorJ8vtF5dRZ0EVjBxkJBtP1
s/XpwbLmXJk/FmwMGCHtnuP6/icJ6tNNHoiqpAs1cU/Mn39ndu5+p4ejNiZf6Cyc
8hwjophrS0ferdAAJp+2Qca7zcp/hn2wgTCoJr/g7pqMNcS0dG65OaEgfvo+Zt/l
p9EUP9eWDejquMWnV1A3asZRRxqoSwuN4eadWA3IRBaW0TlFILyeAgS3S05ptxoI
mDWpb8n8CDl998biOis4vjJkuNb7ZeRB/BGHlLNCdDADXXRbvBLTkruIN4EzlSlg
lfiOMQ04rMSkeOvoguJxrbCfRYEqi8hC6xz+3Nh4Xn1qNa3Xiwx7kulu9g+d8kH/
PvHV5EU5mZz6iO8JAHsFIKEwaGM24TXq4dZECba3f95NgGHlt10Zg3YDoNcG8vCb
O1ZOoic163V7uDp+KJWm1a8eLok8Fhfo2Dd1MXtA3lp757tVzrDN0cIqGVx2DyVF
hl7TrE8Kj+zzGHkKEnXFeojomfF3p5kukYqz6/t3H0UmHnAv4fZqZZEMzRSrTe37
e9YcQCaMw/CG8fx2+EMyLeDHFR7v4MQ3l+nucGeDw2rpzKeB+YILf+x8cOmy6ZkV
kQk7XgN+TTbhz7cONGVMnUk2n22W+K09qEjPhZQdh3bm46qxsaEhn3hIwmLYy0dU
hDdXYL15nk9IqBQ7LOEVMIsGGMgpSfTsmXwK1VzCDCMFzL8iYSQev/Egl+VNoquI
Y49tbPMCM4VNi0FqIyrTKi2w8g0ZUqsVhwsCwDjoK0htAHSKbaFDGr79BuTxKcSp
+7e9yS7Pg0Tffb28fkVajtsjJcrvUONFb07SdT3vra/MYCuvUkBsdmB9KJIAWUkA
OdlgpImtaA5zOk9XfVVTTnjBydBd+SzBhkKeFUNY5CLWRl4zi2+GOkrEkQjd9ywJ
GGmneVBlVYhgudn5xnAymO36Y54TbjpR3IsBR3EgBxu3sKmaL5/xo1DsGE5OX88B
a2ZbhXX9R6jbM84rOC7JIZ+uQaWIEcOafHfyuBY+SVXglw4emi/3kVHl+GwQk/a0
k3+5Uj3qS21yMJuEQ83OLpzVW9s5ie0i6Tu3Op3r49LImEX+DWRTWtKHgmfdh9ez
lDaFZgYx7i0NoEi6aggR/Zg+2n+QDd5zB5ofW9xhW+wxYBF1Qk2GTnq80Jl4bXlL
68+8cceqv/hSKbCMQ3pkbdaNrbS0oMFxNWnXRaFUsVsKWhsQAEQqUVFOYSePfyuh
twvnHCe9iRLpqL9qD2Yq66vg7kxqyErfzlvsIKuL0xIQlxHt1JKQJRhBItJVLI80
NysiRaEQ5spBu+nN8coQGl/a+j+19NJLwTNgGngZ/7ISLjUf4yM7wv+6o9Xf7beu
I81FC/Ohi4L7uC5Fw3miUq1DcB91U9cR6+ozbHjK8gVC61kehz0la4BpdFukJDjZ
H+hUBBgASUGSawZ/PIiSsNpgjfgnfj2G/sRmuwFkwHfLwKSI4klDY0nx5OkYqNps
G6phDj2/jM4jmy+48vlaTx4Js7vlUMyl1Pdw308TuW3H0DZD4n2kW7uryaYch3oQ
WF/7XJkCGsfDOPilvIdjnWjRmkAvlh+dugrSrCb236gBkLf6OB+PsyuwsvG+Q2MH
vDz2QzZ577DxnxcxQOu7oRYvDHiTS/w6pij6LAADbE3vkwtwtZ4adcMFSU+4wb6/
rzf5PnsDVgc+S1ADCakDoGoHlPj2CGTJEzULZW6gtun/V61U2COMGvIE0OwGrpqf
IY8+GtXbG2mlxdcBtsCLZsZiW0VRLq7kPVcBpaIyAAD8ObNn/4+5Tc4zU6DvAVx5
Hfnih669XWOxUb5tTnHlOHJv7RqMa2BTrQvzoiRehZ6eKU3jPZc5RY8uVSTucRWQ
PY2fGvRANKcO0J9ifE0celI77NBbTNUop4746RWS2TVetiJDUonxuLgTXA16r/sS
ZZ84QUN2vJKY2xkSsk0iFHyWB/qiQirTSnavXPNwNPrQbDikZ/inHSHYh0X54n7a
FYu3lyFARztpPqHjOttNK9zewBVneQEBvNMQwK3p2OSs5MamyKhrN1KZOeP+WHTw
v+EHpZOpfA3WJ/kuz9m/xo/NZAIp+tze69/iKBgfARXsMk3Hxn3+LsnEEBL84cYP
IsiEP9glY5JRA/Ixc+neMfVmwer7PKa2RoCKHJXAw2TzwIh07m2oDOQJFkNUO0vr
bHxWFQ4sLfPO8UEd90+m2rYNe8F6jn9pD17nQOv5l9oHIX+n+2PRUYc0RE/eEltn
FWkZxLfAYGe6duuzheKhSpVg1wEbUwu++8qYn87ekhgkWDcgkYDgxwLwRKN3T8ds
Fx8jdBuhYwO7nEQJrK6mItXrfSPmV0EB32b3sbNIkCTeFn6+AGt/yZQSqLaQiQzB
lDFUCkIi5JUi2BpuqUje08jQtdxIErrmkgGnTKDRJ+VMEyIy02MdzUi4AFztSqWT
vEaaNzprPliDv39xiPETF4jFw+/aUh5eYy5LnjZ4L6ZB2GvuXk3qBZlMONoIKAe/
3wiRzThMi4D6dudO1Hx0V/j6GDjP0D80jbr4RgKqLPiT5znNYmWe3Rm3TCRxm4M/
cgZbex9sWqSmGVHjk4gHrjk8SsBaxf6mX/VI0FoCStnqytPhvjJf0o5JYJVnRx3d
ymqbPt6ILlkGRJ2ot6Y0QkaPzF1MkXwj23QOzdCdWX+nIae8L9GNEcHFQB/0ycfF
z/NrZFQM9uwXpACq3BdH5/4woor5pkbkz/0VhUdEpt6eCkHXS5sCWC5jLOef2jz0
qvq6om6kUOFvTezXByUN+aUtNKnRJuaVm87N60tgGxWXT1rE3mwmZZKTPYqM5MGn
O0PhQJ8PjDafAcrcRj+1ExujzPmb6q2Ivt3gItmEPl/QsCJPcADsFoBxttvlcpNZ
sJIEVTunffM1xtE2upVW1qzrU6OIuL+YrugI1hny4ss73F9qYikPBFVz5nG6cnST
3r2RE9I8yvyVQS7byiwFObe3fGb3DWntRLlSvuYSANbFghbk+N2lzqkIbgPj598D
C6A+CWLw94taLlWJXv2W9xKQP7DWrNjQZ8iO3HDvE7s/M3hsjfm11YAKcLs065bm
sW6HZ2/ZcDLfXhvSoLX3iloWMF4IPLv7I7p3udQQjzgjzUmFk6FsptEqm5jLS9FK
viYsKqrSLVhik9oCCoZrJrYyhlm4YfY6jXcfsFMvrkG6WqJSXkHBfV6rEZR/EKmw
elzR6Ug2QpN0ixFTZz8Ey+xro73U6GVdmBQ4P/hM3QFGQ/9X5l+pJwjcz2wGEwR0
rC+TXY8XCJV8LYETR7ruHG+4OHwy5BjQ+bpnry34UX6TY9lfviPBSKwsX0O7qw+C
G8pR9umxZ1XKKa/Or7oKNTAgcblmTfFB6bGKLP54fiecaZ7cQ4EHGdDkdW4iedWV
pnd/VO6i3NrwpSpT30/V+aLYXsIQSQtJVEw4FEIvTrgKlJlJekjgzEczm+050QOu
BDj5VqV2jVCZuYDuRrXLV7NM7N+Thogg0M+JBRvSyIn29vNS8ZOa0Yf/KrbhJzdH
RorfPHU8k6UkWjJGbUtRMflWPxKw+/6poY/TkVf+lP+k8NbTYP+IdpJT61bMQE5C
C2ehbMu0Hj/BFViy1zxYi97krhRFMJ7TB0hQ8HkdLyiRAv5095TK/ZcRs1I+6Lmu
OSVdS7nqidpQeLNlEj5xv4WcY5cl0R9sKxxdfb9/bbVJPaGH18PsmjI1764KP6YE
grjvMkxZYaoZfTneUa/sUVBIG04PmEe8x1L9Z5duGwr9Gob9XPpUa/OVwqJAvCiE
QsuWlxKOjTRJJEA3kQKRalB3FCa8PRf+rQ7c/bc1CLaGbAQj7LLtxd6ZbSMf9bd/
xqlNK83wYrrbl4AIbu2kxKDgkzbmk65rEyx0HrJvyGxtMG3Zbp/QEm5LhiJdJb/N
TI3sUTIMiFEBajIGbDj9K9uLdFKWLZslZ3NKWvUHlpCQkZeIyjuvw+dwH4NNGjMC
/Yq1ZRNpUWAYsKgujHlyKu+qExB1xv6HIC82IpW7dLcI1oTD56jkBhBygX4CXrn9
4b3DAf4HmWosIBhBgvIylYfR0Cr1BgxNyULBsK/Z/7KXDDKy7ZYvybKv+Lg114D8
lX+gMR6nLilnkCx/2hh79ycuk/Q3NJr5+IayYw4C/8jqC7dxQwGpk4i+ESbWK1JF
6zzX6CgPXorqkWj+FdDPWGO4LCcRpr8GDn4imABvTLfAnfnOAdIiq0cDLOuBxn3i
KNJJqx46uTz/BuDAa7fleLlk56dATXoo7S6wDa0LVj9fAKFlQBDyrbGwe/TqyDfX
GwH5AoSHrrYegQaIzS6MtYNnEeWIGCewDQe7eMqQavFheC2+IwRDYGKTFUstFc/i
T/t0KAxG3PyCOlr5iGLsRxrcT8WlqcyO68KEdz3CMLWwKX00okkPZBa0xMeS9tWn
A5xYTBZIWkPkHrMdAqdVj5BLcvTx2e3rcewaNvyhywcMCC0Nn3IHX9j2xpdprSKY
jIj+wsQ8QAoeM0tfDTe+8/l9HzQNUOw9ZO4jcYrcVn2YEy43HzKavySxQngy6gR+
9pzQfKYUd7dNe9Rh+IcUv7tFUvEaBnM1yg+G0/4CCQ2jPacW4RfRnTh4ccg6Woe4
HvEyjI0iW3j+GczDZug7qE7B7yH+V6hvfE6aOWv6/EHTTP8uZgXI1HhB7XdsNy3E
RY4Uh5pOwVPfgpJ98Cmbtwy4Pne0i4EkmYlBwyvg6oAhyAfpMTt14mpX1hri9rEp
Kj6peZO6+mlpXoMyF+yx1DMb2x/RuMkLuP1oOButBmH7Y+7bMEt6+4yZGdK3zeoZ
+4vjNembeei6TGQ/MAFgkuCAhZ38vWDcanzdXOPxE21RbgYULdyJsz/tXBygw9B9
ENMUvbg0Lcod3Y+NkoeVppb0NnM763IWjGiFfzmEWvAnIejpFAee843hi3NdHbpg
5Yt+c0EAISd2q6yN/W2OhnxhphMJR1l5+Mrw0UZM6nWPcaZRmKR5JiywO+Frc61F
0bC0FDw/7cRdNbXvZwxjY0XzDJmkPgeuE3usnOLIXwg+KQWk3Tf1E3elTahkjDCD
VgqfkodTjZorzTh9/I2APZGzxQ4LljrvD9ggyrs8D8HmqYcw2Y4X8qzkCwwKlvKF
vOSgdJT9NTyS2GKKrEg2JaizzZR0t5xahsD080gnsntkO829S355dw9TKEDi99R/
O/TGnklPhBnLrQQ7VVK6SbX/Pqu151R+slOq2DstaiOq4RdRp+4wCOglDZSTPQCK
gcimMYuGFbFgKhvJzu33iQs/0efoMtgm5MAmWVFch1MJEBvn1FdIqVSaAopE2cT5
/qtoog3VcNEcc72AbVpy7+KJOKKMRqzhv6xqDaqCcLwEG/vDsISA7ua9MLI2X0c2
j/45anRCJEgqiVgG35kGfxS6jy6IBVV92pW0Rrgn7VbStkqInECf3lEddJunVquV
4MRAf3UCoIkYfvC/4843I3Y18LCKd5rFLnyYIMXFd8XEhLMsXd89J77rL8Jf0ejG
0AYjFeEShy9wy1G4YlbOr0hWs+3Uy/t3dlTADfFsBKnj2boiWPU+23UaZSxoH4CD
wjV4D+H6S//7hYfDmjQiHl1L3iMah0QM2WC4kVIMbwUNmSKpOiYS5eBIy9ejuJnY
MHf5WRw0E1HpfvsW8u+DVyCBCqBymQoVQTn9m7eKzhUDDnzadxHW6nTQwzju19FJ
EbNAiBSod8+YQaEKiwGkvh6J9uUProLPe6LJlB1myQkJ2rT4N4vr9awuwzh4cR8r
dI19JoSnA+jWXHMz0Jd9iXwoih8CYxU+pGmfDKI9W5fQ3usqNoCq11+YLoxz7Ww+
xaa5udDf5pgb3wXUodf5S6ObAZDJc1bxsdy7GkGpsHFulql4CrlzQ1FROc6dDqqA
07eceYyR+iBXF8vsHQwHJ2dAn3+nyIityLxEWiS0uO1wU12IshIp8VWpMNJhrml5
hx618qGSqeJMJkf9G4APHTyztUXXFyPdRkdyEzh2x75WamhzkMyUbcKF+u8YqVVr
fLnmk4bRKI5W4aOklt2DqjF1ffA4IZfPKbsJ3dnXxJnwvRIh1z2DA2wv23e13e0f
k7iBwBpaWfL77LHWPKCuYXurMIVXjiIjw8kQsheWtM7LvP/t+qKTBTldO0hnbHfr
hPWHrU7wkhS4y/TDBRbBvR+ceSt3p1XAel+/a9BCSb8SSBPvlBKoXL0YcvYnjt76
+7fl7SIapwYm4i4c9715j0+KyYelM0OjRgkIDW6gjz1ZWYVdekSw6pS5byiNxDOv
84jyzxP4PffJy5lEXIu5vYEsXPJPNFPeEsjR5JwGiswV7bOq0/XWMOL+xGJ2tcCJ
Y4sIW9mfXcG/pVTnYHxFrioj2U/rRlL8rZ7YE0hPO8NmXzjewcZhdSnrUp6KVink
NyPSkm6LTWJSoyUNaNm+Tv1ddhQ6PA/UuILiuCeD+dGDREU7G54LdkkU8oIL9fuO
jwclsODP3rfbQg4uKMJibx9DDFtPCJypGVZFprBHk7ixWXwpaHTI/saFZLXaeWkM
LRcnHJ8nc2xiC0pb4lezGxglQYTXqRXnVbQLZup5m1VhOrBDGoX4v7oL1xqRXSXl
vasAgivLtVc3ZQp88LWfpukJHKWm+l2o9WqRlvz17voT4hio/r/fCAAUPKKuYHlK
xmW1l3+pmN8dO0yt/Tds36MyMw39CREZt9XKH2uaOJpOUHoT4kSYMIOG/qbcVS3p
PLmMj6FUiE/FSBKvhupIEuA/rEUDNV9Xtpx3h+P9O94rDntxz5lw+15SfN+q8zBE
8LsLBSvhEy8wgK0vdkBaqXZRL4AUZDQ8RsQ7VDlHw5FnRdyk/Y9AHBW3Nf1g+cSt
JNDNyaV/PH/YiBTZdRHb9WyKlgQOpGxtd4iQ3UUoKOJwrunhIcXrbOUbmIGlDQR3
PCJHGN4ohH2uohDO2/Ch2FACWFu1QQPaqVufof4aWdy37Afq2VoSx9BN8rVQnXiz
1KQC0rdVIrnDt06jIxChnJY4pRdGDprKXX6Ty/uyZMWG9CJAwxAf56i/QKeaOSND
fMwgcUKB2fGK74nR+L7lJ1tdrfyCFqqnH39TJu1h6Ogoh9OAYxgd4492HyzNyPog
MPv9JZ5hzSduHXIQjBQoyr/Y84lr7vHsDRxpCc2rLNU79SjJRZY+vp31C2/y0/wl
qsEeahHCOgR2fU3JvjdVHMV9viSAGEeQ7iz+ta11bZc8m3q0mV0hvn4BWLv7lJSW
8CXcUVEwOF6gTqSvhYJuUfiZFnjGx8qn8J+kGmBHl1i1PGPgzKSmSzC7v12o4i6G
eiarWQqqnH30MTZ+GE1yj6UcE0SXNk1a5A50tH4Q1fcvjYc6D8iJpr46BwZKECLk
lTKVB7J/1N5/WlM4UleobJxgYdx/eyItjO9t7qQNFeKOiowDlc3ILIbalwF3vmKW
3JM6qoGlpq+0klTKqIS1URR+ePt2NFOUErR+XOcvI8aBOT3evU7qTwvoBTHaCcke
2qE9MT5B3Xe26qbKLGiXLnbsuLePK26fIitvDdyCFYoNpch5BJgB7Sd/csB3mGdG
fsfjBYWhH9M9zwMiIQXKG/diewxQvdd7JiirSbDgOuaNFgSJPwWOkkWMDpHvkzCu
+cQBzQxry0yVBWuxRlxOh257wnncCztW81InNgmsFsawuic5YGTGFOWe13cnvUq1
Q7E+sCs2Ep/a2n/u6OIQhWwveGPQbbBsa+tezkE7k2qhnBOwD3Jj2H49PY9znxIw
vEBiVfddk3WJGGhPS+Fv3aHWigBMnG2vM8SMbplgvNjVpE5TPtZC/lpaMdaX86Qe
LKIVXY7pgjGYaVgkRqkfzc8jH55LhIKZS5DEtIFM1s3bC3i9dr0Ep2933w9v2zgz
gUcvMTPCRHDXq7bjuPqHToII38C2CLAALg8LPufiZIXgvmQRgn/vt4muKlaH6qQi
2eDy1RAh7OrVe/3EiT5XHezKGurkl84ymqgIh1BOZPAPTDiqzYKUDYkIWB7QATbu
Mjw516l8IhNsTeiWLrubBiE7rUlK3BlocuH1O4pq5QL81+v2SKO9Vs4mTaxCxhXG
iAs7y1PAhpcld8+9lrWzFlX4WBTvAyzI551VX3Yj0+cTZW+2RfSfNoYlROSGfL2T
KT/JTE5tCfFosiUCEHIn6kzsqETHbFHbsllK6Ymmhc6exxo2YxjYVLUmTvmiFW7X
GyVrwlXe+xUtmPTjv5YcdWv0zlE2EKSq8HwfLuASGgEfw3Ng6P72sIwviIgZcvbn
BNO+K2BG85vHVq39BPdpr9xF3Nr4Zvg599PBh/E0OOxd+Uwnw2qPbkRZWHZpOB6J
KqglyuSmy//dKiRnC0W/PLOwA6+1Gv05DQxyCztDcGlOut7a8Uis9SmrS+WwHk11
MQH4jmQi1ahxbQxJbBA2+yvRart07oNBctcnv5d3YQVULBCM7DqUGfyS+Wjdz63M
EX1DLt3dACCn6/HfeAOSq6/KAsh5yZeDBmIy7Ijcvpe3CImXsr2//iAdQmIGyhkY
+94ypRC/uebwgjq0pHlsQmU0ac3ohI5WnBLgS0A2Y2/9wou2J24Ne4LF07BLXyGX
7UpUj4uehmGJNQE7ODy9ncBpK2YQF09tLIR1QhcXSinU/9lCwQkvnk0/tZX+AtJv
AsD+8lNt4QYgOZjG1QWq6Wn3GS74+2ftjZ2VfbimmhYvBC/OiHd7YB7LOi6AA5va
PuKa4vt9oE9rYIvHP3my/d67t15g0ow81pQzGuVu+gLw3SjVKuFhIpYPbGGq21QY
yiByJJQIneDDSoyRfrgddYlMRrpW8/olJyh06zMhUDyIMOvPFYLATE5jU1mofB0o
l+/vobAx/ibjbBAULETSMWtW+Xi3/UGlgi5rIGKInUVEoZVRbr8zH3Gw/cNBAJ0W
uG33ydC+FOIdPqIF7e91cxdPwJyXwHNBwFTJFdwu5fYDQ30gM28EcWmdSyb6xNMR
6+rtZVzCq+3h/heUF74MndzpbXOJqsBj2LLh7+hznvNkcb6M3Gq8I7ZcBBZjNOR0
B2+96Mgh5OefMAnTh5d6XVXx5doqyPkIdBEhDkdQ5FMRP0VG0eX6yHxH351muQQf
FwbENL8daCvPubtsxy7CN+lMVzZBMEr3Ne06IQiIfDNJI5vUIRrDybksMRNQDArT
jTakZgOEWu4nkWUvQpkSstl5gVCksZcTI5uGw/rdRgwU4tEnNkrzUW0pPtZ9jFrZ
6DBMVO3tubW8FlWZP/dOTyVu5lOBTrpQXTkBkceOR4IMmeS2a3+dXqCMpoVqyw9P
NpKDEKUZQS/11W6hCBgQDQ+erpU9P1kIsF34WlkU7ZbtCc6B7deqfZQFfG2Q+s41
TClGE6vult9w7wKaSrmsLQtAhS3HzjbZybfmcdZ/byCS/8W6Vm0DH0OAXjZlawZA
fWKeUp3g6sJX5vqc+KixNNUNLiC2q5jumewrJ7WnRKRv5bbUy3fdFnumDnDQRs79
qA1C8kgfe/XkqtyK8D7aXcfxaVLr7lWzQ7Rr4JCM5N+YY1rSlLXP4EcNhWxjpppY
BX4JeKRqieV9WJ9jkloMWlnTjcPdnjWy6UIASHCoJG8bTwArnc5KofoN6fj54IM8
gDEzPapM4WfE5u/s+48s2qNcp9kRi+qdLbEImp6vUdMcRFp0sEn/r5XWIA67vazw
sDQMR/0g785kU15bCfHbzyfNNvexL/NwOXBfLBQkn3e7DD8ezwF4d7r+ISqx3zFZ
vgUmMqytTPj4FXTFmlrNi3d9bgyRQJjgI5tm8f+uqCOGpRS/6sqU0Gb6dFy7dBPq
MaT+O0brFBCScUYXaRZof3FM3Nwnvl/8MhDN8iJ/N+1BLO9ULxQzyBN6llDSaEMS
YE48lPrAfVJmynyQZWnSm6ptk39U4RFBxAI3QuF2XSwB3aUW00Xd358FhKyHEv7b
4xi2Fof6k/dfFI30DfbbQAi37SwbmqWBeaA83QE2/GeSF9QzV2YHj9jTgso9c80s
w1HYEjuJQGM5NpdY9IrXg5X7kZFmXPTp3h4+0nhcxy8oBxM0DTf7VasEeb/jxN8L
57ubp9tKMmVf2c8b7UquML/hSaM61zmovFjA95E7riu5MYVZwWa3NLwey94CcYzW
5RO7nrUs85xdpVphd9upTqcWwJ0Mg3luhZYsHZZYgBpo7rzTiXBmA60SqZrDCjuq
yuskXx+YMvHyU2dn1C0CMcDTR6joSRFVsaGToWtuUVlDZdMnWw7gpq7BFTFFk7Mi
tlUv+P+rHRuN/YYufMg/XLY7QANcWAQZ1SwwCp6st/7V5QYLId6Mz700iMj9lbJV
kZrs73yASvtuAZKYKT/uumkAjjyaXH/9Ymq8lgfNKZO3PIzoeL6SD+B+b73ZSE0X
QJdHbaHKYQZ+nJ0CUVsOuBwKATLhU5qsM0C8RIH9P1yf4dc+G6B1N2ss6ezY+MtS
5FSGOj/BrGnXej7BZqMofDKcevu4T+mjuOG9gvNGswtbBCfJ4qy8lefYHtxW8E6c
yCCVv8oQbnWc3xjeVqFALyVxoesu4rJFKVne0Ai4acYGWcEeMiZdIzy8lTz9lzfi
lq77aUdQtO5K0vd7DTWl2UbUSv1Id2M2IWmy/u+LWS/25t34cB7LfktS8y3rOrSs
YL6aeqKy5EfQ27CRSlie7Y7JrWskfjXA+LirYm7RA34EMc2F0sSLUXazqLNSAqhw
I95o+nMzUK69Tk68I1xOIJWBaYiLq6IkzTEprt0P8nx78IS0lqDqnbBIwKwTBoLG
oT2/aB0s+U7cAt7WNc2naSCdwFNeFWCupNA3YpAVpWGuchsGK42sMJs1shdGAvg0
tdAajC1a/3P0b33A7ZW6suDiGAkGkBfUlMdKgioMT+xuD+ozqSP7Edg874JOokG2
jsFcB72Xz/2//oBrL3kL/PRnKCaJXYtxfawH8yKi0NVQqPPoY5ok2/m7Rr/ZYu3V
msg0a0lSW7fEQySJl15E3FCgyksRWXks7Obkh04ASHt9zhmB4AIALTkw1zhdLv1s
G3WOtLRoV6Rmg+CrGBYvQzEYgsCMEiBwkl9ZbTAAQ3MLNnfG42BT6dR78Rh0d8Wb
9wrF3S+IErzRuLJJS97P6W1EH/EPD1gWrqimbi9QduNcboFr0cLMwYVn05293zin
au5vqLrV4aYgRtv51Yxgp3vxcC+nnHLqrsjYJtuTwnXQS+PKbRU4yCuG1D3LVSWz
OTkCmZWxgi7y49VOMaUyeseKPNDPyrkGrsL76aQyqMIpcOWwRgfX0KtljGmPbtJ0
JfwbtTR9GFXyEsWiSH+AjKOd071C+nmTUV2LSmHVTdYMfKP6f8SiPlI2pDhRZ3oB
eGXwsmwzhw7Ir5f9fLSjyjFyEVUxgW8AmKj2h9C5UlYPa35XBJSPwQfs/61xuPcG
Qr1JEqvpE7GWXkiMumkJbu/Ae2vE2CVziaZ+rpJt9d3Yi8fTSqnCVP/ug7Oz+212
+FE9UoogYgP0qAPESLtoJ6ABE80SahkNthwTLX7dmLNU8UfOXcLpFd9IRFNNNpfv
eUfs5IUrFSR/OLage4k70wiX/yQGSmORLNZkfA0wBcGloaUimYn2wEodHn4wEgpG
bHQpyqfnMmiy44SfC6TuoQ3SBivVImHwsCT2wm/l29HDv2ImW7+iixyORMVwy3FA
JI19qC3H/z5K4srsL2n8NKH1rxHNgMHT592BhYjUgqonQgCq3vs60qL4Be2JI7Pm
IX1vr8BE/v9XLYfGmoQhys6g0IKgCI9MVZRj45BDCBh49MxZ/t1eehKoyi1cPnMj
n6H3C0Adz+45aqypKCGJOFY0VGwXPwhfnocnXxvmO0T0pZLRHU+dlzkk5oowcAXM
fcPgQQcu5xjxYcJgjRHgaJ4L78pLrGD0LU6avlEhTU9aGEa1dhDof2zz47JRQ/n+
4wXRmeVBCLUcDil5yfKTw2OWiVdAUTfV1hNdRGn4vFJ96vpKgV2sMENvj5wEb4kw
EEuvtC9kqQ5WZY1q/pBuuvXkItbyr5HBdKKjmfOKuHIibyFM5e8PmWG3zJGok3Ww
kpv+RC85D0AziFPoGgWiKHAtYGGPpCugf6hqdGt7YhsUrySfhcszuQ1XZi2pZ6dv
mj4++qwz+QvW1DRzpsxeBebjVBvFEyTIPLXyLxsOcVirUzDlxFZSeDLRfP3Fdscn
GmR+alqfnAxcq+PaYvU7NttplNTpWSiPhg7dEpxPAL3sOY/tFSgZO3u6Ki+Y1CYu
pIs8mm/xniVr6ow4EVygkGWuzWnw1OOdEQ3OgJ6izh16AcUkSkVoMKPqnlC3yL56
KgnZI1+6E4DPD5sVpoHfSzbdsxUP8KgPn+EUpMoXYIi6Y1ui/SPsT/M2cMLHADAl
/7RLBp7fAW+Z+6jDCEaerSHHVJpUlttDJsRKmZaq2j+lif6/qQ0U7gR2i4lHeuZf
CaUL8lDnw24PX2JmzTRVD2ABTv0Qg6BJK3hwS1pxg1XRAHyGy/ucYABLxiU/ceZU
9qpcTtEzFZBzC8fgZWGHv/EwKwK7Leg3dKwuhaWIQHPKPMINMuu513W4JC4FY1k8
PK8AY3LBiJiz7UYGLBLnArXfJDsRraqMRDw2IGtifs+rvCJv7rPvgyQcHJpKjf9G
DO2vLpqoMaRNvIXKVT7p41BFobXtyS623VVqZ8yTUqEqil/mRS54ftmX8Ou5mHLI
my5io/BC56tgmO7th4Fg0IShJDRROLZk48M7QLc3wXU2XyHnYeYzlaWJ5nndXTiX
lwShl9g6MmisH5rKqrIHFin3pIJMe3PJbtBOURvA9OVUKF5pYN+16a+7LDf5pxYK
rNyMKm1mcpsnjC9Drn0AKZDnWUHDz10uk0jwlkSYT3BU9K4q0JPd9ltOZcGuEZWA
FahOuSe4ZGvycSvnM/ZZfsLUg2Ba4WzO8rMu1Vvm/1REasFefk3N+eV3NEhXS501
WgoK80eB2O3IXeu6Psyjq56RhyjxAbxVkCO6ous7835Bw8oHENkCTXT5pWqMxjWc
wY4iLbaPItHF/2uPD0eiYv03b2rqAy8LkZKeAszHBOF9jY+dEyjbdpovQVWmRjvm
B2NZPkrup4OUOsuPWJ5J2E9QM12zSO/GEzi1YrSpadILG/JUUGjMYbnQsut0EEXn
epoOS2kT551rU1o2q/H3LBws8fLNHKrjv+ho3MlNKHmNtwrfCzCZ/MmafgdIf0XZ
aUgnquq5NWY6qtamkF5iYjDi8E6VIpn5vTLHzWQ3sl+2u6YkhevhGpqcbZKlfVGE
zZb6wPvJafpnZS+BCGPjq5Fvv18OPCGu5Wo6yowGYFeJrUglIxi9rrHu0g8dkF0a
MVudV0V3V9IqpBCOoEQpNF4G0kUN/+ltFIChSFewkeC+HEKw2BhgAyT33HHDiD13
5PGHRtq/FKEkOxPjhlmLFPNmFp5ws9H6SrtDfCW3yJwwB1djtr2BER4ZeqG2oGaT
0hI6BBuUU5woLGvMHUzdhitGbYatLOK1/H96nNSqEDnK55kPQuU9UIqbWVn40qZm
PlNKQy34WALLEUfxGfi7RwkoNmrCsFq1kv1HbrYgQjGw6GimzyKhUFcpOjiI8xQb
jr6N31XViIsWOrzey4LyRSxcU9o7MVhOX7luJp57We/hgEw3Z3vXIU+DA9Xn4d9/
ZNBO8iDwxsNM9GbVa9lv8ZJ21cUHrlb1UMTEOOmN5F5+mlE2WZhRsVsRNJB3CV6t
0XsuYGNquVrpj6CE6bRD/m0RJlJrebQd5RFmrFZUSy6Z2vdlI5hqazfxnfL3cLg6
G+kM9xMYGxWJ71l00gmjWsawUTr3ZixiPLFERQ92J9Swkcd8Q3mhHYpQ+dYKtkgM
a4qDyodWLFGF+ukKrVLuav7rZdGmM5p6D62SXDK+vdhkICJBbzRmmr+GHof9e94i
zwiTah6rLF6FiBrUuMzFN0Oa3IXwl3p/9T8o9StVMojhIpNTQaf1g+soyMYvQLw/
YMZzdmTZeYcYNBHaMxhhNjdX4V/6COh1dGlBcx/zu+NKf9p6dpL1BJl1ZC5SXk2E
ev/7JrAIJK7rAT5Vx+6IVxJ6dzslJVXmBoFv9zVEA4Pd68BzWDpmZU80syuFr4vG
x+zCZVf1+TzzTE+KtWLwtgRctOkLczZqmMqggMlCDmRRNp9exv4qeLIQxpLWb+Br
mmhNwSOvDqm04UOzSDv8NWVTRh+dZ3CuZdF7aI8lgUqrM5gG59m9xABb7AvXKzhu
hsElZxTEROpEMgQRWq5MtKzQcIija3KSd/A0ja5waoeUDOWmA37w7tUTxjfeFCtJ
y5bm8E8pmFlJ5HOJPiIY63mg0skIquWXH7BuUBydqNwsEzVv7zCSa0MksynjaoHO
4Ud/fknOrZFBdD6Cj74I649UkfPhw6Ji8YRRwRAPhSVDBbCbMtfb9klCPT7cSgti
QmhLCDsK7hxguXtrjuc8bdOCRqAxripr9E85dK7v+W8Mt5aX6IdZv7IzIXz5A45C
aZy6BJn4GBe/JRMhsWR8R4Yc1mM9CqoBrhRSyGDvLDF30q9Nc7Q2nujx1dsV/UeI
ezqQHidSYdqXM3rxrk6UlKiYSXJh5w01v9w2+zvQNhBpf8RHa+loErwahj76KZ4v
jvZznA0c7xT1X9j7ZxZG7kVkIWO3HORokQiQFd/wqCfKYcJbe9iSxgYMdeIMAQKc
lNfrHVP21sy/TC1NaRImKKgL1vKzu+1R/KsifcXoguYHIh/j0QgCr1/5HiFKHI/q
X6VSOdXrbBzpLkqKAB0oceDCKXBDQgXGNcHmGSzKxhisr8Yy/yG9lgRynNxX0x0o
LmRPxATxLbumdQ4QmGMhcGWinx2Q5F3o9qdKF5A0HFYKOJdQirK0R2M3lSv0UcmE
KezENaqj4XEr1vKqcvcnXpbVwqA4IEPS2+6CizBGRbToCjyOKDhYvVlISz7ZS4OP
T/67us6keQ3ki3gV3SPkqUkzxaOKqgE/5JnOl5W/DjeIQrly0hHEWYatIFxd1LRl
ycQ8Qpe/8dDqYXMeoNhuHGMWevU4x8yqqQr2P4OICk8gc45iBKTreTeKvmXU9utP
xXRvp8v+fSzFauu51qscX4MEQOcGRnPW0/xly+JWjiAPLUNsOcQ/s3c2M17ZGdeM
zzzv8vm3Qh4csjoMj1GU54xMoJVgGqLF75jiE2Hk0WoWvuTMZHeZ0Ryx2zHI2OcP
oO4fpVOqM3K1Crmurbc6EjTQujyKxY75HnRpL4El3RRcdRp4o2sDWSJkaPb7jIcy
JTenRKd1zAM2Q5AR7KGbQKlzCLu4AkPf4qG1OjDYz+uFXbMsdpkPWO84UzjLkIdo
Q/NxACZkCTGBbVlLBpWAiKqEw6xILtegypcaNbCMOYyL4yB3khGyvF637XVp2EBL
ZCsMc+qzIytLbAQKgQNmxBfFR5iAwMcx9miJyu3f4fXNbiGi16POdSpZcDJMptoA
dGVyH9JeYxVKXgvwLR79kxjs3StKHQa8vBLt5ENrBm4v1L8MzPDLJnb9FPtyLoPm
IMi6Q8qdMAblNWxcqSU2PkX2mCwskrg18tFVUe6di6zTKKjFgiVQlXFO7akpcuCf
lH2n3IKluC7lOOAMZKNxAH4C913InyxAsIeKOGmY9q+G+YZ4pkXEm7B5ibc+yeRJ
/RVJi22pdQO8ruHe0TapNlvQUlJt2ys8kNVvmaAXYUmpAlR1faFr372QaOI5gVtX
Nz9tQz/xPSsFL06GDXnm/QKwlIjMCdmAQGX3idSabJoE7Xqsr8rUUXeMUsNW/SvJ
aZJRfpxS/svspc4omezblB538upaoxjIZPHA1gr4UfwOVyNfC8S/xjHie+p9IU6Z
4LXZLoyNYXasBBaOquzghoC1Sf1SDX5gVeZrylcxU35YsfwxjQO9AcUvc3UbZxWx
Def1DIGPSMRt6SbkhyrCM+GP00wW5QaPxd8mG61dMvBOzUwgTT/rIMM18Y0J4F6J
wbR2j0ZQXxFRnHsARjD+zFSiY2aFH1gBpMH0R0oyC+0NALOzLz0yOKJCQs74iICf
tSZ09htpL+zsot98OmsnPtk0+mFgzikmqykKs0oIa9H96be19zcJd0zhFjD8wlFy
Wcop+0LkOvgolL6o0iQG7RIOJHeTZ8cOCFEY7GbBlPCTcVMKvw+V/FyULOEyb+eQ
y3Slh+FDpX885dvaPcNa7tcGSGA8mzvTdvXUlFSJNzHE90PV+im8Jj0ydxpaOs7H
r5FrzFwvZerSgXK6NhMAIrIqQJLrpaBukqkw99JuZk7uACnnU5EroW1XZ6xeOePO
gU16H3XbJUUi2RO0IJ7syVo9NyuP5O2zV2hvdq1zSc0qbp34gRmt3W7fEDdiJYJy
7vquqXPlQ4TxIrxjDDomaA5NHy58RcA4bdGDo6lZpmkcNxeAR8Kht7EzxWZK5Gh9
P0+dZsZflcPrWdzJNTFP46UKCzdNS9fI+XT6DKB7q76g0EwwdRUbD/GaesL67bjv
XzbdEraCQRx1KYeukLYzGebttp+9egJGIAmOcHPIIrGsiVm6DFfBg0k/VcfGL2Fc
mCRZRTZTs+nDiu8VTMtsXlPiX5R9KjWqs6SV4QtIkm9DuMU97mhavN6HFl1PttC5
nByA/AT5Gp2IpJOI9V6f1Tn1f3+1V3VyKWRK6XKF9RklY9Po7F4l+q80YuYGpONn
TM/J/c3haYHiKParvWy91s6OfE2VeRpomt6Gs2XpU+526plJ9KpY5rVklN6S16PQ
h3vAe+N0sC1RJ7sXKiFmir7k/2+dzgWwbr7T42GyhQz+4KbThOKzlwwRxlMWDjqi
8418tYjpLCoaH8g7hwtPu3LY7Xuila0kq8UEWfJJhneUTE4jBKfAOYOY71VPmm4U
bhjoGBgO+Qe7y9/J3dX3lUBwAKSnN0DIzkNUFWrHcnyG9ClnrI0rYAi9/RymJvcw
4Fa+bRwnFsq0As6IpuOqj348ekb5E5aNAZiHt1CWMdUWKwQW1C5tj3VWH0jSlNcb
yZgmytO4a0jdL2o77EG9hoBuLF77WV4IZLS34G6cp6nP87o7ZU3oCOhQm4ycr9/T
54zAakXs9c5v7kRDvlAYigCUurVJW8hNMNmcB11jXomD/kOUfh8bOznD+mB2cN3h
l+YOAiGZuEeFW9tNfMRk5y2kjOHTQr34GLamdfnI7W6XHN7Jldj+1GUEqk5kdLXc
ua6eIkVLzIm2dwqkPY2AC/aJStMUo4GS57dRxSl1qoJJ/BSA4m0ExlNFKSVhg2vo
C6aQ8rYyI/aDfJzqx88VlCEITZMShejg2j/mexhtpjA6Dkc66vwr8kbfIFOCehSL
+lXDpX5ZSgXmfWefO932UQnYh/zvI4rGNZ2WDI/0jCUZWtqA8f0QNfhJYHaYQugy
Ma/8kfD8l75pZawUDbKS2DOJgyLHm1kRkyiERjVzR0l1q2dmvUpRKHUZcnR5haQD
4I4fC2d7BhmL7wswsFWNpVrV0MTPaINQZ94CCPW92V/ptDWixkJz6UEiR5PwwHK7
AbCQJoIjJl14PKGsiLZNVZhgAmw3bzWC9WVn/e5TEJn1gh04edNm5sL+MES6If2R
9Z2PR33GZtlorOWiKlTeR8WFlKqPNBvG+5tZrK4pkfiSAa7DUJnaLOPofV+C2QRh
3eqVjIUDf1ZWYn2pXhXUuNuEb7QMSC5msKGGdhj+9womZ2eLtiIFb0LtJ9huaiRH
/zVRUmO9saA7GRePhSYg/cyemhY6gVBCPkBk00PKsWVD+D2nRzx1FUWz+QNxsR+e
dbhfFx6sUOo6AHJLgfzaQZd8z8h9aFex83iK5lTgMXQmVHNr/qWKEvkZwThhj/iD
qDa9zlqDLa/+SYELVGh6GEGAMctll7t/W57gArhTiJzpq11a3ubfNd2HULMJpYqj
ar+K/uWYVUjKcnE8XOkkwdp8VG3O2/jWXNJh4Dn2kVhfYWu3ZfJPSWKo0a3hkvuW
zHNdHu9rS54PVv/HVrHQA/bwHpzMtOR6gGG9iCSbGzNCnkm1k+04vRpLCZu1jRdl
sdMaU7Ib+bjluIJlm7TFAkftQGWqXsx2LqgUzaw+g2tlZo/kn8GlQuQLTVYJVq/i
kXnaO5AA6t+Wd9fTi3xkwHTU1QOIrdVzzoRFdaSktXA62KWYwJ2wAwwlumyTr7sE
cuSqzXKeocrpeas6LZaqf01+AYN3+Z/sy+h2lmkErSaVE6cORRLf90IS90JPEIUb
NPbv4/PGzKmbNJdgoByeMew0DlhAaekue0hXIzQDrrCgNcBrs0EJmHx6Q27+YALD
lFWfm7um1fsQduajCd7/lSkgYedX85IlOjVAUTluk6vAk0u6rhYn6QRRlKAx0HC/
GQP05AvBxvq6KrT8KuiGEmJlhLbbY1Ax8KOkEv4WUToVZqPoguk1VdVBPjJ+bWav
EykolVEZ4hN6KDMz+UfedPIkrSlIUNteJQTcSSiIawXp7jfiWzqpQ5Rok1mgvasP
pjX33XE5QD8I8XGjth2fC9QJ2tT+vznoce6hNJVGQFnZXIalPzEG42PhBCUCMSlq
w24hCLJ5dSlNP0jCd6XRUT9dyFk1jMxM8/6KRzrkMsGes3fRESEdqGTcN8cjBsfR
v658wz9QCjHvwpzfZrN2xCeIkbXgd2hnFVpDd8N0lrGrHZ2isaDii0bKCSErplTW
OWYBzaGhN0VHY9vRi7EWiRYA2e4J+UEeZoNUijJa65mPYOl9ravadJwDb6cHN0DU
kiJOHkfsZWiXQZDx+iuxQime8dtyeseu4WcDs0HbZnJTa4LIH77oNkIIkWgJ0Afg
S+1pJfZWNbnRM/z1jaH77kSuP8Qa9+EUf9Wmxn3BcoEvtNU1/JSYIWMc1xD2q5C6
niyzHm1WjQWY0YBmUdsGSz1DQAZR6NnCjQixW5I+0ykwXz5SAamQhhikuz4v9HRh
iSwa8FfomRzucQvVPNiWdt0RNXi4opAX2CqLHzu+eTUNunREyIcFjVYU6U7x8dpO
wkYq67JSht9SG+dUFR/bNsUk4xKcQg6V2ey2tYMljYAqaOzaCCQ/tVY2CVT74NzB
t/v+bjlCsOVTvIFzCJ30s6Vjqh/2ZzhBH7Et4O6vlOxBRd5obTC0iomc5wgf1x5b
TEjLZ78Sew7TT6WZFiIIUMe3oRzB3dL8bgWAdEoY+lm2O5LQ3JwlFUXDX/SkqfrV
OtN1uXf53v5RRx5sS5Nnlh2VcbQ7MeQNZPDIgMTffaKbANJV+vgmGjSc2onKTanN
XL3tRi2ufgvsPivTdgjKHjqu0ldUe26WHvk2qMskwyDVozBVIzqrY9m7Q75zG6Pc
KR1rnAg1X+wCZfr87X49ENB5gKGuQdPg2t8vpTDyegaVfeXe8NWCW239AJ0m45om
EjVRrgn/aC8XHZKZSy1CcxBtZlkxldiqFNS/Oy17v1Xgs+tvuXVpzwtN9BJAr6bh
Hp3W45IjScGptcMf6xBVQs8MqFdENIHefhjhH6kO1nwBhbndhm9jQTCoyHJeUnAY
vpYS764QaItW5ZEqvk/SLZCFLcf7A49helMSISXA7Gv/tQ3YxEmZfBvTUA3aJ1/s
6l/iPOORgfxM4FsNgPmwa1ZVBsVY9s4NABPWHB4py0EABqJwHSVszwk1wrkL9tHY
K3irRX1ZXp/Z3PiRr2z3ZMymS9BILLgLf9JIv2Z3jbQUtDX/Y0VipPWI77fabS8v
XnJ+y55ebbmC4QVQn8EMXVhgb488KcNnMCqtnPQCQKIhlY24x7UyRy2gsL19yAQo
GORt4blza68gln+blPjh7E8QoYN57gc7koD4jvYiOaDytGsx9blWJfLyolvOoW9c
gXyV40ABeXJQWn+hBcxui6xzUZMpYBElsGP050krpyr/VNkWN6Kec/iOH6vK90PZ
DbuuGFCb2dIITcRRPRL23w7d3i4xXyGmBG10HBqVcksSry8sw7c87pacCNtAl6ht
W6NZ4d+1DuRnOm3bI/Q+ycW1A3dT3Je6DyP79Hz3RrL/cASNTr2ysHiTe0lr1YiA
rBFTAldJVgDBc4MJkNLyF8rqSNtANNj0y7lEVQ/LJPzg8vYmV5qnNYvCkjzHF5Vu
8rlcfJi2puaFYM69i2ZNWyrSzxTlQdIlzXr2T6dDinJnfwd2vWTzQVUxMn38V4Xo
6gq8CXPTio4bObVY6QPslSGrgnp5oW6cR0PCUeHrG4E53TgxHwZf9w1G+E09JOKg
zOQt3dLwf2R3D6itvMaSlCxh+xPo3Xg0xIdQwTCouaUkvGGM+V9Jm8IE5gPkYIXm
bKQrE16CEDjiCHH2HZ/2J7tVS0SnKHVzks3xH9H6yn59WFtkVGBKJl+apLjmEmBO
3vx8SgDgu0qX9ycdzjjLvEm5g3Ya/9K2qUHbElksaUE9m/q7fhD5Ckh9VEmvwKTy
ShBdQePvQTGbINd+ANhJXiqcOIi1FiCKwgyw+QKAQncPFzStEictVyR0MX4RmQA9
RDseoSK83keNTf4pDyKoECgcYvY3DygrCXXH+Zq2cbXzL049e28R47BZCEjF6xTZ
xOFPNbyeTuZf+BoOiK0huHLRvIhTtA9+xTAUJgu8P/xpxM+aaTviIgR9Q7ejcQJ6
C0R2GQ8bQkUPAg3FjWRSuTaTGcoZLYWFgN10TPy9KBPAPVy5kBx3QD54BHG6cwXr
Zq/Rbi0mMFAciSxzeuh8RnwDyPr9nY9h3VkuhykbQADNwAUtfguwMP2qOaDHHmft
0o8vNhU0v8AH6qoBQEFZFP6HKgWh/mtbevJoPCvKzpoCYrUDC5ObR+iXD2G5+mat
flIelKuVKaSu+PmoTq9R8Y5wRKThV6rwPt6jeYCdAPx/+fII6nQKaSfIxPUagAMI
5KDK1TltnSX1vtGyc2cu3dHzPEV6n951pRrp+inHNSlGmancdMqPeyGjYi64ifqo
4x5tn4qMEJ6QgleiMhWYipmkdq26SrYP6DJ2QISA57mFwERJTvTpLBge/XxB0dZd
w/TY9lNcINjleasOEKNMbRuM5I6dknGByOziKvg8N+WycfRWz0azcgn5SO/1PQoG
Ltk1PSUePKL/woRzyVSGa1P2JBDoqtAO1UJzpxeh1RQWmIkhuHDUeOAahND7dK83
fYek1q/SttsqjUdZuWWezfEuLhoTm9Mk6bBTxJRKCJVmlXm5VgCYMd3Gn7T7+xfn
EcQc2nAd0YL/d34QAQYRC2hjmINLyQvA5Z19Me/0Pm0rV11XvnXFXRo29ciKRmtG
Fn22aAUj/CEh05/zVm7OPjByDrWmxf5E4AqJoQCCfAQoB++fpA0bgI3klvA+2ouU
IJSyEA9VDGbi+FtmLXw/P8D6O2J08bQA4AxQud5KjWxHm4WuJnvo/ApnXuJIWzkz
fSauBHPsFDhISXqVmDNFbHSKntw/CTp4aFloC7A/fg1YzZCCwrd9wOHj7Qyex33l
eg/ZHEeRzUyjPID983jJleKDTzEaHsTrQ9JaZstZDoYxEx2PhUWwTfNU2YVcdXYB
ItbmTQ0AFzHXxNKttcmj7BpHOHvBd6Qz+grruDjgvzfF7rlPt0dnJdLKszGxhGNk
Q/zx3/AD9CQpPd3/uZLSQaSv2p06WE2Ynlsn5E38V77PBCtu++qCwp0wdx41+gfV
mrWZrLwqZGdXuZOpPU3yIcZTFjOXJULPyomllN9zSy7x+WKa7oReCUQG+y4qiuK0
A9+GxUNsvPl9+xQf7SCnCAlVd95RKsfgWLweH/5UMlC2oi0jnFNLtSrDVxoQJwle
EgFrP1oJgT2lk+TJ93KJkKDLc2+x4CayHtIlEkPhIq4qdKXi4bUbPXVr0z2fmuJh
+w1RNbQALuT+cNNSAK1S0Eu1wIJWejRU7b98So9nXBoZp5Bfs9p8wwOHiv/6+LoE
2A8NB9No619xAoJJzqOgY13b3S7bdxbIb67OSTC6Ol55r1hWbM1m8e/9cLZk33mW
GriVQN16lJM4Wj1mlxWlJ/yT8sXc4vLmh+aHgXkwU87rAeGQ91KPpclV4Em3gs16
dTP7jn4mc5uUMSdR7oPi1U3B9dYC1IvNZ67LdUZV4s4Um92N7ujLSFc0ZFSZaa1s
mq14RfFTKGQKMfUaP4nFjbpkknsEZitcRCZv/vMCmi0bXkNR5vRiZs8+ZrgDnUtd
9r3KcFqZ0COZuLJHAiSEziaWCNobjybB3WBfnMjVStKwfYyL6eo5U+4wpz7pFeBw
jHmo2EFpphWQ7xuxu6DB8AWs5UlAOCIUrMaat887RYo5EW7HNRJbLl4yga4yOlIB
GrE5yDggjhh3PxPu95U5PgTOetyJQ5ut5aBXI8eicdF4AaO4gNSlBP0oi/H1R64s
tijrqZl+JddbeMxXHPK50ZhjB+IQ7dlhNt9l+kMTOgRHMI1oPmuWwySIqzhUPNSC
k/pdjEOoFDI8Hphm7aT0Mxfdx8TpUtgHzLmLOkiUu4PzoXI3HTT+MpiPbbdeqEW9
s8nPpb+9l6iwEPKV5BcrsRuCmuv6s9vAoitgt1N9a8xqZFq+LeYNbwayepxO/VHY
m1LbHBCP1ax+xmrfNcH/VSDUxunuU6tvwtv6N0ZAiTNO5RQ8aKRVCNtx2EpvBexO
MobUAvcX0zR0v1v12cUKodjNEIl/YuB0Ado+tncMc4GJRxux4nC+iqKIF3rIg9pU
AX7jPQHunSIAM+U9iZ3kF7+owdbmjGuGivOrvaMnD1ht5pI/BAPwucJa3UfI2TxF
Tysg299/V+VR2mQgZHH5BgAS2xZB9Ye0WctDseokT0jY0Sl3ZGmG8gr4ERxuOYzv
rFv7WcSghQBNeQRbw9WaQsxC/zEqJeikA9eUUsqks7cgUV8y5Xmcytn1FbCx8J+y
ewRGoPlt16VkwQ169vfCfLjj4DgJfpWqQYQfEJBKihaCE+/wh2g+kr3jCtVzX2zw
QqlVsQi9aGXTn2UpOA7rWV+UR9X1ILX7vZ9hVknKGdxYSkIshq7Od7abwx9fZnd5
tfkFSbcvY3fRu7elihbSHCGjunHsRez0+Nb4r47e/eb3C9kzlhv8sCv5v5hce0WJ
DMzIyZTiJiNF3TaSa1t1GkZPXxdBq6vygvZ/3CCgz8sd62clGNB//uup1qjTU4AT
9PKJUH0ESiOQxIEBdayg/3MDRg6DNRqpo7mntGrSQwMvwU8Olw5yqKOuS1UHqCXx
kQxhuoeCXduIU2LQlic2Zkgn5OrEjD+HO+rYiydPhKdJQSm60Anieqp9lQ6fUBac
xToc0j9JiYCmF/+Ie1svX9J7zlsAUBjghSQGYdwr/iAsO4vYjQ5lkUbngqhsfayv
uDTKMKuOiOTrwU3fDr7bTpuoL7D7X/O7wAbIc355tqX8T6m64DkHfdjxds7rhbYL
8g4/noJvpVrBI4dUfUUdCcfIlGR5Xh4wPNrhAAVWLMBO269/RJQF5d9jOAyvW+MA
QmTXDmBkoihezmSqeWmlJpmk9AjVSHwD9xeBIi2te9WJa6z83duvsoXsLuJbzvSF
wUvLH0TSs88/HJwsAvvBtlmAi2N6sXUAa26DMJyaeG7YVgdDbMiftgTtNLOfWs6M
7XJLP/ARS9qUaqkFAco7AQ4T8cL/DjOFUlmJhkFnQrFTvB7oGQu+EH7qMTVfrJC5
k44Ez4LzWUoR6WslQJhxypVejaIMt0/+02ztGPV+4tydg+emuoc/xbz7s3Xp7KZn
kkqcAnK+Y4RMB3nxCptzeESeEiHCohsleZ045t4vkThFxlW7jydBJmrx0iVo/DGm
r6J2NOL9Vc3b2RlAb+t0Es05OB7iaCexJTGAxV/PwVfgsW0QyyA1RjFomlrp5Uzp
HwbD7yacOYeWrOXUMksqH4jllVznWEXPLyEQ70h0nNH/mbrdOVPTjeaGI8WBC0uk
ABoson77sxaHMKNPnGqjVWVfiyQBrB3GVOyD8Wp3+pwDtC51o2OCgyrSqC+2t0c9
oVzdrh9S/T8Y9ghHT1nha/63+ifeqvBqi9ym1AurjMS8PzKqURT7eAZCG64Jrqld
fafLvK/DKKtcFwyK6Red5UMMQHJ5FWidQkmGdaH2PMXqGyvK7XCuMQIFVHJaRkpb
5BD+/+ixaRGT6SbCiYPvuSISTycSDXIF2WcqzOniyn8wmvvmiE6itCdeC4G7NsQv
5itrld761w0Bdk6Af+7geSbQgQjyty9hRfEwGMCNFiCyV/wi2l+ovVwDqSpvXIRL
sxWFgKjxcAIkhdQWGV+AlyRqEWqjlwFGQUYZHd/V7dZAwm5x+2JeJNP7NhdTMoD/
IDJkUOrCpVmDG1IxBKa8QQxnGpY53HTc7nF2+zySkDL5OmGd2ynV7RpjVR7EsNx/
jfP1RPRi8prlvUHk37e+Y7TcI0hfESSqJM3d1KOxcXzi8xBy1VADfKD12IaQdz6i
wYN2xxEd7eYqKsVoH3yQ+XpQCPJwVUqvXbVtNecuBB04Pj4u+NxRf2LfEq70sQcY
hSQy6oJxyY/ppcXge87jJ/dhN59mJxEHJGecNnYKoQNUYmXGHDGa5U7IHFeTCN6O
6pbWDwzDVdzMJ0cNSLrIZLUhbllMQHq2TTIvqAq+EeASzeQGffYMd1YwK/mqj7h5
Rgz5JI4csmhPPY4txnG6ioN54Wns8lTuiM9LIXTwIpZ1RE7lsxJ/PdUPiaE9o943
5bNOO72AcHmtlSrp4fu7wklocUtLtXpOQ5Y5yVVGzM6X8WGuSZ0lkgqkh0haojR8
L9D9/08hWV/sC0BPF/u26s1pDgE+GU5rPPsbGbrpChdDb7fzqZtSj0ArKs5uWRc6
7jy/XX7GgwRJp7dpVtN9+zEjemCgoqaUMKnvuh/L5Slu19d7nrdiDHpzAFbTp+cV
6AozM+vpQS413ED/kt1pFjSKCNHByiiTrMH9oAggXi5ZgqDVMxirq+mSkfbaXYr8
sTWWBX2c/vhTQ8YQQMinYZuDYjSTTuXjsCqicjiKnE0nGX1oJku3Prgbey6UX7tK
ujZuPp5tW83hQaLC1acjbMV37pvVAKTQr7S8/6j/yn4b2EuJYjEd7nWQWhuCFhMi
42PRpCfzAWdGNBeSs5//GCd+dzTKLrIpSvR7xap7WfDq84iVRhki0//TBxXYLKsi
lTljyQaStgaqVEE+n+YFt0I7yO+3r9QDYFCVXyLM+XWELP+KR3FoBwenYjcolQwm
+hOncw3j/uFfJYqtzqT6uCgGSglPbRvO6DNoZ2LNVVTS5MyST5QS7rDGHMjabhtx
TU6l7iyyHvanX2ezWH1A7KwwIlRs9hAKyzGEexseqd51q5bD0MrGUiozYw8LR7xX
GrN7WnZDiLIOADpvX+8B1Bqsg91lM6lonlmsWu8Rdcr8yQAlER4cnhZfIPJGW0Zt
kXHshMmYQ4kP3QmHIoqemYUBB9OuZPITdL7/06OrwafjGUFk+UNGq5v24EGJ9wCC
5a5tkHZ5Ry4QKN422Tc8+XAB34k13WtU1Q+RfOfrvQQrmlouukg9uD/y6U9nDSv4
Fb4B2e5/0UyrdGK8Xu0clo0IgA8F/acX9dTlLDf+5M2X6dXjJiG0a9ul2SK2KOE8
yfdVObQoa+M9DzZgfd9yL3lvHBdXL5b1NCb4u2Cc6blypQtZlRKR2jJ6eFQAGw70
u0u+xM4990+CJuB9TOYNqaepVo0ihMDMlFHl0B0IEWeeYi5+2JYcq+KHad/tgQi5
44qhmSA1Rrs5MMel4uIdn+hAiFtlZVtoTv+ydEGS7R9AArRqIJAkSDnTSpV2h5HA
mH7wT1drtjnNStDnPdjmxh4YkUewul+0/o1Refc8YEJxwY28DhZF6lxJOB7Hp2Bd
NzEK/E+b5qvclbckA/9e5Uv3P0XzfcNl/bXV+wGu79QSKKimE5F8lrhzJmpwxcNA
wOu0knKrtYwd3ZIEe5yZVLs0K421F4TYLlfg7UniBe/6E3r7I6ZY7UXJ+MN8AK6S
16RH7U+DHnGcXlYs/TBNvejTlg/Poo0P/Vswx01D8UTI5t9TAU//9KyG7J3i5I1N
d07rF27y76Mz+sm6V4sVILsmD2zPNJlmjXgampYaM2R+HgZ3XiwoWBb6JywW4gGZ
dHLek0jCmdd0ihhJOdN+YfNEzkdwax3PD4lf6Bu7s2lbBj6tfzEBtS27QsLpkLBR
BTDCIH9NADzauqZpRAG+1iqsx3mLDUWsc0qax4qeOF3kLgqv6jrvg63o0LMH3PNI
1NGfMIjwB4El9BVxJbKQN5fPoRu8AZAQzpR7Z12VXqEpAIs95di8YdXrgc0lzHjj
CoZmeoFbrUWDGxqZ/ShAtgm5p4s+KAc/86Qc9ip8odurokHnNu2rl+aAMu9TUSNY
vOX7vssgonmQmxoTb79cDrO+zclp+9VnqsZx/C4qFs1AAc3GQVBD5r6c9gxUXDei
Uo+UqjRID1ad+cNSYeifXuD8iXe8re7ADkrZV9UKTO+IHw30S3DyPRocUMhFuTic
vzGXw2r8YrV/HaD3QCjZKG2PYPO/L8H/ytRM5UhtE+/GPb+bnt5KGxWS4skFcH2N
kb4T6C4yWHkvyBCUXC6jmkza/xLcqdtxUqQ/aqbFVWdKE7a4GAp48nTsTK6W6247
jZDPfGcjTM81B7KMDoKQM774lKL3JDPgY4jkxfZRwK0d7i0ZL0/XEJicux5ZeqJm
MqQsxx7o3pNNRJSYyZVqS1l+KWkT9uf7vCGclKuRE0fYpdxIRKBzfNV9k5z/MlgK
Rkiq6VcjxaFpff1thuty6uYE58w9DNvlGHGuRSgWuERznG/xn9m0i5fZ6iX1BJSo
s7BU+Pxh/tnkI4kHFytZjg8WEe4x7ZcEvGkXB2Vw9zOqcFeAAmlBHy/0M0xsGfWf
O5y2X1ZbdHPGZyZ32djSrUcCywEQJghRneHCZAtG8VJqH+rbb39de5jy8F5EIZBx
pfb/pTu7jngmoo3qj8S5wcgcOOKd2EwarvGBmSlBE56I2at+MF676wQMgJZgryqI
VMdlTgOAKi/9GLO8Z4JGUPZt/B+O5gLA2oApK0z/MYUdhk4y4LcPb3UN+g8FFyDh
lbXtZb3Wl3uYWQeNPm4yiIagR+167KM6NY6LFE72P/r/tiKwWG/R5OGAt0JDXIsb
Rv37nmnoszGeK/YciOVs4armds4PYI6OdXYSqhGL7tdzheo8V3hpjWlq+OlwVvAd
Ka6gvNI2LWWPPVC8lvPPHP6lkE1CcyiANjku3Uzdt/FrHJEqy4BRr6dG94BwNvsj
r+XJUSjQIeC9G3XorarrIOtqvyMOhq3X5ihbqnXmaOZtOpgWYzbaHSVhtJcaWoTE
223niX0m3lsCd5EP+WW2vuy0eo7TZZ1pm3Wx59saDsj4hz8wHqZgy1P44Rmt6A3a
EzD+olj5ygBMrElkpp9fUTpBgDrn5KtwHAaUX6jhKzbWeasHbg+smY4HubKJgjij
FJZzmCCSlCR+0F2vggpQf4FUG7TpjE379v5TfLNhquWu8SPlExXkmEQ8glKzrQFg
llzcmhJSWiWbcG2YjOaZ5QKf/Be9XRrJOJaTlUy27vaEfKkIUH46i/kcltBsTT0/
Js4pxwmCZguUDtjMFPlN+WqrEpDSX51y96m+5nK5ctL5tSMuC1TwKiYYAtwZtF/B
9YdxZp7qv1Dr8h/t4qx3nUuGs3x6yi1Su6RCqso22D4XnD3jDLIubYwaddf7VPtf
oHUP1p7hcKc9re7ikx1XQTEhIhSKw4I2iIthFJiv7a8TgL2AaAtQluVOsQ8MalsK
9bA1MwiWO6IqKc0qmYBuU+7ESl8WIuhSZyvFhym9mQ9BPolhWbNH8YrbtO5+tvP5
RWfkvZk0WdjOKLYbUVb4YlPluzekL8PuSQpsmWCOfuGTJY32UBqRZI9APRnzA5jr
TEbsE36HACJoE3foH5wHOPTtNtdaz92uUE7KAt8jrgeCiOjXCSFGbn9paRS47qrt
R7c9/YZtESXi/CRTvASExAGs7aSwjL54NFM+LwRteyeiDAL0a1khwzUlFuKyjBbn
19J4yoJVarYFXtNG2GUIEiRm1AqCI+c47G8T93DVELCBqZawsTb2pGfQXESDh2yU
2Zu6ycxo82jIcxbVCN3sbSl3KGQOmZ5/mHgd0zpyCaWH0g3iwlkzeAU9jgY6e/xP
ubO0xQax5NBYqWElQB8IbUpV5HPvuWl9Q0oCTmgSggTX0EtDyLoEsUiqec0CxRa2
BA45ZUeenU98lEEhE5BgjAL2dCPfuO0REEaZz+DXDuDeQ3HL2pnO7GxSROO1FbO3
0YWUbJ/zh1TibaSlzCjC7ZTHeJEqAD/82pE47iWbTuNQ/iMsgiQmXL8jfn/c0v+c
wIF7dqZiUM7fp3yFjqu8Akt5OWdQJE0UgYAE2zCUziBQVKT9pgy+no55rk/OLvml
GH6ewZ22W8quEwn2E4wndCrCsDcek1jok59C1S0au/VOxQPWnOyOh9e5TEsEiI63
z3gK9sY+8tc2v0BngA6OTnctrgUGoKU2AeXnInK0NeJ07tWe9zykRjd4aw5GG6av
yGpoA/k3V1ZRrdBmebRe7mMspRclSHbpU1hOkRq3/6eBtwj8tHyGSGtykR0ILbhG
lbQmOThp6Lb24DChX3iiNL6oVAYkSAIwMudOSVl1TIxD1TmCdKcDXdiTR5HuaZrQ
5wExf8oefhOCErA7LJ/++KHKjfmRs8fH28wDA+WnmhZRz+YFvxVk3OviFl4sHJs4
PRBwIiOvzyl0x3hbXYDoqT6x+Ltmg/nwcYZy69xaos3GynGsTzqFm6ebOnKXlxsj
h8Kj4GznPNOiEaQwvQBmLD2zooKpdR9+1KutNB8oDSzXlu7EM08+4zAIp1CPKqwa
6nTCQFKux+wMSIbvn2OGNxe/shXPrirIRs4EOcDIlYvEVywU24nrdxQXGkWnS7il
srMAbHgmJwLlxaJZEUSkF4otk8m9WPWcJLgFDXHIkuhQ/g7hBRzmWWypin7cbSHI
1QA9voXzyVohuyaatjtZSjx3CJAuDpO/lUfeoTVHYDx4zlFSgRsCalE9/KwylBTH
Q+Plhz5GHcnBz+0NXIgFGKSHOOVaH4fSSFnj9w5jZo3rm0bzvyxAmAzSyifnSBf2
UoDRQYW2i6Q6JLJsAcvavvJbM2P3YaOn5RvDfQqvpqEce4eXmeFgcWFb/JyeDGDv
Stoi8nSr75/9yWf9/TltFEKvIZi8533XgMjPY3Kqza9oHmTl+/eVwPBOxCAosFvV
XY2VYhd0KttEf69mC32szuOl4XXpJZzQ7mov8KLjW1dInkxqccGhWkjVWJM9r3Um
0KyR0sYZnnd5+9Ii4M64nZZdg8ZIafIcFxDM6JxKqnnTHJdHQHBXKiu+5O/EL3ya
Hw7URZkKaE4S4hQ6DovAiqUz5NAq1B+EeUH/wPNkg+5Z2/tK3Hw1eMugXU2ObL70
HL+GI6sle+rh2Y7DJ2HfCSC2o5QvPOMahtQO1QrcUpRtv7umd/DqMZ31UAyaXZI7
c2XLUgLSurje1wPGpMwl3xZnNP3gKS4CgIfAT86ivrz9gOU+zy7uqAWren9TkJas
n36NpOHsk307ZH+sARYnUBzJj3pBhEuH9zGmtX86Bzo23PoeRgOhtE5a6JxIwrdC
qyR5oFp1I8sv7sovWxtzuUDnR0trnswJQM8fi+W2aRbKWUXRVk2CBJ4dy5G+a+ci
j/90SV/VIfjlxc7N9AjBQMl6uIZREi7dGDJAQDK9XVlrgHztd7xXq4VaJLTUXZXc
LkL4XD3ni7Xz2ya99eM1aOcUywSTi+CEXzTPkteci/hYDZgQvMiM2dXDPiBAe9FC
97qgYKnzYUwr7CUP1BRlwEYPPabub63JUVGKoMxKg4L9DpH55LZFJ7cpaDht9NkU
pYrnVQgzt1Z9im1FGFsXOP4roM+GX9rVaYNhpDcGU3huZDlnLBMn1u8+HNzvUe+Z
9IYeZtXoh/GPJ/PXCRjU23NvEDLW3vtVPEemod355kWTbKT87szQlFQyyDv2jTsr
WI9Jj/UocQM7v3lIBVH+1xGjZmZuXrE9+UmYIs5+m86JjAdHZb6Nkc4rXOJr/1bE
qXt7i6H3XYI33KJz+/ohaTEVQXrcJJKZ1r24vUqwwUrGmPX7Tkfp7DTyXYTncGqW
Gdu0Noym7HIqU+OD7KFsjqH2gzOF9y54x2CqWrmw2Wb9MNBzaPahAsz8nFnFKTYw
lBq1w8b0Ks1HsoaDz0ZPVksiZoMAG3SWEgubdI8SDHZPjie//UHFJKJC/AQtuN5D
rLvzT8kfjxrRyTODFXRxIAB/+jYgQ2XlcbSRxH8ItBb1yzmESp3AGzux1IbSCiNT
8n5INt7+wWUHmuw1bPO/iWXXCKL/i7dVKgvJ+6oB9p97H83zrxGB3QarbccBupZW
oCW8paYbKolrK8RnFp1HFJ1JLnkAM72LOM++wSbpJzgVVm/dgybj01u6y/OgH3mM
paajsm0bS02QYZIJYEZcLfgMrb7kF3wIpCXlnYj16oHbRoIPxhShoaLkAHAacAcC
uF0VZdoh1ludp//7iz0/HfjgQD4NlaOBqRK9peXjJxdMYT8qG9Xd/0XaycAemCXX
dhRVyArMiPO1jRFns/JEqLjOFbYretLO8xsSbmMFPmzaUCIlJB5R3GuNEc0MDF65
4PIZlo2T86yda/AM7i+O7edhVreu/79eSJqlP3OVfJSB48T4SNqDypLqGz1Hvi7m
sAvayOKb5DhrSc+tnoahXYCxMPYreF8C4U1d4Vie5RsdScEuSv2hl2zW1sOe3r24
FB0GxTVWxgkzJApGyVZ5c9Yt/90DiYEgXYzl467VSwHaL8ajOR1BWvV+chTc+LLm
qXBdBOeGbOGunNn8/gksRvCjmUIV/IFK7CwimwTYwlKwldS+Mbt6AfrqhcP/QSIp
WU4Hij+VrC2D/aG8+0Wsm9R1BiOWHKYaf3jaa5Rhjd+1bCd8e9MUG0/9x/9p6y4s
cyY50KFwmF2llWCaLDa0ueLOfgy9gMBEy4AHd5LCK/PaThQztfHXuNwld27f1aG1
mqkHPYWbIja2sQGyd+Noqd1fmD2h3R+IjfcAX/xVOhlHPwQgLjOYgLAxfGtRT3E2
6jksHKRQjh1OysDR8LLUt6icyq9mpVp28B4I0+RTJUz4Z3jloTttLJN0CcvJ0eI5
rMwUuyDfAsSjr4qeipLj7duVg1cTd81zh/DxmFmW2hhLxupiZsWs2Nf1blzSCPlI
hKyPc9M918rgHvmhbmQFyC9OWKEBLnzDzlI75nvF/hQmjPU4PZywYgkwpkJK66Ea
x5V2XPRXkMbOJn5eNTpZ424guqTBqyvxye/SnPvn+dY/sXe2Qh0wCgbT3sLclmyE
fYADGZlGiR5JuY4BvSm7Z+O3Qgaw+FBP8tyWMmzWt5pVkX+/DeogGcGTXURWh42o
kvBh4CW1/u46LGaKjt+qKgBydcn18iSL9hsn+fMKJ2iTpbd3y/6fLBJng7bd7Up9
KX3bLJ+Ie+omrCqmzIchooya5dqQhlFVC3uKxixLZa3fjoPNLBwyy6/+uEDZzM+p
EzPVj3jbFAA/WLODEuLqFpXUXz2rK1OW6eZpnPogHbX08dExqss3nTsdf44QWNOe
jw5DXHNJLgmOhwPva0YKoheCSTXmk7BpzDSV8WLyCpyOC8sf4VyY6jFOr+5ojpbR
Tr7rR4Sd2p8cBOazdYZHpl2Uk3Qe14fVNne89JMQdeaewQf5gBhNwkcp+I5BUt0o
HQV6T18hVJuy80TueONaEEoPpFFeg4Gx/46DOyz8gCqAIm659gqiIF9Lln1dvcjm
I7fR4mWXyxywn6Oy0Rnc4Fi/pAxXYHnf5G0qERaBvaLagKkppq6BypzYxy3vjHeR
gixtcqai9dEPUewQ5emWSt2a1C5hKVWevBywlcCn7Zw4MtQ2A3v+mNiuTKtBxGJh
UQnD33QmjmLgMgiWe3MuTDfSDJUtBHOGLgThXE5hc7Z9HWzKcIC8AixDmqh8daD6
oQOqqfvM2PTnTUCaJxBlu5sUXVy4J50YpSLp+AUg2s69lymCC/5SPVxvwiOLHf/8
69jj8gNA916aXNFsv2otphLJ5ckrwRq/jlHg9avc/zPzqlXb/caf9DH+gXSKRl6Z
YWJUdz9xuDweqEoDb881dt8yz3j1A2Aq3aljT4Qa64rrp9jE3Qo3w8xIxap7nd3u
g05lyMinDgWVz/ZuGPZSM79z/bC855fdLONQh3DkpFSwYdZ46ePT6cK0Gwf7C1nt
f+EH7twBCdpLvyi7TaJXm0AL9eHZQq59qBnOftRm04Azx/hEsH9IKWmMlDf5L6KD
M3BJ0NLahgGD2DVZ9Fm/tYt3LC3ERXxwEGRnr+QwCOyHrLxUNkCv8mQJbGEK+X2q
hLECZh53qaoudrgz42DX1G++/L3n80iyZDId/2nJ3+Ne+eJUuZ4TdfmjiU4BCEiH
mXOwg7oO4ZlhqibOY780SSV1wxc1ooxpjhoVb8uKClqg+K2y6IIxvmJdBqDWtQAr
dlOPaCElewfbM3bJ2Jf80BYiDCvVT2ufbk/brn43zrEzPp20qoyrKx1Qrm0pxMD3
b9APol1EK4NE68hsb7kBGd6eaDHIlSETTIm+QaLTip/dEfvRfmflHRlUt/sa6sRc
c1MSyzR1SRrUvIYG5fUnZUQtby9C+ma0CDXVc8SKp7J6V3BMpB8/GLn4aR+dXOW6
rUli2J0S/pldn67tKQ2oHtuG0EaycUkadAplxGyq9VaStB8lf2Fu0nOYLb2E5ea6
z1YnCuIxIzV0L3A7/sorzSS+oJP1APdNFAWaBQkxyaMY4AmbuMkPZ2auOCz0qA6k
NVs+KZuemlG0E/dXMC6gnbXne/zGIAGa9pJQJ0Z89Ptj4LnW4AlrVZaC/m7OlHRu
7QwMw1Id8YNjzOqbcdmhRlVML5gQ7TAS4CNlzYjaZRM9P5OMeM7dgpiaM2QfiJBe
dRbEHYvhqSNr7CNzxlW/RvkkPiRKBbd8d6p4ayfWFW4zKUpcomT7F3n1fXSUEQx3
9/hxE0VRuZ1C/3GGMGCNUEJgdqfARVD0oC0NDek9xGrgbp6+GtnkwJX4lBSJNXgx
ItM4tV+6PPm8Hrrdpf1EzNp8JqGmW71Jq6wmO6zDl2tZfj7P0Tzcbh9yD5nSGWXK
I41/wbv2kjFwt0hD2WlnCsFkVVJvrj6dlp/MibbuEEQ3uMRLNTFF5H8vvMaIyyhB
vbACfd+BRoHv4NjPp3kaPH8YwA9GN7kQdBbpvcVT7YBoV+wwdRs7DIpMkQNCJ51Y
1LfPbxq3S7pMkYNusxlEka8QGQigBcbHLWBdjdt1VIejLQlDMc3ZfcpL11DXItdz
pfzWzISQ59I0y9polZxRyIZJOQJ97EcvKwB1iOOH+7b02nN/NyqpmcPiyTnawxro
yF4zrBv9/f3ewUe+jtRJq5+2x5o0kAlTkFKp4Ee+jz8ZaTRox+EjoykmG1qmIhMY
p62PqbfE7nJh0973baTWk+NxMBkRWrSb7J/lxhi4uDN5yYR7slk91CI01EmXjDsw
jfq4vWDsyv3nKvv7qBSsub0j/ge8K6QOQe4t2RuunkCO+xXPaeZhAqzGz12QDcGN
Ng36wryaWq3XPxjvAQjSZrBoLdwIdPbabWxu4vfRnxFmFk15/8+b4YoGAwDDWjsr
VHLPXmdR3sMdIUo/fFcng4rwtsKHvpXR7Qw4Jjru5utySR6Ua/2ZgS4UgJavA2VR
a7pz0oyP+LyB5GCEfOtlzdRoM+/z/HICfJvlwMHUIOsu5GzwqNoB8rFvOvxaNlSn
yi9DxmtDc6WFI1ee9lATI9C1ULXkK50AC1xOf+zF2a3cVYdqZ+YkTsj6iwj73aRr
cwAMbKARXsxgzljuW9TJarkovT1xSif6CLxaqsngY2JrYnNys8Znx+BjifLwyoCX
Aom849WFeIybYKtXV56xcprS8COR4KYtHWLS5eOL+Tf7FN9pNEQAKF8R09yFSzYG
Jy9BeyQ0wcF6G4aH498PiYADtgpPKuK9U1oi3K6sxSYN5WmOPkysm9Xspdm/zIXH
+HM2pyQDY+F71weqEh418LlU1sxmGTJ0AYnqz+iK/h0kt7lx3gK3lhFshrnWEL+B
119KBmzAnSlN7hpn0Vi3kGAg55I5L2H4n6ZiuGKOFS+HPO7mTn/71aFTWp7LxmXx
wfnnh16oMfbOLN7nQFXTsrKrBtS3qis27cNxvhgG4OiKHElG6IlDCWeg3Nn8B/Ua
4xEvvQS8U+ZTfo9u6Z41+MnAXtpiSFeIRVyn6rJM0mVxYljztCx4MwVI42/fDSbS
2sollmDYWqfQzrxktuhRtvEPLiOEWTokntS8MaUGHZMMHDSK+SRk53eQoY8bgJh6
weZX2IlX1Mxc+35xZeAWnHhd07oXc923VVN9fu0R6ijZ5QwxhBXUqTN8wdI87idf
i5vCTgLgtrpOOw0DqTw+swbww5ixSTNanpq01WcPlrquu0hm2NRXfgfOTBeV4QQ9
x9h9w7emdqvMyEXHWaWtg+s3z7B2/2RHQhgDoS0l3drAnGh/nDlCfd+RNho30aSV
RChVxErNY7jtiqngTbEWV39EYwA7xYjWKDRDwU4gIj66slpO4RIyTEnXJ+m+F01G
c5KZtfc2FAriv6+vY8fv5kPFF/nHGbL6UXY7mjXl7WFbIRkWNTDkfy2K/t47GPj0
Vt6KxcNwCkvo4WWAaHZ22Br3WGDn3DjHV2a7ENZifqwnW6c3IGZjhUgaZlt/N8oX
9+igmCM3MHlu3nTmPDk/EfSdTDEHguAY87DZgRCyEG20otEHix77OSLN4a/+pwLp
1gK27VRdi22BEvGLEGFnxI6cwtF1GpcWnmTRisyjIu9Gkp2I29XPzZsl9R7xOvyl
aa8grZtx2vEsAbyU9coY3iL3LjoTCdNk2WHx4teMq501JZy9mujc+EY5t5+YMyX8
gF7L+Fsh48PG7Xnuw6MiQZuiBX7yRninNPkXmLHo6gB8Q2LM1leWjGVZxKIUX3XU
1FX8/DXnF29BCSxoDS6dXIN7SV1giWB4AI2kQSGJpqUDoP4knqJiiudRD4w3cfJS
8UfjcCSriUVVTwjSp+E8d0opBCE+DzgpRq9DEwgGzcQG8WgKBV+qGzlUdNOxELd8
MqaAOEWcZ28Hbvo7EsYrmXS6ZpFnqEiB+mR8ISXJZ73pJTHrOMtPsg2NLXdr3YYr
8oOHqYmDHNh5llt4QlED8F/k8IIifiB+8Wlp9PaVKkf3JBrPl2JJhOwAZcd2LCN9
Q/df5TeeGXrIPJE4EoycNehRWf2YoDxQipRAtFFvDuUEGXTmSsMonpjMBdxytQ1k
B76HS2v7hUPzzODPGppnE09hwtIrijZVA8vy45tadLLN7uNQbmN0LiXxfg6EpMca
qV8IcPypAA1FtrIBnqOKt3AZ80DPM7lvULqXqK9bw7//BYveXAU8siOs0301tZLU
47cBo6vkOvHGRi0g1I3YYDrpy2ZCCEb2JZAdLtkb5yDaLvEe1ewJmre2NfoLO0yn
N0OVBTMlCgqji/q9yJTtGx0lsFa/AhPFlJxu6EIGSr7AgB4vFJdWhxTpsWx4jS2z
6FNx6QcxREBDfUBIVjPuFG+zW4fZi1wFc5iyB3ysvDTbs3iMwPBpcupRXnOIS+AR
tUOQ0t3QohhUaxeqXaTi0N7GI5MoAxBQD30PS0saIiebkk6Pl4G5X6iwV1mdSL+j
zAWk0HhVQcLGA2IV17YaktlLPGIDKW9AOkRC3gtCGRL7Q3GqNHTZPuittnfKqyEI
K9Un4YwYCof73J/bLT2vOoeOnQTluc6tf40KhuReOMvf0CZORPww4zEdl1Gt5PdR
CwIpEpeCdMOSCXNJ0i8BU9h9fCbrz8fSz0T+5yuBkRL6bMFuMEzXVq79b7gq2EXH
DJPXzCBXxGEkUjibF9midHedUSJvASSSRdoTlRNlikyCcMW6NCw0jJyUdj2MRvZW
KgVluJdtUXw3Vy0wO6zXWgBpDIZK0P7aJZkqiRxcnduN8gTnE4wOBjP9vXO7CAQN
hd9ynPkQjkqALSQvmnlokKJ5c/3nM/xZDTdTlLxZdPIm4XwqKWDaJ70yKriY6B++
p7Cdy38JnEY4FIW5vH0hLN1gj2TUtm6OI6/Qs660/mV4+sEbImmGtVcF+rDILdG5
n/YeVVKS1j2Pqn7dA7Dvt2RiczMgVlwabA2LAZEP4bTY81zCuKc5b0tucRqyNj0h
xwFXI6P934yzsnzROgrG4mxwzeB0VOdQCmDPH7tyO+bSA6bPegcsZ69PAfKHckSD
4Taj5qE+pJzbIS4L3x1ZsHS+pLSy8KtIITWiB8/L9w0pwrNcCSFsWVoVCV/M6qB1
Av3LFyaOmiv95RGmnuXka3kett9vCdjK+ss433raRrnOoLg2aSvsLrjjp8j43w0K
kNV4oxI8SSqPy0jdwsd5DmbnauaI5Rr+3cJ2eaJXbzcLFT/QB55xVg9JaeehSEkn
d4PO2Ek1ViqP9EU0wpqo59/B+3ti5xMWVHmfeZcYKBmbZIN/Oz+C2gS8nzQomxsZ
qMlAhIE+MGT9ldL1cN+7OYnFab89C59Ae2qjZE/VWcpEc9Coe9bN4gL+0pX9fBek
WbWVIyozi1S8eyXaUmCktKwyPoisKG+dm0/7KFD2O3xIFcWpCeE0VIbtTZIDJ1es
la0Yc1DZBzi966wfcIBsq5TeeFGDsCJSPUewvrSBgFEf5dg7gbzaFkgTLWubzegd
i0Tc90gOF4zXa9sUHzI5nlUfkIa62W5PyIEfFObrweuilztZlwxzHCSYQFhv335y
8fndOmsND30SyUCEPCLo9iKngPp0I39W0ENDV6b707es49m+Lm1LTNB0SWTgdDxK
eUJ58i0vYulu3P05dnvBENwveSlUNwtFgriaPYYciFcrN8BTDMc1yTEJMcsYJ00q
zYIWNq7uQCOBOtUt78vpJmPsr0AfMQpKS+fLE11osMOqFr412be6FKC1uvnrcpgV
LfF74s66nfmxek+w7aDIbBHJ/dWauGTfyRHxXi6Pa9/QE/i42K7/uxPn3b8VK/Er
0ZZFyY+1oaUu1M9t7OJ4OcNwhEWQfMJqqcedTMH0a6tHOok3fh1QnqaF3r48lFUW
IeY63yHj1Xa0kJz/vLJ/bGODuoaUiA9nWEf++3ehmEyBfeG6saogl7y70dPYf3s0
7h+WTCUdzvWX+cdy9CM1I/gpzX6HpmZ0WZnj5zqlFJlNtASrrrjbwFnEF4a12YWo
B4qU5wFQwLW48HSNvM0ViooN02CdnIj0y3uacnz/mgpEUK7K51VvF97eOrgAllYF
qWVUwugNpoizNfpYsOHyy9D3N338Gt7uD82NIc0tKY8K6QvVt022m8/P9ENH0aye
hbjZeACmqosZGF+GofILQe4tiQkya4CdI6XVjv3CDmZym6tVICgB/g9rfq7ofHxV
QSPuUZYqyk5PsVXudAC7A1n9uoI0fHnteOGsoOky55kt0uPMIhFy/Qa1K/cJs7fU
/QPZiFEdoNpfEFdtDFzvMsLqyPoSC5FyH6eS5A532FpEWk7RggjxrrT4FtPdkCIR
IQ1zXem5DWXSwQVCr+Gh8+Y/xzAc1oOuK8+KmdPobJ2QeIdRA081hTnz45GrZHUh
KuL0UHT7+743OEI/IXSZRk8HNReADBN7BSFk0QOstbTEpUp1nta0UtD7QBNWziHH
qmsSCBpo9Rl+sXy8GVzEe/zIIA/qH8MHyJE2qDWccPzc/Nh062/SR4YoC9xO/1k1
flk8GMxoTycqeSK/q63PiAgzy3KPVmNhegzv/PFmjYsDPWHIOmeC0kI7g3w9jlas
zHTIXX4Vo44XDizfHSt5IZp0s26exRvLxnqum2/LhBJ1c2owaa+ORKuLokluyim1
DU5NzPwanVuJWenJScVIFspm+nJ3lZOHFPFh3hyvdibhIp/dpbkmd3ElxArTJz+a
5WKb4JbjjKgyurMH0SRIqOYicT1cZmHBV0yewAcqeClla7MFP1eB8ZIz+DSdjsrl
uQ3QL+h3TSNGkxXq/gatJfrbCZvasdQU296VitO7AChSUhfgYKHr7gb+ILcc/8Df
OLs95LCa7YdWBafh7LeeL+w0UIUkROonpeB+4O0/NTcKm6MwsY0AJiA2uo4oQohx
x6GFsEfMll1J4fdy6/Jx0pER+joX4Y0WyGc/vRZPPmG6QZxS3b0pajWsJ2jmZT9B
7bWn3XROhhvbDbM7gjI8Nndd0DtDrtsaF/QwDAyQqndhvF2XieounMNd2axu7v8B
HThD/faSKYsBLHrWr1cc//l6NFyRIhzxcfTA9XDtmdidAZyHvqoSAUJv2G4KOY6M
JhrZtB7oad08+Qj70M+21LIKBZHJgDw6N8by7B2uZeNMQ5C8wH1MYYAKzA2Nbja3
/s86mSoySzptRCEjbgXJFTg11HkT3wejQkObv9n9XCp2bZiq7A7za5M6m3/AyLs9
5QE/NrQjreA3QR6uxHkwdylOrr5/T0XFpU3ibn3zPTEJy8TD35D+2iXuM3PuIN4C
/1ANXFx2y/zt3PWjv9t8bIc7kMLRXJgqcc2HaApGRmFDymxTjR6tVoPK8GpFMoGb
fVjBCocdhkZnmYOFrTwV2uuc2og8Dj5NnioJIJQhuRtAsfKIoVYQJQNMrdrZ/T5+
dLC5BcXi9+f4xz/SzZIpXGEyKXSe7habXaPm3/329mcveGZLZhPYsQ9wmEEQ9UdA
dggsKEaIBtgQSC4TdiDDzE0l5eZf/kn5mcvtsI7/RY9wf+QphZMNOJU8EczV6K0P
Xs4hfGWzxk3a+cG8lCJxVuGKMqAuIiLF+IHli9qyl49hy4bK3kWIgfNMa0dVK2f2
NaQpmPH1WQxApcIcV7pLcH7Y5FkcTLh+/grmnx/e4VKqPAA0mZfEpR5IqGFVtE0/
uzyFoej85GeN8v91zRW0ahtvT1tdBwE9CB1lHSTD/RxW2ztywKArHPfXOa52FVzo
FFSEAsK3wpyaban5nXbfXxSE2zYPwQsSi6s8Cej9Y1OSedQkp5m/hIeOf4qlMSr4
4IeFVL5ecCWvd7Gr9AuiegSDJVLa0ufDU2mBJtscaIbJq/PwmJsxaJ7HcfTMjBHO
vYl77umk7TxNsKuGKcypUrqOZfWevdEzEkrPZa7RFR/jbvPT3pxJWwmgXa7OYf3E
VP6dWqMBDyv4wOiDxmKYSHo+nvHJlbKvgFr+EkVxARIFy6E5t0BNpGIZW8+EFpdE
m3BxDG6xwjwza4h4ur+X7oZQ2TtqLk5UDwSltXbmH5hsDqpRUlsJPtTpXDuwYc3V
2lfvWwjFhD7yH3XGJYU0m4zwStXlRChDkAum86SQvHMVvLaWKzD5JBvyEiT3aQZP
VGH0H5sszwGcYVWSowXTE3S3LZNc2z7wN0kxPOrU/ayT/OTviPq4oCJg9Gll8gEh
TADsDI2z4KdYGvpVrKoIaugdO1hrOpEuG0YllfSlj+PeYSepxEKTHuCAV7lP7EzH
aH21swrOQKfx7pZ4hqMnz1Ipv2hfREaOie+IguoFHr7W5T0b8VZdDMsSH4iPEa6r
kDs1xbInQ6CjapqkIwnEAVVyq6TMfQS/2ssBZkiuifHynQZ3/iRwUYNkgJ3o19E6
D1qUM/L2QAvlKkNWgurZGd4eCaBfaL8NxamzlUQ6ODpd8bLeCfRdh3/u6+VKcjil
WRjBdOXJAs3P6x8mSfw5ts8GL40QnoG5Ux6xrV9lC0gt8+oPvuSyP47zXJdu9iqN
ScDTTmacMWzKF5zpkVdWCp29L3Em/NLGoB1AnYtLYeiXnz//NS59GVX5jLg5mOf5
n+tX8mOt3rYbrTvC89oXJRs5/j8eKZOnmXhRhP8zQzDanCDDvDndhRcoo/vuTx0N
cINMyKa332rgPXNCQj7XRsR49nM1R1h35rj2tG49IkTgnLtK8GgyjTvDb9Aa/DNN
Me5+/42khRWnI/ij1tf786XLS+VsCoSCtlSqkul0BeUdkgzsvaxsAlwAoH2FBMEA
8uwSFqkZNkmkNDFzjqRdwkVlSOaLBpl1Rr87/7/OwsTIcWAzs5oEqHk0Sw1pJQwV
DwsdN95KSCuE3FguZHdrCYY6uZtOstNPneR3IMH7E1zCh+1lnUAl4fcsT95ERxhL
6M2oFZpcqA7bm1vFNzTBzC6rHRjuna1zn+FK3oUFVfYUxXefyviId5kyuRZYDuWo
PY5129ZuJEDhgOD2A+nWWTcMwFnBFFui+8J9bCkluiCW3fykjMdMQzoxtXvLuEvZ
cC68pp2hmBi9SYIDlSEBlNc48c6sy0gHIi+CW9RTOW93HfORSpZzhZyf/F/nCDnt
URTbToLGiMJhKgDEZritBp1wCeOdM25S9PEApGt64Tj22zdTmGKjfUGilyA76U61
XFU2DMQMuwt+AYHWGgm4vnl5iaymd+NjkQjP6ekoPRXq0MGs5XDOGcXxm246JEQ2
+wF4x9xrGtPsK/CgiL6mCx83vOa4WWsjrmhSgLJyCONo64LzN+EsdMhSXjKKAMKl
NP00RQ/wwIqKsUfxZQxfYzmGRCkoiq4tf6LQgW9Rkyx1mwA/gsJ8644+Bo0KqyNX
w9/aYW6z+PZmIsbtwRgoNslct1xyD5PVpYZZzfynx3/wKgNX0l/oX0PpfeEQh9RZ
LGNz38gNWvaROK4Ru4aHERzCrXt2DQpF9BAaDJwLmg+mojL25Pi+h34G8RK0U2/N
GUfBaR5ghj6l6dVSDm/fuUGsx7JHjcRvfTy3dkcCx1k8zfMZsr0qJKW3C8/yB6kQ
7eywPAPA2RoO73HQSkxn/1gFUkvhpQbQmGvVErx7zaSHSZ1/AplOwG3w1dtjOfB+
GgzwnSR7wBhSEXINTZ9uqBoaYUG+ErqDLDmJZlwJiGDCeW8aiMf7C+A6m/wFxBiy
s3jMSTdZ9jtYk1VUTpxQ0w3HLE39h9js2OkHpGPJ+/A0Tki9oYGpux1g2zGJMEJh
WTURnm9g9RsK8l7ks5DAX9RfXGSkDfGm7ItpeYOc3jYnquhuaSBMXGjyHJlhM/+1
W5VJvF/7fAoZ7OlnLTj0PrJd4VDO02KFNMJyhkXOBGKa2qa6Po4yeIpGmPXrz7bd
Xw8SZZ7RfPrUFxrNdrBfgck5uL3SF5Klf6xIQP5QzmtTY1tQ9DFWDpBX1I/qrfe8
StJ4JN5w9p2544BBPfXITRCc4SmXhgiwgJR1zUZZ6JFu9wvKtiukm9a3EXFntkkC
0sLiWNAC32CWZxTmK0YuB/Os5FyemcV21EMFwn1B1XgF2C2e+mViV8EibFJmaqUq
8nLHgol+lE+EKR7aRoGr/Xs/mETxl5nStA45f1mcbKoDaV8uBjf9RVGobzTruSfg
ROJhMxdnnCOOa2xiid//jwT3NH7e/k0VHFvT82dwV8QeSGbT6ldGOKzqUMH5GTrA
rRYHQxx1plHL2e517rM7MBjW1GGcapy8R1hxDfG+GqRnlYn9x1385GYelf1smmJD
U4mFK498TbUQhv/TE3PDW6V2JKHAftbSIF9PyU4k24y2K7DI+JRFro8CN0DSMJdR
s6OFpLvr8rua0Mg50B12QRE1QNgqEYEhgC7fL/HHd5drlCTaOaQSC7VltJdxdS/I
iPH6CazBVYSlT4O+g93bxzhz6NkiwxJxrXMT0XmSzUY7kSsHmEkkIahGaZFKuFxO
iV2o/ZA9updVVnLp3gEZzVN29gkE4RlpQXWEVSJYNKvfBeSImuOxSR/3UVSlMbUS
mh+6n7hv8lN3VIUcBQTmodQyeaxQxkfI4+WDX+g0/9Q5BccIsRzHRU1uuSRp+0gB
8clHsH6XSNqy/Syd0XIjQjbceRPC4S6q62tWT9DHpwwdF43yYFvq8k9394txjYTP
LNgqsrSa3x3T5Bvt1AVfBsBd6I9Nu8WOJuKz8+ltLbzkTuJbma0X+fmSXJjXZkeh
qCti1Yltz6TYlVZ+1HroLbriTz6Q0q/P9G4hp7edbpCxxu/PEHo1Kz/BGJvs7LNv
L+dCpJbP+sF2EGtHY0tTc9XUekeSPD/TkWsH502Av7V+EJscDXM1mJre0+cOimus
WoCMzygN3UCIRnAzidHxGln7nIpyyl8/aYGKbdhj6xDw7dMRUbGd6FknU1V9atwb
5MkdhJvCdlsm7g9Tim4ePzQcWOlSViQEOQ7ppt1HeFfhxRIRu6QmDDdKJlSsHcSX
xeTF+NBklnPRZsBcfhOg9f3RhfMwyXaZHWnJ4ul0z/wxOuJqnKDsJx+6tJB3x1vk
Ne1eCFPksCcxehcRPaRCM8DdZXMaqWXowIFlna5ukBbVVsa9e6g36ACM/sLCIqR+
16WjRSnd4k7JLQonVHbHG0LQllBgMAg4uNRyEzY3TH+qXZvA2zDBguMYioAufdz3
JSAWaarkKQoRg0wlNmRUgN9bDQQMZT75+glt8qV/oRZ8LILNKUZqlTDa2KTWkMwf
AksLgIq5FPTmIw4KN89NUf1aAJunzv0nNwvwMCDJ5eX/4ubRaqIiUae6x+UFzm7K
QDWIkj8Ye/gYOJfjjKum0zpP5vjCrhD1eb+lY8EmuwHJstOuv21OGCiqMEKZhSJr
EdazQ2d0/JFV9tsSk7PRfY4Lx/4sx2bDBAvoBlOP0Ahlpg9KJsIchCd2PE1p9TSi
+EL7qovRih0YaVBEGim6g6moy+zw7Xz2soneOmQjuadVU4z2boaLREWOegq90uzF
KXs32UrmvxWu8lwDA2LEuTCwXyqC/T8HloC3UkGMtFixZUEHwq2uEMYPJtMw6sOf
BTKk8hxX5dYYkP7hxah+hJhagw0WSlFyWFFnspz1TabQ7KuLWtmGj3M11lIK1Xnd
tUXz8teIdSkMQh4vXLyJRo5uYaFHVioqbb6jyPt6luj3HVsaQujm8gnkt7aEHRCs
jVtnPwOj9NRUbACxoVy/SOd6jD11gUH6877lnbvnLIqvwadrB6gdBFHhTBw5a4vk
DF3E0dTSdpK19miCyRr1V6rAgP0xyFm7wrSbFy5WtoBEyefLue7p2KGYbH7OB9fN
1B+CclafKxpkXHT694yDlK6jYGGoob5RthRAz5gj9nrjQuaEAVFEqMTPnh5hr2OW
zz1iTmKdl3lw8kNO54tnId6sMSgi5BZw4BInoOFygGMSGgKIPcBISq/A7dm2PpvI
PKpE8bbE6fkV6HphiTlro8XQKajGE8/fMTL1bzARImk01BlZhlzCPYFKLCpPLUlz
+nATZbJfNEUrZ88iqFo052X4mFss+jr5BH6KQr83JQ7Yq1RmnZHKM98XK556VtvG
PfJqZ7LLfYwO6mkfV1s5WD/bIaZVqXrPROgsbVBBLrcHpBGdkpGOWvBYcN3aSRf1
u8tARZDTvmZGsm2CPORiEDCxlBR1VhANmqHeZ9dCM0oboM71N69zyB5WAoBm2SoI
cx6nh1ajF0XbHGFvvuY791UHZKEMfk0pkvoRAEarpbFQW0DHpRVNRsJ+AkekcU3u
s3kkNcvQEREP9WN8BXRebBP4Ep4cyyLhIhF5D2Uc/nZj4bM7mDb317h7tqNNFTbo
ch3hVDhJf4Ayj46EvVaOi23YkjX14ZFCZgL+fYepqZYImSS+9cCRwV3kgZb5ce9o
cAvU0hdeQIR3wSb0P62zIWWKx+KB2jOxqaC2WyVrmvyH5EoH9OW9igy3nMamrbbs
F32SW5MikFG3W0aRNA45clZn1vX3JdKWQhVx4eSizXT6VPbF/oJuFVYwnvdZdfic
yBRgzGY4H+fAPxPCie2uWFY++OUiq75lTf568aTu/C2m+1R89yIlPMorea3c7jE0
7lrGteWEynQ7EKf2Esu4/q7hNLbc2469lmuIjA8uGLmIxhbNy25wDnTbIBwkJX9Z
+HnQg2pheL8NqlcDhzoJsL/2mVVlx2HxQSnPX4S9YBrFW5rlyxnMwqz8ZR8CLMBF
wPQ0uTUKR6Sv+LUpd6mbR8GB2oATo4iDBQwN+9BhqRuWeOdfK9b+0I08weNbGB/A
WiBoXDA82Ow70bgG5ss5Oj8j1OYU8nz3STZcOp2Hhr3hE38Z2mfVAIzwtS2BwgXN
P6o8v7wDzJU1XnKoyVgjvaBYXHVJWGedH5c3yVmou0ma/B4J+vxBrWor+MrG8QpC
TX908SeugIIg+vevzf0Bqm3KqzUEisTplOChoUVo13T07PZKc4CQSyKHiqPFJ9kd
5wxldE1WAxRucsG7YoeHkWJMXV/8d+so0UQ8kT2+mxWG3RNLH5o9hCsfuLmg64Qg
M5xME3v5XtDGBF22g/5WF15UnSR2oTRQF0sIoNTrYvwoicErPwUIytQ+DcF//SYe
Mc/CGta6zkrSxDyjG3urJnrM5GA6qjKi/REOE3FTjxGxEglvhjizSDc24OtdGiQr
joY+CWl+oOuwyv4YlHqXf1vXRWfZaE8iK4AyiRd4kSFQpSCAhwS65w9ZCijnooT3
c2RSacghMF1Yq38CEOEinNNULr5xUVHJVbiZJvMoH5/XPd2t7I/4XxRZJqlI1KzW
dBpm57V48pEl/Y4MvhU0i/q93Uk5dgMb+XZIFxElSNJ9wQSYmls0f/ltGArFTHk8
NzBRr8x7uB6AVZWbYPJvXFtIQRRNGM0GvTTTeDx/lypDW35oOfG/Jr9Qngl1jrhZ
OJnG8Vcsf8Hp0NmzTe2qvFBLIZGbiCquc+RNSnRA1hpr+de3XOZoudjyhYK3/QMe
wP9H4v0ouMZXhTsLo8ecAa8q7TxXpUYe1zm9tbb86IuT8V8OKlzo/YDPO9bnDB9V
hq11TxHeJ8tmi5JqF63qXmQxcuBLF9tyR67SjYGi0s03KLb/uxV0jwpDdedo25y5
gcy1oS+7od3RNWQKkUIyMwCuD5nDPcThxPzF68m7le0hOVlYoLIStYT3DTCuCz8x
wVyqQZJ/oQ8mV8Dhjujs62H2GfuOCVSdJtuxutYkCdUR2ug1rOlu0iN7cfhIpf6A
lrKTGAKJ/DBs5JLaVzFnWNQVeXVHMT30FvHSczHfst0ObD1hoRY1IZA/fYtvV6jl
4e96nLW+KlRgZFdsCU5niMdaGO90hvHi9oOorbAOyyGqiJzMLRwPFYEc06fLIeT/
wlVTTPswdYjyY78b10fu2iBl3oEatr49O33fdRlq7eXFAd7AFPrKJ3GlG2yz0lLQ
F8EQf21tzCEhiqtEhNyhYcc2547dZ8wmfv2JELjAg2QE9N7bIDtKnNpokmBwRut9
O+kxMFQMEaE5X5x/wOpSqCbDFnTFT37iW5UhgIpezBzPuUAq5864k0F6fDWhsOcx
1a9lp/FmwmfTrJ+2ji0YDFs7i8z7EJgCRS83RhaM/UL5BgX2E49YNp/hgimFXb/h
tqnNgfAtpqtAYtXXYD1F02QkTjTMAbKfmXnK0958G22263wwNVVdlkLR1/5QQjos
MqcInhoyp4geG9CPWpmgaOmCBOWmLCmJTi614CXO8+2tyKJ9EP3Zs9+yRC+WwiaM
1YDXXSSAlKJONCkhPw+Jwigp9E7Vpe9oEFY7MBQtcxe+9BlVJGivFETtkFPNLe74
SOR6AQkZikh7Qu8pw5lk6T5yzFSv6PzREL9ySHKOO8DgACv7/x72XSQRYNS7HGTz
WGhXkbXdVWCVqQ2Qdd3xMSEaIXy68rns+Y7dJORMWrrq0UN9dk3GUItsM/uHrPXX
mi2gJ6z0rV1KmggBKrIxsKyB2xU9ElLovx0g44LSni/vqONRP7xKKwondV4zva2f
RzfpX+OuqWC4PNzI2zoytLr0ULWJX0rK4EHGo1z2TP654L8uw/skEpt+U5/ht9ZY
IMo93//a2l5rosQLIw8fdAHaZwq6Asn1Knol3pua8gnCY5OZujWaZ58tMweyM1lE
aQi/lcD+HrjcW2pzq77L9xAH7rfPWTfvDcRWXrxVjMWG3kqpb+eqsAeqD1S2dNQb
2/zADtjay8ZFr7+XnfvQY/Zq3Rjt5fkiKBXBlaWg3WDASJQaK53R9yrpcGVzjavI
LaaEdjfovwiAy0f2tFkh7mZLKfHo5DLXoc6pD1vkCPNkE0S0VSiW9KkOYL9MPPiY
lx5YOOJgZZrmr4OoonhpGJBCOtjCYgzdCJGt/sFd1rW4Vqfj211Ivc44e42Q5Ssr
//z+KCIYxliEyKvQsm6So4OluUTH7yhatP01eXpzfQng306jZoeiMuZ5w8b6aSZs
cUPg6rjdIUV5Y8DbDdHKWMkJ5vygkXUljBPrbrA+KPOqvpX54NwARm+RVu5w23+J
GVUvY5MjgAYDzkdKCArhtfWMMpo2tylHgAHhfyWpwNKro9N5owkrVjkq/PAHD7r0
JiYLBSnMb269ogC+h5KQxPh9x5YnELYKiD+8NczU+9uo1ZoX7CbIXGfMdVyzydG0
IdiihU1ruCitgnY3OsRXwXncXA+Dh5cxrLZqhUe6Ih0unj2eqliIzWInvvK3npL/
QT9+rYy4M1jqzlMh3q1CCPNSPilScZGpjPlvvH6fYF6vRYP4V3/f/oh7anonE1fk
AimokLpZaaEKItuSRoBru3a5A1TbpMw+fAQedZWaMrYXFuXy5MKa68PJI9NQrB9l
QZrQiZMVQq+3X6rVoRKJjBMukztSM+88Pn2lmZgz8Tjh682C3DjgIxu7Fn8pnnTH
c3jKZExo+WaEI00fxfAKrHq+dDwc6BpCPYjGHAwwQ554qRNe7/HaWFc7Fexb/Vsi
1SGzXV32EVzacP7AbxpeEEDjL9cmpcL1GkyiJnjAf6dvYiqtfyA6bZnCpw1auHBo
HR1leWrMOFozpFaNMVhg1peDlib/T7RYSQN14t9MWttiBdKbwI+ZPePUN1/gvSAZ
rbcgrDyS2ns+S1S0h9quHRZzVRjDs/qhoA5mHlRuH6PCdwMZ/4d8fdB579n55J2T
62El2CrJedqTf1MyXidCvmqDDdSDIlHEGvpj8Pv5Qbam0VB1MSyCQvdn18Lxe/ff
dtyd6FUb14W4AzhRiBHROfbahUIv0jR0hh6/eoWwAq+Fq0KDz1LJrYuWIgc6EeCT
GH2PlGNyytb7SeQB7aVGmHBlMSlwa0shG/mBTUe9aPVlcDpbwyqvwuciOB8LijZa
uyxRgHMntp2m1Aa8XFCiNE3Zwp0BQciWoOKfQA+arPmGF3lPHCHJOkfMdxZ5yzmY
avAnIH+MvkfOWsYGBCARZjkB5TTpvg4gUx7o900DMQv+yZG2SPckKbehg+kq9JSy
1amVqkIDedDqSPuYo+cXckIliURtZVoCxvcWcxNs90ht/4XSgcWE3vRUaPJaEQ9B
rNyXK2fgHIBJ7GKr1TtdW5QIsoxUBb2k74vQav0yo8F1U8LKUFn3gnemf1HErjPt
NPgYgu1xIgYCiXTiZrJ9cMZ0HcvfdnYZRt6P+t6WbI6VK9ZChtzN3dcmAPwPDZOw
DQHeLaQ0RfkPBP/jYQ5pri5UFtZd601qo5vM628YhhOuvU9rJrD2Z/Gewi+8lrD9
tkdwN87/zcbbNIp4AyYIgdPwVhlZtTfnrkez38rhv9EjhaUMPfLHzGreTqBcQ68b
Ko4wESWDiAotJSH2+IFpgZPVRezcQylyd8cU6/FlcKGSzzL6kgZzXRu7TChXue6U
v/tyePe3Cu5A7R+bzj02fgd5cSunBZ4foHKTr7GM53nw7ojTlpTslkRhQB9WP4AF
QzShcBpdx/12HQnT2ghtda2kzQe67mOKycH1AAyYj+x8BmJvZNHMNW8FKh45Pz+k
5di16O+jtI7vKgDZ5ETKLJSwtzzsUVp6RFFp+O0ymA51sOx9Pakh+KCiPxdzSlZB
vc2tZFi8osUHJM+gbZhji5jh7imCVW7ggOi2tSTkiJRAlN17B8R4apF0hn9w6qhN
9cDKi7Wo+CMA+4xPyoQsmdLcmMbUmY9asMSVk2WlSElBIcYgpT7i6/KMYVvfaTpX
/c++5YL5PKdySz539zcKJyg2HrQVhmLPw04eE7NS3yXesd5iBaUfuIQPi1rTOLsT
sXb9+OfFlP5A/66i3BfH4kgTkgHv4xxuV+VvwiEX+L7qflGFiwbBsiwOzgV9n23c
Sbgy4jQiz9PCaszGPQdooELyAozUrW2QUwX16PMs0uruVWraR5uV5NlZgGletZiV
CwnzlY0+6AkXv1t9oR7aLmJxMkMtgQN3PQ6JMNl6UyXbsUJKwcVwVf36QGsM3O39
v4Yvlmym8t5ojvHw5P3aGKH4onkRbqAI7ffzyy9xvO5DIcpoBPjp6P9q6mzvXYHw
ZTQZm5E2waCOki81JX83Js/MVo2jgVEj8ctWPKOdG2cK5Z8t4/DyYa8ZuS2YAAmS
BEj9m1Y+klTunwguBH3SwjNvkIIjqzyjHl+GfATLx+v0MfokMZrCojtvrSyqTR+R
szqGVVQrXWqh7tMbZBx4tousPQQBrGK3J4qoLtPQ5t3G3EeqiaR1a42rlTmek+0D
o7cl3e7D//nWozTJ1GO5ZW4MGJ6me9hIFGTEEZZNkSj1jPb+XdEkkdZDns3pkj3m
6cgwlqhaLBobc5MVW5+qUyAKd7fKcgMgi1gBcrHSx3ge8cxzSYuB5AoJflaRO9aj
Bh973fx6JM1G5CtfJgeaWwIkxb1JTUCZqQ4+Y5WE7CVaFyAz1HoH4IuQs/mrsXkP
tTQ8hv4v7dG30+iBPPn5euodurlHlkhIoD6pTySqNHGWzVUegfVclrMvhxEjck02
z4d/dCOvakt9A+L3FWIgylLbGB0g4xqhcVOSOp4MYRvVU1DnFuWmrOTbWpxBTQXH
wlmTMDiDZna5f6JTuItlnzNpuIbzqrxQPWzo5eZnXccp+auX2FOfnEPU+LBRJ68y
1jF8eqRGdtdstrWbrNGvJgIi8b7rHrS9FXumguHTzEdPWXRFOf7aEKyVbSZLJ0GR
4D8HkkGOstVpHCaRgZ95ZYpBeMVP6Gd102Z3kbKadNyNKU/v4oKgC3YVBceDtwwf
CVKXhfJRv8vrcSsHy/z5XVek6H5oemjbhj6Uv035N2Uz/hjz9m3S5up7OsHafI1l
XnKOiEV41gW6EQ7GzA5JE10m53tkawSED6uHgJDXNpzV+jmAnsW2CPQXhd533vza
pUmv2yPG79I60CrNWPm0VyXzrKrnvf0zLT4+j1T7HfzzoRX5b1Jr+6bxX2A31nDx
Vy1068UwXnFOYyz//RCW37yWwSzg6ixPpQXMi9XC9c/93ddLUvMw2asrz+yA1t1e
wNWNt3ctkJNtvk4GiFkxjsgbVwvVgKkTp7UOwz5E0+DO5JMk40VtMJBpYY1gc/Kx
Jrb5+/vLqHWlbKkMk6I47+qRrfSDQvu58MfVCwHvwa8Jbhr+d9CZ3CZbtrZcDB7V
w/gNcEi7Qg3lW2UxsL646haJx9OQtWheibm+eeS7bdfuRI2Q5/hIjPbfCtwR/OFD
u/rxAhc5z689s69nxmf2rZNkC2OWLOJLEE8PFZQm3Su1LwFsDhg+4yNSLurGwYom
nfuw4it7wKZ4jFH7aJIkUBksQqfHr0Zw3md8uK8vpNZINxH++17qz02+tlJHgEmY
hWhQvTVJzHs6D/zYLrPveycO7zBEtKtpdfkUsnOyBrP8iKYU/Cm8l+don8FRMlBG
5OM1e25awsw9Fp5rQjkjIuBArv8/E6h70tsSc0u07bZf4N6t9LvuImX6a6VN4FoM
QuKg/htW1AFRDZeeXcUdXH7LTH/aD7fqpayPnEAuq1VyMrJm15o8TId10ndIjxAw
2IKnI0A08J1RSNZaCe81HeeEoaQh0kguSSLlb30+0U36xTWKAJ5tslPMsR+FRZU/
+6SkwBPwkXUYHC/YzOuyw7MhF5ZU2j+bkyBoJlAxxPQl6A8s95S83ks6BNmYjIK+
52XQLBRPvycvtjHOEsS2mfHoqWfnOU9aQYARFn5AwlD5DpNtTqFTyF/XFQGxeDtM
xFaLmGnSqCPpkfCzXOLkdtLC80071cQlY4aQa7sQfa2vrrXhnToS29HsxaqPE/FN
9PpUpoTHJyOCMlBKQI3anZUUQITV9T9TPKIPpolnaxiYqZ3S4KoJW6FsGvrSgLk7
w3RzzBYrctIw3bhI5VIdRO8SHQSR5zgrepLihgoUioUztDlcZ2bIJstV26yudh9n
FJGO4s0UEQkP1SQFNw9iKwCIvikDdfDYfq+yjPk3Oq2wHMgaAYc5/ICol2hyuXKg
UGgr9gwgOPSkMJ8FgNuB0eiZSOznRpe9CpYCm7xCwR+tvMVZWo4P1HY9opjRjRAS
qUTZqjGm2VrLuOe4aqYxZnl4uUOQtpqcM78Xelr+emxWng8Szae32gVDND2uvmiI
IdAXBXYcfjIr0sBAwstSdfj8XBbna8z9vAh2246odxlkpc5JcejW1kNrmvoFJm8/
KNMlIS+i+jtLdRHcTC7T6dEaFYo6KHb3ZlUT0QfpYKryOIqkdP+U0fqxs1+jJSOb
L4zfycTA9LBb3NqGUrajcgEUbh6+xP7YpwnpW9pphJ4uqP9inmYFwhFPWPzzRp3R
gZyVlbU1QKQPp5KvsFSX16Px1lqTbQxaj8PjLrWwXmUKvigXVlhw3MTlhJ2pEdkp
6/4nWfO8Q7MV4x4nSNRcsdDaCmbmZja4Kq9LSOeCGnNeWoHBvBP7rf2yuWOOC1w6
zIc2LjGjbOvsUjgVimWOljwEiedp69Xj3QnFTPXoNKhh8emdYMTENhjchFXg0+lF
9FeYOY1ixhdTSZLfgVMklpOM4aFKerADAV9DoWDQCPbpqDGggg1NU+y6INQt/6EW
YraqXu401gLrpUcq061X3Hn2t7EVgmvVOlRxwP62T0dcqA6DLiDSNyn0wUj86FfQ
4ypmDwWUxo4z2lPJ79MN8iVQRiGianxX/Of6Rg1UB9lNaQ2mEPWrkIJXiylJATWZ
1/PMT2tvEMWOJcOhhYhCGKc8W2mmVZSdGa6s7Lylu7hrViC8hF9tZzFDR9RxoSG7
H09A/Yw43eIJEGeg59BQLUFmhht9XJtadQsrYiq+QdAS/nA9GDdkHpkr+p9aeWON
BZzYiWfI9rZFaFAY70/CxK3gDRp3jnBILXdrx+ITJjL0pP4MQ6/Psf/hQEl8Axjy
w7aht5ovaO0HE/lPyItdfKVpGNoPJtL2wOpGpQQ60dUmx8yCHowC4Nl13xZV9fER
Xr9+eI7tMCtOQTsGoG2o99mWxzoQutNrxf6bRQ8GktL7tFjgj9uoaYddE8t6EfR9
Y2J27q+MjIOK9HLY4lB64sDEZJitsLtLHy61Zb72+neyEDVR74p2iF8gWm81HS2B
oc+V168vXP3AN5BqGSsOhayGgJuOSYs6RiBFjEFvPr77a5edKKGiQgd33GydtHqT
aHOVd9vQiJV+MYBqMSvs8/VPgQvmbNtoATbiOY+vXtNIObldxZfDHNb7CW6GrxN6
C6r5fh66rmA2N3OXWF9wP9hYYuCaw/Nqob8naSJ5xk+JHEKvuOv1eZI2LobtbEtM
d3KjjpeeQaaxYrKwQBRzui/Mo5PgxhY3pDtOiW6rnXXtK8K5CIqzCqaEPqf/njf7
b8/DAInPmDPrXWJ7dZHty60uhgvJSkT8/wqaZN09euh2KjiqYE7wuoaPxE9V3ncI
XbwlOROoJJXss82efbIYkw0em5zngaHmb/vw/p3EUfA1Fuoy3Yz2FUi4GMFL1hlt
wcM0KM+VDrQDiTw2V1G0DBkaQngYBfrsQb59AGYrFXkVQ/jjKYNg+GD6dYUYxDAn
Rngr+wo7Jsh+rz7uRuNuVMGZn2mBA/wcH6rS3LOgfAAxl3ai05KNODf+3nnFxF3W
lA41LDUCwyiKkSyzCAFCF9l26kRuzzeTtbt6+6JaT7Vci5Noz43JmTX2IZRGMrs4
amjBlkHnsDKbBvVIc3j+ydhvJWqc/8mOz5IDEpUu+rZGRAAVRrxq42/7nthey9jS
uc5wgEVpbc8VjI84g6kesx8L7KtZqoL37iePsgc/O0pSS7zMHQVE2LgVjR7qUbiP
lIntqjTyktq3Kz+xnG5vMkp/a7u1xP/+sJr2xjDxazhz/4brcZkYP65WweSsD/p+
HD2pCYwzbo3+xOLRbNbNuyNZntqtaWmJAec8YjWUy2naqB4l0r35NtMMW8n6p1CR
MARyizli1e2sDmftaJ+EcY5b7lHmR/LAFYr9ZouuYO2N92zgoj0kkmgOmounjohg
hdIar3YHimsULJFRPhphtnp/L6SKXIvjPn5+7MHJL1dfVXT30PEHvZhLk5eAW8BO
Jk5rQeiuzFofFS0Y5bwNR+CD7+irFTBrQlsI27DcTF1eKYwe9xbzyBiHrPMhgMoS
2Hba0m6TS+zBQxAWHsR5H5PrZaH0xSDRB/zIpjgztQmi8PIW/ID90eyDgg+MQOoF
IYoUO58QEHGs1nOzwn5aKD3/OZgA9WFz58NILVaG5Y4lLtwKAUZp5yhziiU+wInY
KHsM1rS4l4OrpfA7uOOAu/CdGjL8POQw4BnP2YaAKkkqtQSryQzZPbP9+0n2pKLF
RbC3prorOwk22L9ONtii01PJLRICFohZ0gGe1QaQPUsHT1haFod6I2T37B6XHyfm
Kret2xDg7P1GHaq/hmPKNnu2c5uHfJ17AD5TQEFWdY/hPaxAG4+a3uktlRKa/sA4
DAkLNkbISNo/CHK+KbOfAcd9bRjkm6bb1IXGdfsPKB3AwDOqOdDG+49nY6F8JUny
zL4lxi4zbXq6hE0Wv4QzbfsZPON088IPNmGZNpV175CJY/34mwnTNC0wTxMXiGDX
cLj4DpXIlQJbtSc/DBLJ+UD0eqotz7cCJBzK5aDH+EZCnusfvvvuJCUDifkGATXg
t8P/aoIXrOZQ1zkwzu3LiqWEav0Ws++3eoMDALum6ldJDKFxfYCQju8KO3jDES15
WIETH3eXp3zQUN52i9QSNSkHstVeXzpSZFJhUQU/hLd86bgWS3xLrw5xXM4KRGYk
a963ZXjOJg+H1QEeDl5rfvakjWNSQn1JhPoUSqXVw+NyybjLg3PP5Car1ht0DLML
BNH9C+IPn4XZ0lGxk8wjUMFczd9L+A0nQa8R2pkNcpYTuDYxIWWc4fS37I8i8eXp
OTiwCFN7X+c2Nc5egD0XQVHNL8HPdgMhVI5/dts1pExD5ybEOe/RW5EcSyVJGE07
HRwV6QtNXhXtKVFqRzEHFNUyy1yqbgMqJ1vzzfpHfPPVauwKSnH4VYRJi6ECLrys
Hp5I/D9bgdp3mo0ZjBK/ATxSXGJY2BLoaQXisPup1dOOHDhvX5PrmaGfcSMKGRGE
vs4Wf3Uk91SLTlFGBrlTRXzxW9qYNmBG/oonvDG9ocqeFWsXjoeySyN5KwlTiXf7
976rbeXBK2lxJY5vU5tRIxyZFFIgdYeAMN0es5h1mODmuasZeagM3oa5pOYVwmP8
Qhv7sefHO4G8VsLBgVc2kMcQfcFurMzV3sdijILgN7dNcdI1q8dKhjXdH0x/57z3
VzcsUaracUZ//iO5c+Q/Uor+2U1xJg6aqSnRLrlMzUrBgSAExIIXOMnY/dJzBZI0
OyuwTqXjtkkvj683ktrquTXf0ZFqj9MX2j0I+EFKBfIqDtuGZ+6BfowJ5XT417xq
cWEokiJn5oL6FJ3YJCVaC7Bf83i+j+776LWPpt+xPDoszMZ1v+n1q7U1OYb3fjol
2d29d6s2O3vMjeLNcrCWU4msZn+2YhktYygRyQM/tJZfRVRcxElZkbAWU+RSSG1G
xIAo13zZRsUNN6kYGzzxySFbi+B7UdqZKid7vu/JaNu1my6/zVSZVlO2NPD/ugqW
nxGwuRWNbKk6T30Mj9pifO6zkNSllAyea/lzZB5cxYm4lsNWxUVqJ7ol4FGQBQap
6H08XMBqxN6QzgBVain6GiwmEhaL+OFPoneYnYRO4d7bucAh118MFdFPrqY4umAn
OElVO2zBOFnNeNylvKrzozne/KGd77mlhyU8RVaKocHHAlSE3ZHgcf4RllogISuF
wWK5X8jYbhW8kpPk4o+jk2ZYUcytGrfzAROB5KCcAR2c83fxBX/G5svR0zZMFf0q
RlFkvfgH1rBoqm9mM3w2phk/9yVwFd5s8wz1lhZSrLDwGGobJX/Zep6SbR9pfv86
xhaIsiTJuJylMh/o+1nvuuevrcaCcKF8FqGGlz2v30jSV9Rdaw/gFDMI0U789h+d
5Gwj3jMA08i1qr8jRvhZljvlfU0Z637sbxaR/9CSEGJS/TQdzE6vuJWu3zDiLW26
3dSpImQFXxhXPZdo9e3Z8/jVKDbmduCd94KMQPwdUZLtWbc9koV1vBoucq9Jg/fF
wH3kU44hmOLX9azldZrCHBhTzZRCtDbLW3f7r9JYbfak+KpFLyugq6Vya8RL5RaW
HkXgBhQhASNMRd6mBwOgkivKzt13x6X3WFf0zcNhV3CBInvr2Q1GPPwbugTHsgDi
vZrEyQ2cdo36lQQHYzA5D1q7MKP5rYVzIgC1YYiqChHaRCLY3UgiRnaSOYQ7qwV/
5sKxY6QN/LCAcfor488twkjUKL9WGcIOvb5M7bZenNEAFUCWH6v9WV7qFvlXPBsz
i1e3xxaxXFECFWZUATyqV/LVA7hq2ko+vZlMwcbMl4iYzxnSdaXS2JKDaNTfy2LF
DWph0jWSpOexV5/mEsf138mSPGMdab4KOhJ+Zi2xSk3qQ5D1XVNeXtRJvTj10pwI
KejEYrCUzgngGBGpR8pgRn76TqjIOJJDXWc7KXf5GbFddOyIVC2C1BwdC0EubmbV
8u5i06LvOsWBGQ9mZYrDIGr6TFboXTpTC6irEasIP3QdZg0U//ruY1X+d/KwKNHg
ZLcwQ8sLFJoa1X7WUVhw4JMaL7XHZfawEc7T3+EgfLZxkx62+pZYF4Qw+Q+SFO9Y
TylWR1Bh1UU+7prDpEjVtosXM39C1L3HrnWdw/a6kxGhCdEbmuHuDBkWdmvrBPCa
mwcW1itpeHVKu6JtYfOA++94fw6imt+fcQT/k3prp8d50y0/USHoZlSQwSUBWNa0
icyQO6jbxz28Ru0qQjl8xvUJgicp5WEOzXGOuzFnhRWOu0JH422hRtuevV6pm8h3
abxRHIWrhc8H2ueYYNW3EgH+uUNncICxwcu8xRWm3hdca6krw7Svk8kzJQky8+OY
V3m6jekHS73SOS/5W3S3B+PrmALgHHxzlV/dHAyEDuGC4Be3ZnGNXPwvdCrhQHKI
S7dfHsTJKCaNoQ067b/yrzU+7tyfVhUDiWgukpZArdh6+43u4udFT8HVXwMI7hTO
2NFjYx+RRn8D0A1hqKVLt43FZQkrjJEnb7mu9J7MvpgWewYDx59b66BW+2El1vL+
8KUl6UdrSGWd4VRZBcBz8YOyNhL5ik0OmqiZD53qNoWQyRJ2tK/U/TtgAK1DQraB
c4+9RE4j6+VZ0VFRV9YaecDTcqaViHeei/hHuoOYgMu/kxQjkz6Og9xEMMHXYqEX
vskT2Xrz3k2q7kzzj0nLjUoUH9Hu/6UMTR1p1gt7Pq7hguvdDFsiFe+EK7jqUuXN
2ZaBRbVjV1/S8yR7vWRuZKQwU9UQ+ynZeAPeZ3ItMZbDNQKyRFMPIWWcaXaFYUFx
udOZUy51NTVdLTxC3wKo4yOM3BqtV/FJMun0BpuVFnU6ScLBvvgfJTfwsRC3ZWFp
j58GiDlYDbzBvjr0HFfdE7oaT5/qfob1SeeXVPZ66/POQR8B848k/yP73k6IB4pF
q+Y4/LGehFjODu3DLdQf6j43KDquULR6Tk/QLpOzAkTx2FAZUTpPgDCS8dmEIPjg
cm849umxi7V8cE67t/FVkRIdwlX7HjBvNbuBMaKo9hM+yu8ARm+Q8vIr5h5KExVw
c3Yuu8h/BEZGFj3m6getJ6j6bg+kv4QZhz+IygxyFC+usjXHfeq1M8nSbgm3B5rN
nal0ijHl/KlK9diIT98EKoudhmMkG6hP8zu+Od3ydGz9/JSZlUKa/jwGUaEXvgCD
Shv9hdcggjBiZoC27mpsyvsprhVhPfr9HuZBCPZeKp45ys5PNpgoFqU3RPiNbx2U
qbTKIt6tqfHeD6UspFO0zcJnzia/DHCoUeHmHRKiPWOkkYD29h2AzWhPDU5MSpVy
5DoQ/bK6ybL6bvK3qOp0xUSJKonSzVerSsq+Sqw1AZaLpTgF6cpgsLExl3KHb0z9
kmSVFTGLKmsE4Xchz9cSmyfCO46XAa7Jduxj6IwsOB/PUfzts5F5B2qaoymILqWn
bzjQw4gPyi4MhXELryryg+WRyHrOWQ7tcSsnCO+Sr60g9IBh5F+jXBJC4Ewm77xO
Dbd0xY0JJbIP4j5+odl3J8C+O0HbygH5eGRa8wRW1V7rHVdA4ur3SQl3z7npMFa1
5SO3rkHazQqCUbiIRePXT6Qv4aSuYlXskEKXREhgUxgXzLDXlRuN9Laf1gFTIhgc
Q3tVv+rEnn2d1XomBiXJap1+/pvEzW4LdHMw9xiBRMAPrjidI9X8KC4zjygTwDY5
BHS7c6bRGO4eg2ovEjYZ6jMn2IPikiQIMXeJ53C19iLzZJ38nIZnShUfXHpPpExk
SJ6kpB6egnMHkLjqklWq5bDy/1SzdG1bMpH8sATmvU1usttR6D/zIfkPMn3qO7De
P/hlqnEy800COT/Exo748hRaBlV2bx2CsyBizj6Eu1IFaCDAmghFXOOsnxQNeN9h
Ux2eUEkBaKFldTDl/SZhXIISUJovuJnW/NdqMcXllT6v7lW5NkJa+Nd2i21hCSIM
YcFbM0WbjTAjz7Rw9vJfRXa1cvBvmTLZNnHbR2K5jj3xZABCy6n5+IH+q1hH+vRi
ISq0/FVijcfnuDc8R0gbVobDF+TzH0xi39+t7vB/3XbSVcFf5kFRTDSjkEkw/TSN
qeP9/k3RERUPCsQIsdZBtNeKOxFHq57hUVvyGrLQURT1fFuyRPsiAmxfsKOTUYdJ
KxqCs8nV6HAH/Uv8Lxi6d1GPU0ngzVXZxqS5x4C5mH/3dc6QcDBKmkEI0GVLeUix
bqimX69oZ6AvK5YkG2G3ar+1tHmD1kyfcC5Ecom09vK2PSzQhvfLO5xw1gl0I7YQ
Dn3nibBTGYNHnoHCXVO+TkfS9M1DymYEO5G+TTrAdrpT4k5mg8GwmunhqnA3PcQa
wzK0ZXG5UhsG0IfVW4OR02EdVhBD7AgNLUrrRHujePg/lgQZCbiBt96FSF4vahGQ
8Dn/0x/Ds68mgeoJYt3esJ4n1y+5mL0nJSFRL/p4UWNBAE4TGgHbALeKwLLxsQho
ziKDhL3oCPpP8TpVBiYf/GMbtCiq3+DZIqyg8ow4yMaf4cX/Mpg84jIYMVcPrfSy
aZ1hy5it1W9BeMunB9Gjkgky2Om8dvQJ5iFcidAVE0bcniZt8FvQdsVnsa63FCNb
5HC2ngFNsZfHh8xb8SOd+QpNalR/8OpBgyyofx2/sHi/ZfyjtUmHQlaypWuR0XAE
Hdzhwn8iFnJUUgv7oNXGkPIPfqlC56nMzRAISojCehkq/cYUcP44wYOKgI7OTnFa
ro3Y60AqHLhXC2zkLMb8m2dps/IO19EbvR3qQUuBrWegpBe3xDrxbgWc+SN+SOoH
YoPOmlWLBs8M2NLmnQrSR0l4UYCjERaYuRN0Lc1ZzzxL4j8QcF2Nitsp1zMwLiCG
j1+B5DNDSEP7boaDODn9pkah+Ua4Vms/FY2DiqKSWq0GEw9stl3vC95WtLV7uR61
l3qj3PDuz73y9Whnl1ZONMF+j5I0GT3rCvpUFAB0CVHT95VcF3MpJtEyJ+BIIpKt
N3ZK2ozgI8Kee/K6AK79sFzA9nwt4qdtIQcr9rC2kJtdaeA/qjgIHuLL8uKkMdnB
/kOd8hgrP1WSGrwFjhgDa5fknv7BybZdNdZcl6RjTs9L87rOsy7oZhdZ+o7Gf50U
vuseO6lLtLFi0kE7Kl578OrWEhZIYWt0+B/N+j/m4mF4kfF6EaKkwl/u3MUAsmRB
jrGIYwUObTM0FGl36x2JT/jOG5h3GgPq2Myw9bSRN06I6HOEwtx21V+EeyZIZ6pr
6cntHv4Gwo/B5ta1/40U33WuMx7ZeVO8rBTGqFuhR5otJo2Pf2RAeXeSWztfvGNX
guPRvUObxB5guYsCzToPJvh2mnXswLlZov3JSWsX+w+giL/bZjkptObnNwQ2je2u
EwIRlbX+fONcMixItZALFgkLMEeISx0lxqIq+zGJDXeHV+FQqsLiMZyPolDx8gXW
WsgA100KW9slN921FdgejvBQc7J/yB9Gdzru8Qabk1U0xQI/YBL7p2ovm42Tfxgm
hBQsZ1Z6HUFvhAgMH/zY9tCmR2jnk5iqQGBMaSiQSi15I/oSdovkOLGPXJDujWHV
AnAPd35LP+sRphXHdKKFW5o8Kai/Oh7YJE3BMWgpabEAoXTMfy1biT2f6faq7n43
c40N5rAfpA7VhziFV2pouwJbn/WwFyyYI8hm+vUiHQZEsauLSuje6BGJZp5OuaQZ
+8SxLMKeRAusAh2CW0wupH7eIny1N3loZFWeKm5cAG905dARLJz4A9i+AemheGZ4
fxMEaq3o/FN5Xa16D41424mWN0LfeI4dZYLViV8jIqUF7i68D1z9EPJMrEVB5WWO
cuDU61ZsDw7/bNoLWamw2j+Dot8b/Vz8ge/+a5oHkGTF7eALi3jFgLr9R2Xy7tHn
IeOKc3B8mqvi1Zgrsh0/y0EObYp6uGDmXwVDlDU/ob6iWW24zJhpObsH/+bS9C6D
QgXGa8X2OkiVRDHpQ+4AfWQzJIsUijvKwbx3iYxwG4uclNJwD9lO07Apmfa/AJFv
w1Ng4nmPBpD1x9GOjI0EI5OFzKCVotEdTNS+PxJE2SDnkqsUb5wiQeVDd65CxYEA
r4Lwll7CUp/vwwV23ErVG3Gq0mhWmEOyofkjSxdEBCW5EmABP1V18m05AHYbKXGJ
K+640LaR0C7JueOhZUp63latcCMPky6+tUNmZwnKup5Sm6QxZEeqAsbW1fA8uytR
+f8DcZrzU9LeAEVhsims8Qwe1RJ8yM4ePVShy+cpMk1WMVNt/EF58fRj1wRL4Y5Z
RmsdsW7hPqmZz0sJtqnGFt1dJ1zm+Xjr0gQKJYJdgNwZkOOEw1eM5gpdCAMur+9+
tzeq4LZfCQviN0eDdcF0E17fyUBHkbkFYu61bGsSJfpDVT1nQy7HifSOfXRnrV2C
9WZe4skwsNKv/J5nLbk79NL1at5UVxgGfpjTPTc6OLD+//Vbb7JokeKViuLXw3Lr
zwBtVk6IEQQFf1MqkyiqZrcP4VG0xaReYUVQuj7TjSj4f7YhY72hyqzUGnkBfAzf
0CFqiGRTIFxnF224SP1GeXtA3CLGXPVWxU2fC1f5QIp2rmVxvctVvt/CHQJAYlxR
/96ScR8yxVjqs7M0je0nWw7KXvnSXaknhHUgsjKhTtATvuyMU3v1w6f0DhSiJmll
UyArMIzHk26bHJLHxUepA8aIfMKUlOF2swUGe09VKocBNutIsn//qEyh0GGh/Y5H
IUeyySAxsJlfGyZujMUxw3psN8munlB4TjUcpRJ26NZ1eQ/DL1OjZgrEf8Y6VD/N
bV8/FDpHrBXugkJpXGPHihleJ6Ql4O2pn1LxPI3ziBwrOCZ5FhANNSFoYNw1HdQj
U80wSCkBUr0MdHCtNGUQlGBSeFtrLLDFN5eWiABi39HQDa6ZNWPLSYIhV7XjLctv
S2kPCGCeQ19qQDJM6ue1PzJB1NgTS40M7T23YjAO7IeX5x1ZpDXj9v638LqNrxxU
41k5GL0FZ079LkIBRwx86Bahdg4ShKJ5E1PE6pamoib0kTWvWJwEbmte75PXco5q
sZlnYmJlagDZngp8/LCsZMGws9bw+SqXvZIxru5Twi/2BwvaJnM51t/aXWZzF5HF
WvrZ48SqLHTIS0UBKffioa913dt3pmdlQ2rrVz868WlgIiEGzQ2Ap8iOpl60F73k
y5AFKEzzU0IZpibsDiCwlp+BRONxQE8JOJOIyPky2nWotQ26fm1ICpU60un8zguv
ysaMmwwpMUm2W6p6p4aIFyT9vvBlQcu3Gw7KfWT9+9qbqcCnW5tFhwCuILk1V2lY
kPUk7dNq3TRwWwRY73H4tKfgxLRHoegpn6dVzAoMFhA0jMdIAblXx2T3j1A6+XX1
OtwZs9us/KL/UzgUPzvQhnmr3RtDraU45CMEMsofPA69eSjVqy1XQPahG8lEmbEQ
cjpEpNDP3Cr93zYhiib4IACrlcnPmfRPiw1WVMfluWnduIp8//NdVYmsoDDDxvg0
gz1bcyfchBRWfsIBjiUbWvStido0Bv6urAHlPacDw+MG7oqGmya5O8nkCvdIEu8h
bw8nwlFSe4+PjXBAM+joyVX3WhWUCgsjDW1bcfb5IZw0i3/Yj8qIRtN9vP54XNca
/73ymSHSwtYTMdLkN7OUDcsZzL+vU8bPECZ2l5KYHs1I7UVR3TivPfFemp9k9Qyn
hj0sQ3Vdv2VLtg/jyn1HfBsQhfq9rvda2Z+1GVOED4QGlgOFNJljiwQjIhfT8TgN
siMtwsd2/aKjQVhSuLbUzXj3suoepK1yMmnofTrxWEROpItHH/vCGMAVVkVwkz/b
a/My8i6BAfajsNu15Jwd/WZsqpWEfGiUhZwkr6vpja2gHcoUgwxtYJ7DFHJRzWTH
R6y4NkH99XJTKZAftbuZ5x2TkrJeYgrTz1ZF9XrldCzRXOx8x3NBK+rrNNTwcon1
pN/7I/CSNuJ0jJXeVaClmnnL99aEIU+V8+hjWgIewazShOYqB7HH7pzYvHLGp+d6
UM/e2Sz6NVlTcAzvFPAiQ4cZJ40XT7xO6BIRenBHO9IZ4fNXF9DvMMbYAveIFbRe
GZz1ICZ2z8a73XNo9M/ueFzRJ4bnRyEUQqecbfeTrbaKN8eiR2lA0cxlM2iOe/D8
uuC5tke041wpWLdNXBqyclPzsiyJSP0XkU9mJFiBIGa1aEs2J8OfVJG7ONppvVUA
Iebc/l4DKQIvxyZ86vIzrL2QxCOB65jQJa69BnG2FU1+7PWGgyfi5Yg0GiTsE859
Ss6zjXAorTt3HMqZzbn9kvO/+MUN7ZzPfg5rrJDD4SmfEwDQmYI/6bMnigNXqNlb
Hcd8gCGDrvjx35OjXQKXE0ynj5UTVkhZxVcd9He2BFxeqMdFJXfC5R5tq1hGfqZw
Ws9xb1utv5Nn9BojkcG6hKUDJySaYR4FKfHfRW5hgpziV7KN5fzPBSRmsWsBY3Fi
mkrZahXDb178uyiggo92/IgzgzkKBhE30f89CQ1qSirVGkclFxBzVs91eRmSOF31
9eq9CJlvk+hY1kRj+6j2NC/UJaT6gHbzaZrt2LnkQFVa8zrsI+LdSTfkOdHO/4IR
sLdxlGYbBI26V8VjMkcmljZyS9xQXbC3zABXdkbEYoN2OI1SyXxfarncWlP8wFob
VK3F0YYxc9TNYWzZ6O6exNIfw9Z2Bi8FmTwM5uArDAmXD56TNGRRsWIdQXTyatae
ACW1HHgbPNC3qrTlmaULQVRmyscx/Wll7T1/i7dk8hBTODJkbYJoPfeI3G/4HdIe
DbX1hYpp89lWC8fdUnUb+BabQz7GqEzwCqfqECQxyS/iOhaOFqITJpCff76uBfIq
ESs0n3j9c150b6GdHSzgAvhWe0DLnv8Wj7Y2vY2bRi4F7MikkLiT9Bt5Jpay6+Hx
MvEFyoJ/f1uMZeR8lVZaP6fmhv1hXJsgsNFyjYipOpM9KqBU3U/6Z89KvPPRKLHS
FKiSwNb/zSotKPuekHb5jg6cOcWmf4jpezpJlztCQ1zqBB3duZj1B3GG6l63gPHd
LS6UMkfKQHaPApLS8BxsUoh0cWRth5kkf8VAwcGp7firMDZV6zi/CAHu+s5G/w/4
ghgr3WgHngM1j1/5GvtFstJ6bfCsPrBoVD8cu94W1Jl5GXCqW1yWPh87qtNx7bf8
QwysY6PbYVq6BCiTnBvm1bfb63HJf6w61hyVThRHtHaU266IvTNlPGqezcwyrZyT
jCryHjTZe0Xvj5flf2WDzHcQ+SfJolUYQYou6XkX9mw22lc/HNVLSAYjdyQUCQNK
Anm6U0ad4GOcB56U61GR2n1JgZAyuLzVn9EgYdajic0CBzSsiBSMFW0SNsTW2oCV
n3CujfokKpHBWJbe12lZaTUXVk02w0vw2KiRqgznNzd8yHbfeMyIL7XJufHKE7E8
NLmDwbAyCF3jWS9/A5IQHbAwEudIqw3XO1DM27TpbN9aYrwpBZaK5r68P++6WG4u
ZJV6OpJBaf2uxWV3/G/hhtE4IB7pbF3YIaIt/72D2jSJ54vw0WH3sVPscYm3AWmT
8PfGs4HSlZI57ddge7CJePCYDoz+9Del+LPjNGBaS9GlyyRsM/yPiRow9bsYfOh8
aAGcpaDstbVmeMZ78s8buQWddmL/DVsnLOZeKKWqMBR09NhMavcB+gGrDX7W+8k9
nEv+1Ev7dk9ky4cGKRzxPhFOgGVjM2ki0AbOucejPpZ27/o1WOIvUDpUFCQ6Zu43
qH1qmygkb/C/jg9UOJbsVg5/QMezpOBfbDb6CsWJLLIMBv+W6eWpaMwvoXNH7Gij
xksys12rQ/K23VGditOHVFgnNinhq9KP0krZ80zsEAQLm971UmzpdcvxNo/RixO3
WajsxMMO40mGKCg96pZ7vS1JnsLdJyAjLtfg/UhYwRT7qLUBfqEZdBb8P0LEguwt
DbKJ2XgTffo3Jk5DKASBsHAUO0lYvLn2MtJsd+F0oPUTY9mmZUvwDylvArHTVe+C
LNNQQy5XEPzyuP+t6hZKQSi79JIm5G8/4o5KPyPWGhg3u08El27OpFDKQQfonrDv
Jw10N5aCLK1LQyC1ETCgOQiJcn6IGDPXWBvxlh4gNmVkKgjUqLVqmP+atM42EP4D
r0Q1l8NFKww5z+SIGBvHu6qtP1hf7I4x9DCCMVVjnWFsPvYR4f3wF8CDwe6e3SL1
O5Co7lVCNqaWHo1Ajxge6wLEdfXYueueqsTgBHYB0q3FT9wHVTCRZa3QhT6nx4oJ
NMgIl27up5wnII18zh91SdmSXlSaz2rjradZE8AW7L+3rCok1kBA8pA9IicfE3O6
209wmvIuFkv1KNhyE32MgldOa2rbtg74pr9nWEReZ/67ac4qTVCO7qdfc/qdcYCU
JwP39LMnDYB3CdV+ZXoPj48l6s5yFouL45yo7hLhyKd5eQsGrdcGtYo3PFL8NqXx
RiGI3Oe2s1mHPQYwkfv9qkRCDmSD4dgP7Vb0MHmvugtBf5tN6DO6jVnDYfc1eWBq
o9vPV4X84sidMk2M+SoOm2MZxD/Kse1CVY0X04j+jJpbDZRCIky3V7nqe9qOSTQX
gMUMa6zPgcJ9OdWpZLvvLL0FZl4ofJ7a5bVCwQ9YRG3Ak9unNHB8W0DIBUJUpe+w
ZvKqJJu61iRP5oUR1DRLwWPqFP/5LNckrO/86tN7nEd5dApEDVZzKtzKpQqrRAxx
aD5fOWp8kKm9eFEIoEDwAdvPRkViU6qF2BbQNKJTSlLwwrCZbRtS1tNOASvlkSBS
/FaaxiqjkGAX4t7or7WUwF8GdxzxKIKv9ptkJH67PGycEDPeLugP2ZXJuiLNnFWr
WaRX+YPIj7+4CBdJ5+bmZTLMX/p4l4asWKabxxFGhs7S6Hb5uk+BgZUpNa4AzhCy
/MqnfyFbmAb0MUg/E2liZzmH+MaQMh+LwZqg7/vjRV7PFrhUf8TIW4pzxpm6iRPa
L1CTyDHQC/BrwBukFdt8dl7yecC7+u0EuVrY6QCN+bXqzx6inW8R/FrsKnPtog1M
9MmUtWkZMQuJJX3DASQyRVAE/Si8zwZOeeORsmwfS27rIvXrZvrDGrXPCNeYkx7d
bMDoSq54GIQ3M+aWQhoH33l2E8YGjfq8nZyZ/2kuu+cwm9uF9zabthzTgUH9BauR
XrqVx3q1RBE/tee9ZkNC7FBscTXgF4UwybeXeA548/yYfDMjPpaGO3mv5syN7l62
3M36LCAIRASao0dcYRnVkpGkLmXg1/aDp3AEeeeFyzcQmCEvKL4zWtdrPvo7W/oG
OiLaoyvU0++3NO4c0oSQrTF9SFs+2T25CKPAZ2+3Vzq5aRiJhTngAALTBGXuEsNr
ZJAirzVV2/baQmv3YW0xP3iRShSD5NjlZA4x7MOmk09OTAZg2MQ/WSu6BSORWa5i
2sISM4xCucXqlzgO2WmrKZ3ZEF5iTsFlE6tK54nrJf45Wmcr98mNM0634FrBc218
tdj4/XWNEJIEJMItkYMRMT/wLxmIKSxJQjsjI61Pp3tKAnv0zvSLmvzUR03hJQwQ
7PcbNpAKMNTkqA3QiIQ34fzG6mTrpuCksdgiAPBe02IjIBGF3cK0wfYxYI7zf0Sd
6BxfInwo9aHbXH3JGxPaG5akoLs/pAl0KQ5NOCcXJ6UfRetDF4mTtnBbZCrk6XRZ
e1vvdLSaRIzjDUCC+2SNpC3g1Oz25D0hiyy2disv//zQUD7ar7/oRq403ajk/17a
8X0Xu47y94/kUo9b0OClhHAUCI8XEThCZ1nKWVtvKgkZwK2xBiDScTHD2SbRhpaX
RR42a7MW25RG5jPf/l6w7keq0Zg243q4RfUz6GMP7J9c+25sUq6XtRuyds2qJVzH
EoY0v4fMCdHBdj8D1Vic2F2E5O7x+6+ooutbii4EEG1GqAMpLJiNKQnSg8beFU6j
u4XKSpMehl6I1fZnfIvR10cWae/W1FZdI6jG3wuJB/38teVkuCQVa4BefjOkXqLy
a7IuII/YVYr5K/SzAvauo7KxhcGsN1ml7uM4VTsu88NDErd/G+wf/6Le5WCodWj2
lw8LHmUOKSKyxeahhd5ZMkFPWb9nTzOLCHuoT7MedJ2Fz8e8l5avb3u8isgxu4gm
M33gGIb/IFztacNzqQFpsMmEsw9UYKCGI7iauYZtJ+sp63iM4m/LgISL5Yr2M8HD
vecK/+VJRp3InfbnStcKr4ksQDM9/t2ddGiArywzVGmo72y24OiGBBh/iMjXrcDn
BMoAl3qSS9wx5c+m6wv4R71zJcfb9ffoTq3yEYlQ14CQcBd9pDUrRXvKHb9tuX1J
tbo9FEGf5lC26kyI0cM3KZzy2fYOg6+1YnJ5WdZTg5JHoDRr2Y3XuyPTiLTiRsiQ
2s1W3ef9zLTCnOj9pxSNPT8U0M4vfkviicXle7VgLTq/Q6Xndn3PKZyNmuD4avUd
wDm8Q5EdIiiBtoeiZa+GMY0grdAR1iIuLPYGOxa+TKHrSSqB6lblmr6pa3btQCwz
PQmpTK9207d/Pl2EScF7Ka8zgBhOIk7FdpFlZzCc6q5+obYYbdJDTVKeemqGGZ5O
o1pkxHIe8FrM8krAlgsLP210ccVZKbqP4fP/cvi4c2kgxdKV2emnE0wzUTm9kJYu
BCQpDTZKNXuF0aWzZVLbTQuXiEdW1SSfhp5q1mb7SlkpkDl6XivQd/6kMhC0dDHx
K31E41S155ZX63QMQqGHFh4NtaGa3RtaO6zT3FJ7oRY+xmkMQj7HT6yXAOXBkj1c
fqp+xB0ZTIoBpfV0bB4D7w+uKoEhFAC9dnqcUB/xA24htNnJiH4jb7Obdud5civg
kwBXkVBDdk2S/Kn1vyzsKkqTOEp6gL9VUFHgl0R0to9S/nNC+hr7nK9ZCrwVde9c
SM84qoaMyYR+SsdJ0TrsKGn9vsIQ4KkGkm65f48yrYHWCMhh2vz3v/dR1YkbUfM+
zefhRdIp7VttdJVgBsDKRL7F7QCa+3zDo7RQpw15gcsUyUjyVLEFkZlsalVwZoLd
KABY5ZbcPjNG+36EgtYfjMjyjDlRqpDf4ySlZBIvwItC/lk6lxz2fOwjctf693AH
Wvs9P2ZMGwboIQyF96+B+dqWVIPRxqC2xaZQfcB1/VcEWGgNR2hZaEC9eSbOnalH
+IcrUn2soEisFJ/IzIQfMzYx7/EFvzCBKC+cRC+7nzye6QW5Jy/Ag23ipEFOfHRp
Vmhu961+5BceU5017HsWGMwK+tLEV494J0HDdFLAgcC6ddx1qxUkf6Ut1p7i4ky2
iB1rCSc0ceMY7lGakXe/b7KHjXlWTPD8q37sYQk9hszUVv1k3sVfdttSeOF3S2GG
5wKKWjSctag2Ihc6/9pflA+wSluyqYLuQ/nbBdD4qvC1EqTI24YUw95sabv8M0Ga
bLw4e7qXvYCI3RxQ/GV5YiU0z5cx2X4UQSWWLr3ym9Td3TppHfaMvmfoUeivx0LV
X1HrJvKB9BjvgYekFDA1IjO0n4uuVdF9NgqIwXN23iYIf1DuyiEIzgcc67JSZtB7
qZMyBM3U6ltGNpkRpAgf0FAHj7OpdbopOBQoiSMTIhSnVxojU/Tv+9Wzju62QYdp
bEdoHfT/Ap/VnVH26p5M6+aZFgK4rT2Z73mgufJk45imnT/rbmBssUTCptd69lqm
6QBeT7J+eJwlT7YFVzAXKGlDFHr5cG52fTiLCzi/quL+vObqNx+dW5QkHd5cFETO
W3EPpTQhcgq4/FOhsVFxo5Lipb+SOvI5DSFzVDGHTU16tmRqliOspYDqabf73dMp
LE5pcbm3SE/H1r11vs9sEDDiqnDpNs0AJjmuYYQhPFy78926IBFQGRWsn8kAGVRv
zI0ZNAhDqKiBDwQv1RQNJ+xfKjSIBh5pt5Kb4kj7iOr+9PqFH1RowaprpsYOInEO
EKWq1ElHILMdHWeRihA0jmqlk7Llxc6jbL8VNyC3sDWrn3MMmMysL4fSOw1kVocJ
tZ+puPGnpi2pRYnCQqjqeLNqa6jX/9bgpgt2u53nQjGk5sla4s7D+nWeMn2/0xle
OEzJ8gvhVGvVH09a3GmCiui3J8vGdTdDBQZNOTJakV8yRUMLbEsQmLKUquEDXH+z
kxURms+tpOxHsLWJh6YiE4ik5A68F9hY83E17uH9gOdabnCHX1UpyzevEzAj7VAT
INPvUG83LGqvNZh7XRwx/CgGYpnTOu0J+2pQAEoRroj/fgB2MJO9Al+bUWSeLa0J
27WmNB6ryjbDCRedsTFHNWQ6v2bJfAFxbLJjsop+9LwJinhg0QrGfzbklAsjkyUh
IhsjxbO3aAIbF03XetlRcA4gn7Pym6A/wK/doCRSjgRTvop5VV9IlEbw3YjNpDm1
aw6W5YtHwgHwTNt8AtFD/1sN98aPpFtTq3ng4AndBcd0YSlhMBxINHuAYYzvkHJN
cVBevco5SvzFwEb5TVdHYA2i1bPnoZrlzOB1E/Pew59YvdWNhB2NSr+fc3bc5bkI
diQgsottFdPLkBrAbZl7KUaJxkv4p3AOeyv9gSxO1VjXemx6OLJtsoeffiv2cugO
s3L/BiIY0Hf7eSKjr1kj+/BB9iYTUI9iALwiHbbB3xdV3BylCMfLhEY5GNf4hMYw
CdOmSUzwXAz3UThI/l17mvpVgLAtiwVAnrapYozWVVv/i2e78E6vOCcNjm79C7h7
hTqtrqMjOoTpTeGbAV+uZ9OAWz3x4+8xl8NSn9boj/gSAk+JZ0kD/Movz9Qca2y/
lUnfvcmU1WkGI7JsUqgI/4inoAtj3OZSWWQwEowAvuR8qGISR+/CJLi7lvuGDjES
v5LR1OrsVsOa6AJm9D7cSBiYM2VXpMs9or6Y+gW1jLXz3zjnkVGTeIPbXFh54j6P
ySI0Vtfb/UaXBa2zmMYpcJTCvvzB2p6Dc3ZcTZGYU3YeI7TRF3YBkwxNt+q0/r6m
p3HUqGMyPgcGS2ypAt3VA51NQp9Cx7Y/2mzuHdWWhUV5Mssd92+fsDGv+esD6fyb
IDCUpfOfG1d5ACD92vfApC27TYAcjIXTswLxeVgaGqdxP7V0tKnYF53eG7NuB3IF
WqpUFk/imym5CbiCzEi13fELV9RxtY3Be165RDLUpRMQnXe+2h/hz8ByMjGNgEHn
JfWQvvcGK/RVwoGMFxM9tmju3DO59QJpdNuB9fJ30dE0d4/JR8k7iF+VFkB92cFA
TzuJAVkEX21NAYBWjJh7ds400yMOXQ9YZXiKSd6vKGbc+EBwofcs6iwflODGhZHj
BIAyamKu2v1dIaEyTvDfmOUYQtZsn+frfQ6TItQKO5bJ2hm/vhHZ6+IYmi+5SDxv
3Oa05skYv7lWjHD3YPtj6B6BcBQfFfsSk3cg6vLj5lLnpuBycq3EI3xIw3qBMaeF
qsdker2dFhPYoOdOdX3DvfP8D6opakoiKNxFf5jR2Z4ackG22CDTrpraIn75F/Qi
bwPWxfUCn12GdNqokbN+kVZJOyfTWAqSQ/qW7u/GjQbdlKL3wub9SN5klQuihb0y
Q7YDnGEBKt6+mGb2qFUR9N70Y4NRJ0LSnlHcqIOzD+Vtptf6xUqYYnS9IlU7rZrg
9pyMyBcihiAmr39DeX5vjipRrbOq8umAWTLvbnxVvVP/d35hB8SyW546dNYiWboA
bSRry9FRL23jYVXfjGXQPbgKZX2VGhsvBcvpGR3qcCkGIBKxpZursBpLYfW76k1Q
mecoVRXQXcwThfbj70IDa/P18f90AzviC8pX6ZLoCEP5esAYnCHI34t/NiUHM3Td
YWJccKp4tWo5l5zj7DRXe9wdxIycurjF0nqa3L3WWHoC+OnDe+6CLIz3Co4kp5lo
J4M/8i1T3kNL/95tHoXkTrSoGtuBtNYulqVafdO+JuQ52QYYyjKOHO4EIVo/3tAA
YqO1BmjyPmH7uvVy0nP5FJcdSDQbHbUj6gQeSjtubYMVKta6IbJX1KTA1OXMMuyQ
/84wxG6Rz/6qba11tX+temM4I03VAo/YD+yoP21kBcQiys8TjBDC1huFEu4QAYQ5
Usbz1cGlbWDbgtzLxVAE7/wRg26KPRn0cRGOAgmhKElB/3LPmg/p+9Xk61kOkUQR
L7LBWW7lg7bxbTY8hLbq/Xc9Dkzn8vmTGEWvtD5JlHQ9GDRnAOXhwEVH8RQ5aCPY
R78PDsZa/90+DTOvNBODTVUsO3SCYcsZVSi+HtpYh06PNza5FxpM3igY69Rkb9O9
zSmLqhEvScc1/5FMv5hqu/fNYlCyi50mu787E4/whjthL3eocGgoilwUkFVT2BCN
WHFUlKRZdXsBUoOoN9ziyCIfp9G0ZFs7sbJ94gohv8kr7Z9YX8DYZRlf7tpxpj/t
OHkLXJy+ETqArYlMjDGO2+eOaFO3OHqwXO8we+8xpu1aCWbQSwLxm4bhz8go42hX
3lx598r4gkgxxV72uf1/hD028yRJ+RD6qFJSQtIK0U/qHC6lDLnO5R3JcNU1Hd9M
l2/o7SCAJ5HD8ViGy3O/ktz0sozpunbnwSg9mDAg/apsirAT2D/C5I83/q7GXm9Z
PdYsfGFdy+kWXdalFoGAygf9X59OaQS20xcncQ6hgrQPZJCL7bRkjcYxfdW4Q8oz
KEy3GKPVyUOdD9BvdUhZSpxntanNhCXBEQ3Jnu5t7fHcaVK6nPqKeue3pFEjHMPx
ZIVN+u1NasVXtbRjKSEg3ZLeZEMK8DWfDra0/qyR0KXNXlm4vnrNUD97H2m24m0v
U9JtAMyF9oRJcvVmWy1ywT+PbLs5mLQQQgpCzOx20+LRpjKA+EoY0SnYiHyXFlj1
tJ/hP3ULeoPZoXSHMnZXs5PjGXzGDfZMs1/0Pi7A0jIBK5RH5qbgKNXTrcEVDUFc
DJlyQWG1gKKQLok6EjREO5IzoV9fu0jVIO0R+4u57cjPIBvb/8gqAHo/OyzIEqe6
CMJ7DUx3NzDn7WQ4/bINY8vvIRdIgqrbzfLvgpD8ej0nrEcISiZlenX2PAZkKKgp
yDgLbJy6L/PB1X2+4Q6IvnrzuQea3Y9gci4NbHBB8A/6OMHH6LRgiWff2R/xZwZN
It5kkfe4h8DQr33JUVTIEALQ2u+DvtT8MAhoL3P+qHSTydqzn9VEf0Vy0FIry58G
gNtbo1tKomvJurA5S0yPWQrpDU9m/sFPK3/4JVsAVKZxojAdRuzQCoai/7yYCri9
lo2Awk67UX7z4HRRoq9szHspIsetYj6vK4lzr6ZFfwyvU9OzQpeQAi6p802JF0lN
ZZTjt166GTxOkeyPKcPcQM+bVEtMItwB8Yxs0SqR/RdT9FkZGuSbwCUUTLuse0go
GJpv9o1Q/mi1i5INRTg7/WY2vvbDZSzgFSJ8lSpHt7Ina73KxQvZibdvdQvLBYJB
HVFGTuOCtG/v9whs8bmc8wTBilQVVwUpQ4F3NlaFOtSqTrB9bHImDRFtHIwGOyP6
ooHV8gA4aqNSlsUbFWTc5hjiwOnHtnFdZ9Sl7lisGRzp+q83E3ATmEFSbjCTY8D6
xeTU8paJIq45G4sxdAxDIaBnicvZyyIliU4sCFnyf1C0r2uRa8wMHdctwM+Iw8WH
3h5HVzWWxaRVpfq4YEdCd92mSUxlrKx+dfk+EefV1RmGgCcR0ZqJ99XArtZ3O+WC
kgbELVTZ1MXsng2eLhq6N6RuurmQyFzA+NcCKSjCegZVCdhwqY+C2LodYXDj+We9
NgkxYYGx81aBWl97a/r7x57jWgiyKwA2hO9AFl4j2E1xol0uDoMWIomLtQgpShOp
HjTko/SaImc4cFpKXnTmbodhWGjMxkVgyPrfnCBmODnKdUW1vQr5KWwDwGWAAPa6
os4nTJap4CXPghpoLSEmAV303XmTOVKP7mP+DJxt34sKR3kHdN8tCYTKUoyZwPNG
LpESlirPHdc5CXtmDkogV1Y6UkjrYVez0QRbdtt/3iFGJp4sirhjaNpSoNY117IP
AvWUMAxtMwq0ZROcLMPYpbesv4ZZ2B1en038BQkct0YyERXOtm2c2PhQ/eGh4WUd
J9NDvRJwLRrqQcOutdsSusPShOrYLdPJdtGhx+jsSn9kc2GY3VCoRVmaVVuKQaFY
J6dtA+p1IyET83m/NRWaNM6vmP51Xn0JfVFLLGtNYuVsZPK+F8MFGpGzWLCW5XbK
GSY86DKyv+ashvEgNJMEWW6soPKvqatlAtDLFhDAyk4EYVwIgAw+58eUVRRhYPok
Dh4m9BVUf1h4OZR0PDXUjol8ZW3bDYba9yHRvaFsqmEqHDt7IJMaqc/T+GzG6b70
LQQnj3GrUt3OV4grz6epdEU7l2wJEhuPes86KdacaIeH59lOclnk+JZV+Ii17alK
hmFUGQfP/V7vdi/i3p00nHbxsqt1k+FTULVZMa/zX7TMXtTe/K7oWDd7YbTEjcYB
CPejp2ur6OgsnkUFBCsnNA+SfOrZNHtCW0ZV4OTj53ss6uBS6LIqAi/H31zRos9q
dHDDotGxdBvQvxo3wsI5eQPDmxTNOkKe1sOyRe07Rh6+ot/HkU5z2iMqphIEhs9o
0A+Vn+KrbP6/iuxXOdU+texxeDMKRqlgwrTFNsKOP/pMNoHEghiAfGnMkd/rXqNR
w5ktKNtBiDmtn8CA5miN2/9M832mWO1c/dYysCWdzEIPy6wArEGI9rvMh/aIgeEJ
hSptEm6fas59Dcu1ph5EMy+y5RPBhQMiLMKHBoaCSq+cqPc42hXEaG8GoHQ7gLX6
Z4AbJThDundCfnd5ZXhQYMZO4QbEru71FMeNP9pIFnBeGeMu2b6rXY8haxdbipA+
QwCb3fzvuvgtU07kpxcTDcywSkZzGsivoS7gyNAJ5IcehO0E/hbA9TWzfQHMOKJ5
psKayAv2Pjks5xsXkQQxIRLHaI4QVr8fg9EWr3E2v60kp6v6rylb4JUkwRmY9uy5
1Icm1R5hAuYbzDGu+3Kl/5JTiUfK1ga+nmpTMtNqzyzkebawZ7fyE6C9O2CDkual
dYhF5BajFn1sl+NIBab7LOx1lpx+d8KNR3YdNofozHxFjpopVchpb/4074joJY0K
W/XhUeONeGqb4z9dSXg6LbuEZP+7feKXrBZpdECWNU1atk2G74Ruw1LA2LTdUqND
bvWr9Aq2Y4nYlfyq9ywhYQk6jAWZ6jjVKPgDLqUD2oThiGYPsjhALFOsCYZ0bEN2
/vLmH7QJW2jIbbDciV0uNxS7GYSJhCfgQFyvzjPKvX5d879gKVGWA544K8p6bk6F
J/rndg5q00AtsmFN1kBXbowklvkFt76LlIt1oF5OTdbEEnqNnKXdzlrM0glmvYVr
OA50ZEPehpkb0/r+O1T4I9HiCIKBpznlj7oypdD8MvpRR7NFIwCWtjUA5oEbOrfs
o3jYmYrQAVZgbJpQgE5yK3s+INSgFXK/foKml9N83Q7auflq8gx5ZUj7AYIYAzAx
0pCUcUMhKFoA4Ovepfx9NPFLODtykLyEHca2Fk8a21ZaCDynKzf7PuZVYCmsu7My
xfF0YigwY7XE/RRSzhhjD+YdBd+PhYkPSO78vrkBqxQzwfGyN636L6fGYRw1rxiS
eGIGY2U7GJLBEG1GWkCVo+uFrh2sstKRUZVByyE1BPHlsk5tZd9/5b8VVDYxux/y
ntRYV1/YnK6WK1LevmNrc/AgQFjmqiqIuDqY5Z6ZSGBJ6Sbkni/KLq6G+TZ6GfXu
sGMvZjItqZmnR0RtQsRLXxnEccwsM6PulKH6eKm7SpXEhAu/OrLjx1r+bX89plIl
K8yMYLkM5LpYNUUOGWul39NMn2QxfZAR0POoDNiriSvyifnrrKx65jVDBOVvnDQi
ugc0+eKRoiKBTo6qEAXUTZurLpPnKlPEKcu2TkRA2nCb9YW/JLbBoF8il4q9yD8L
jLawoy7Jq39IVi4zCsMa0xwgJwcIvqRBKnBgwwTT3+bct9aQnzSbisE/SJgJ2p2Q
qAGtwUue51bpZ5U8X/WTyflZiHPkujCrF/Vq6YN6dC4f/NfTB11h9zKGFj2wWQxZ
QPQ/mzSbGy3g3y3mOEka0udZl6A0EQEPs8LMUOD/Z7Tb6BfJfKVf2qdEAlJwkBAn
XXxd9A+qdk1JrdKLeHKQkjAi9blS+r/9asU/Jr2blwlIS4xmtLehDiCTjIDJQai3
7ZeWRDPi8Dn/oqbKcBMAVy4pDC7U8OHh2X79WJUTAh5xI5EvtiUr7ScAsOWvUP5J
him7yj8ekkMha6APJcLfyIAjUPTkF7/aXfsp/1Uhcu8Jr4rVA0v1n2v7IXmcX1Ul
xuo5iQ83bgBkUYK/tfa2zewMrXTZgAc6eQW9/plKnKJg1YSpnfbznOgftrK7n/V4
0OGjaCubGnQwtLl2v7WAIUXiwJd4wnyGOeyWUSeYCyObyFwuLXEMdXvYCVZnZ3eF
5WyGUcXz495RuieO2i1vo/XtgpRwH4NeFvGefuJewzJF4HtHbuO0qmsrfW3rdXL9
3xgP5a3KrME2Q/8OlF1ip2i9lxbw4rqRLWiHZyqPkmzppUxXErRP3ek+tCDidaEE
UUseO/OGkjWl7X2K+xEqcqDKgzidra0uburUpKW5KXOnupM2e2x65TzNQaHBpjQL
1sDRuWy3EYpsJqwKt5fneooUpXn5sAYs8AJWhq0AFsPadn/vSNe0gjwNQqb4SH93
kQQsDib+Bk32GJ/q+vQFpShgw1rYtFjvQcqsbY2WbOyqgyPf4vWgNSO9mcPSYz4a
BwkqKeUdQU2AXeF6TH9fU6kRH/hYL36CXzQrVEQUNx9mnIsu3J75LDrPA3OwUHb6
5I1C5Hho2kYMuHxBT3XLQcLc7CJGAeFX6eWHfWMmBLyBzo/eWhGds2HGg7m4pyCr
1sCF6G425gynCTjSltzVjfDZeB3eilSEBEBl9c7kY3VixicCn6YtMb6YQrjP33gS
fFHCtwAiyF2p1qUJcc7mVS3mbrxQguf3qC5esU8RUUhKpwwzjUYDDGSpsqmxwyCM
bV+hah+5IDde0XDsIPAiqeKoob7IICPjbuIRvf2v+3Kjc9EIOpKmJCen8q8BFIEj
yqwToK17oFZe6qFQruVtqNw+qzqxr10kHumZndzPU5cT6VaYfWwgCk78aA2CK43R
g7XD8IXeV3iLUwS80H7eAQviPB+zWE1UC7wgVjMiSMxxvAaInw9BQ8BGvtiIVBCi
4CZ9rBN7c5pSUJTwhqLSvPgqn9e/4WazE5ii9W9xJsvR6RBAIMYD+hMdzDU1lOEM
TvoVhVmdzndzM1l2mxAktc0MPamSQdQO/Lo7xJ15QWJvaF9sWeboPZT44T8Bsc/N
ZpfXu2SGLyPa9bNb5SM8KopXll+WGV2cqUh+8LSReI4K3HGO+C0ZPrCuEcp0Ut7Q
ibHECHUdr+9a3SKgHp/9lh9ksQHT8T69QU8Bza4O5MEAuFlNJgVd6/gRbWGWBxCT
9cpQyDEwO6s7A0NgSbW+DK8j4IOfyCzwjwRt7OLq34X9wUp2Jnmwl0smS4GTnO38
Y0AbQtlqmt781E3cCXigKP+97OyhyghXB/dFVjp99F6Uq9MFaNzNNhzF3Om5jKue
oV6vUCWGim4lwsunX3a+PzayxsWIiLIMJpSchf+jJMellRZvFC6Xizqg7CbwcjGJ
5wGQQJOslnsnwbbNw6ApI/4hEZaa2oxQ3gzSvJYlS9iVLvthScEZGHGKitTNVz8T
B8iDPUc0aR9FWfr2O38OiBc2djzyUxXYgaeMX7AudLcpm+S8JujwAJuOxqCbjR4/
hBfLd9lqn8kEC+U00JTqaKY4O4ITe77IQzxcb6BT0Rg2IFU07D0Fm4IZNHKsCJ5r
11wQzfD5UjmjHTu7QcCnzcZE6tlIvOBBW7NdD+BTTn72j+V9SiOm6zTxGmtlp8Ca
yCZ7qBZ09bkpH/bAlahKdonSfxHUeeegzIojFb7ByRY8KYsjEbuUUtV7tsm3zLN3
GCvCcOtEyoL/lRA9zj1jPmNLipsa5lcTYys6GGCZpFOxHNFnImPM4uctgaHFRGA9
XeiWrrwB3NJdTy7vqzXrF1tX7pgQ6PSGKrkD1kq98YM7xeQzKTTRIMsqvc5OrFI2
AwZGAyJssPm8OTFIS2+wt8DXDtGaVX/+5bMo2B0yK6laf7iuV3HyQZAcbD6C960B
KJDlUKb62/9+p9uTDdI2UKthhCD/5iJxjsfjC96PlXIGJ5hs1nb1e4MOxtRE+Kvr
yddLtymtZ5nkGcH0yi9iUlKPeprlE5qkXbvtl5nseAoTj2NAru5msSbCd711TTLY
oaUQXFGdeG2Dy1wxJpnSS93Bl+1BemJGznA4YDRAy61Q2hV8Hwwj6/Wg4NPQqbd6
zgAgCB05+0Nxsq723ZkVZ24Y2GQT+rceUh2MgWfQptzZfzcDhy0ndUJs4EqF5rwW
CF32qk0nEp5RZFGvlzcMgCb4M9zvRZt/fOo2BWxowjaSXURi4SlyvGqjrTjKn28M
/z74AdywCvAiyqFEmEmgWIMNhfno87qSQEyHa9YBwy1tOzqHm2kELG81PIW1yV7e
/cCRRQqZt9L4gSbG/zEEXjhSW4nZBrjtVZodp2rf3k43/HNCIRO7ACzJE3T9qqCY
nUFjmc8lqe8/Y8yPsNG+kVXUw/2JnVxVnWxnztUOsIhRUzpjBgGoKxP3BUNtSjyN
7hvFaYbcoXm7TOypCoXcyLH1f01Dbc+UnrucBSP0p8kLe4dMxy1zE9haD4V9Y4nE
x0u6lcE4dVI4ziI64/JBaN1ZY9o/9fk0AizCbz1I/vCJhVqIIs1pPz8Xj3/JFwgV
qf4Ynfe9s5iUErK5M053vXKgYTf4sUxqC6iSf51ZCdPrjtQqu7NuxiCWF0S1WbOK
ZwQipbyz9kEukJMNnPQ/EWEiZzkga/hi9T9CTuQWJSZ/YtPYTf0nKlMeN1z9Ff+W
9hfnqcmsKfuEP9zz1v1vURkG12Fhat9E7AigtOsn0OmUvw00bzJvUwH/qVxizDZY
acYYDrlYZqwjdMl/y+gP02d9B9rzbVIqXjm82dCvQbLFQfNKZZXqYelsro7lHzc0
a4f9U58sEU7TX7UC5pMg29Jyiag8Vnd2uG7D2JDA7AyInRXpOFA2IPI6ACMEGJLV
2+tNJifeHabI8GkF6hV4GlHBrLsyw6aBG7Kile/KmaGgtgoQDFQWnLUfKGe/xDbr
OefxhQDZUvPwOQFE7GelWvppKk+JJan3et8sSu9zem06lm7twkIx1tQ/oJ/ELZsf
tlFNXs/wS0su/3D3UcGhH9UHlDrVGeI9sVFMmAsiL9nheKPmrdSNqhfVi598Cwae
ou1mVGoFXdL9u2rkAHH3/+YrIOpFM63MCslQJEGiDgjSWDW0L2pGxNj/tVnf9xVt
/9pgm9xg4XFbbyESd+hEyHlIaUuTdecNBucfNG08gRzy1GjynHbWuCkLZts/GnwS
9sid8DLftiV6hAIN5jt5RVJEHeFlRvOwaZ0g24ALcZ+kIVBI+LotGwKHmFQoOtC4
pgNMZJb4TVGE1cJBoGea2aeJlkACNkNC6/G0pRqdG7YppohZLdwZ/4lcKkMinuwz
MnkdWhhWY5sqW0IMG/5R5hb+ONHUTR9YryjI6KfUxc5jBhqRZ4kIuM64VWxj63RX
Tj4ubd7OxSwotnUdn2qs0ygk/7RFbEjaBa6bDDlRKCnib99bHA5e0nI3ly+7PWN6
n+ZQGp0DZ57dl/b/XR/s3P1YQIWHgoFiNSFH9I37PI7lXq/R5rLa8f3qLGeKCdto
BUQvDrwmuTCXjHMLtYETAvWexdhgRmh9gf9kYHoubRBdY81u4l6+Miy6+oPwCyfL
9j3V2weBxeA3DbY+wWQVal9AL8IAOm05Hu59ZZG9dpiywLPwSRbqunhWlLhIOJLy
NkG/SzJOUeRzNCyP5JHUMb2DhH8yhcRF9iNQFbHHkmgXRXCkG32v62sRR19gOBrU
gRf+ha818RAjKCL0YE6XzJYYkvdZwgKdHbPzukAogMzfIuoBkPwop1nWNPMIk5HF
bwYoUhu5mCv0s0cD3XrLNQ6epxz4Qy/55iw6/QS2EVr0OwkxP1f1rXhxzabzPa/y
Z1dTy/txp8Hcmgl5sd0HQ34Q2Jpfkxzo/nM0BlhPtvT17oJcL4xVmLxpE0E0AS0j
ThcxZkURnFLSoCVXlcTvahQh2z0TAkWRdcYG06wHmtbzNM/bC0Uhzdou5xeoIex+
kPar/hcci50fNc27aiPg7+I+7ywX2jpm6c3gAksZMficIlrEa+kYJzm2hSLNU9oH
axt7yJim53zwQnRdhzjDDxjPJpb4lfR3TButNN1rMxk2t5IJa3a4Zp1WzWhys9lB
jiSo08q7PvLzi+iS5WurU0AM0ti2XONxRszQW8bP4DrjYUikWZMvq2KhvZ0d7zHj
pPs9CLbJXmbvBvP1dov/dDiA9BCUOAAt7yqdWJ5PEpfnWPwNW6gN/CQZvtkw1Azw
Tjs770XL48RZ1/BM0LameDJF5776EYfe6IwpQcxN4uGIr5l1eISv543ohyp//Dax
ys6TKaTS8h8YeK0KqwE9smwHv/G+lCG5WDDivrNxo0yDWouxFD1Jq8EaPwLDGNc/
Ja41Z2p3YoHRVt/DaonwpNWU12UVarI1p6PdcCPc4qtWVZd1/zeFLOMfopRL3h0u
dwV9+h5zhoZOoCg/bDPRMy82GYCIsgMlBNYiNNcfWYLiZPnYMwTnKtHQ8k0uKL0Z
sdzf8iSk5hlz0RkRK9FQwiiz37yNsbvwyXZa0297wXSp1g19r0iX/4i4kN/g+jJ9
cztvSeD3OjzBd7IlsH+1koAK9ZfdczGsE0s/M0Y3NUNkF2CxL9i4h+wRSwhF1+/n
gQxDt/Lx4JlEAkDK/TEG7wu/8eqKGcEs5WukguZuoqRJrEwatKhfhx3ihqqG2N6N
cAQMPykU7eH63Ypgi8Vdrc9ZTpm0ZQpYFdXsFNPG3k1301JXtmktxuRI6NxnjIU/
VMo8Wupk0dHbf+01a+Q3AmWHqd6HxIkCPcO0WkdCdeQLlWQQLz+ObEVn0DTh2fNw
cJi9BOtRO5/DgRg4wM+HAIFzf/1/i7cWptD8rQ7lmxIaH+ZD2qGXMIim947pilNS
rbpcUPvaIrxhBwJwH0XusoyfWO1KFjFHPmM5fx2OV7I4uYX4m6YF4LNLBtGaoxR7
9HyeWwUd8+fkAPHKpxl5QQfQlDpEWMtLI4/xL3Hki3KkIUdIuXtk1Wd5Efmqx35S
HIStP3UD/RC5Op65rdcF/za6Pozw77tQVyxIyegfohY1Fz/B72B/MzLydwP5aKIE
jdyT95UmOrGNkY29rNuWw5PihkiFknrBvgIGaDnum2qQjPIU5kXwtWEqccg7deAv
92Xe1/1UPGdm3aiWIgXQcLfGlU1HGRVbg4nbryf4twltw1p8dUhUULVgno2pnpsA
Mljgy9K/k9fW1la0ioFxFbVI9woIWHgoRBR0s6Pf8QHiQEeSmzEvXftOXXh0lo1X
MIBFhOee1ufWsaI1kGuSMsCHZwqpmZIvqo88ubKlj/INVmrJpJZSYaoJuEg+uCWE
m+GD3wfnWUJ3eb7dCs0AHZabSTQlwN2BpBqEcJgbYWcbVATDBLbiiduqI2clNASR
uz/spShw1V3K8CTZndB7NHCycDgz66Mh0v755sidQqGKUbX3ggZCQxQEWEUsRYTC
QhHxHweAu7EaGqVMiaF74b3+DDtlxsXZlad6AOdFTvx0L292e7gmyppDX2AIGBQj
4F/p1ED6yZQoSOdPzPj7AdI0Z0vojX2ffxdy8uqo3DnaaBL1nYiLm1VRh226rCVX
C5Q9XkID4fyoEgHL1TK63cvMxLFVHeWlJ47mWqp0ngSdftwpFiveH8YnUh/zG4IW
iYeWejD27W3rP+KCQCHg70JYqX4dtKDErVO5X0KLGHXIYVCuazLb4Hej6bQZQour
SMt0jhmFT5Njzav1zOJSFbHyzAkpS6IJDka4/xMcqNUYmRJEVL3f9c97kazt3i8D
+yswvsDsmHMq66j7E+ZVYVmqmO+15GwNosuw8O+YLAIshh6TYJLUByuCUGXNRxXN
C/tDGR1UEez+a0tG715TLkDJJLCBVhzZexZThB7VuyLK55AODwDirdUWJys8p+6X
ayV6KWK2NC01P4BhgBOzVx64wA8oQ0+jauxWK9ts92g6a7DmyyH1SlcGikHC1UME
XgfPFIi4Xz9VWW9lGa0Q+B/dM+rxG242/P7hgCdNfZDP0aAZvIqEnaavCa5cZOCj
gKQi9gkAzbt2F9ViYhHoPTeJ6TH5e3E4PqT5MM1i+2K/Vbmb16MprV2voUEf9OJh
bOCyXrSaJ4i0JyzvJXIXK1a38arIHP8yrg/Cq6S9Uc92mkISUI1u9Y/PPI0uSZTR
AlYS6fk508xcPIIye9XIM9qI82b7ai2komOGzjfCEh9VVRGFHkr0XBDAUqY/Vyse
7THJ3JJ9su0UJkPgsuJPKedqNgMlLova1JJrYJYkcm/t0yjh+MHBNRNCABttrk18
GMnf7qbyAzqmrdvA3P5dPWhPtjFjPm3C9oJBfKss6smPu067Nql/W/+HfR3YIH7C
N2JC7whmZrvz+KjMGYC5TU3/nUtjl6l3dhpOCxI3/xuYszUu9vJWZPmCALvz5LRt
4LxZFJ2OBFi5g2rcvhI97ZfJ+C4rN1/ZP8gH4hqrDIVLqGc4Rxqorp7KpE30ByhF
Q1I9zgn4IIWWmk7D2Qngt8Yfxo7ZlsJixumPynKXlnRiKLxMHfIXIXv77t5NlyLf
PP0RCeiMi596ZPsBiYEspc6AsYmHonEyCXDooYCmMYHB/If3z/V/q4lNtV7eg18j
L2sgK/vU0QYlDmPouIS5GffQooYRxU3/N32V7uPdQWQELGfhS2nf4D6K0RAss3tp
/e9YwrN1hVwoD+ZD6Lzx42FCrPTTOX+BND88I2abCE890CzlT45Jg7W4wcmSOWvB
AV+P7ZF2RPi3cJBphF5PpL5psxV8Si6Eq0JYh0Ir/oaDesY66vk8IqwEUZSpdSSE
s5I2b5bMAjq/h9KhkzYfIYi0V8aE8yfAV5NOJj+5wPWaL9j7Kh3ptm0yBbAFcXKh
jEFRkAPHlzbnsvckQm+RfObYZT31Tmof9HARiZedtZwZSQ7W+UiVGXA4sBLry5ey
dznl9snZHes221+/3a6lYffGqWloHbQDe5JVocQpTsw0tyqhya4/tfXd+PxJ6LSN
FDtZv7SST2cBrzUXZIRDHxYm3JtxIQX8Ynt7HoH0QfMNOE3oqF/xcW9VPlrChxgh
WbVjvHGOuCRRGzvOx3kKPyD1ibuPlVcjXP7MqxM/BAfbU5/u7kLiQCXe76KSfwH1
3jBzMFcT+XQWFksJ7vN//nnZDPScxVTRbcm3jrNmaMhPXZG73SJpWgbQ7i4tj4V5
RL1eloOqLxjMUuE3jj1IETKCVMAQ4y3jxofieHGMUU198AYQo6y4uXMneArpQAoz
rFNZNqkItJKg7qsBvWIyA8nh0HM/soUBfjRoHD/LApvT6id6bh7wNBdjK/IxjCi3
pkZIYTBe5Xg7v45Om7x9hZLv1SWH6aMCU1E+vxGFqxwXnF98X2H3g1n2FFpk9rCm
LjDtllWahi2q+WwkSRvgDO0Kbwcnf0ADzlJraFS/gYIg3bcnsVGcVWhzTm8Q87dv
ghw+LWNM0ZtLaDjnUHtHfcIHN360L6HuCC2DYT4zQfjCjOZt2G1hBI0NHugSXWZX
52wTgbV2s6kwK4sb/TBhwsJlRqr12l4EWV1Voc5UKyGEQRGGrYm3/GJYVSw2/m2m
f5acJfSfCP78ZWq5AyB2ep+0k8A6/Y12Q6MzFjAKgGL5S9L6ChmYOFw7Nr8B08hE
Lfossah3r7irkae0/2twG/eP6i+Xb1uucZAPfbIfl3CWflzDtQLv3JzQX6s6cA+X
4t8Oc4yIGaBfpwgAv1QLHsRLGFQTM1Q5MiSafyAbsqf+IO7aE4HHvF0k1Qio3PQD
msBmvd8/XcgYNcq4wYycFkvJdVDJPtpE9NOZYcg1UzQeLkwIs9HSJMzcoqtYdNO9
Nn54AWTJsDYX4Lty0GVhgqbVlmeAGLRfCKHS0P68X84+K4qjICKupeed3xZqpWAO
wCOfbbzlRWMSw0wAMjZ0fwYINVssIzSeyb1Jf9Xr4baW2+UzdVf40pQS/8Sy6faJ
gs65LQ4A4sZlF3cqWS8GEz4D+WSKaBZOcQ1o6ramIwj/atQpuwRjOI0BTL8aWVzL
1MXb0gzJ3XFidUZ17aGm575y0PinH4jRhlOB/lvOWd0sMMONw674ENNaMM3RcxqZ
kvKC4mxGmQgnPUpGNR8rmVU4dLDb/DpxAZLlkimr32/vzOnkIOqJjbZVXT/1pdxf
X5Z0r3SRTTUReISUNV+Sc2nYZBIAS/Dlco+32CVnc+l1U1FTOyDRo6rwZZgjJm7w
6Rflyss7ShY1KdOOgFhIzVBe0bQ/PEeNsh7lLG5iqIHWTsqX5oT2T1lrBnWgKHcI
iv/IBnfFwDClRFohIZ4YAqfQzleZ9JWrxOYkYd+fNlLFVR7qJ0kP3Wubt3osXhMU
KQXKFf4refkvddfgHxEKOGT3ft5+l5Ub/pRCfg8cbD/9C3++E19fNV4N6JZKT0zk
AEWSMxYIINexCqIVjuUAvRpOWhq5mGbn1TG2UDzzyQQWYzWkvkwv/xyaB2n+Yw0P
wtQbGceBV6iFXHiXW8FcEI5z+kRiLm0GsrRUw3Brp8HFqEqeg2l5BJDdnwNJgdBe
5V7a9sIMP3nPOcAdyoEW5c+Rk7U5naFamIfHlcdYlKF8CDN/1T5R9nzg/sT97NNj
rj1y9UDyv2ZwIxro/NegvFQsIAbHP6smocEJHlQ0ojWDQ+/OarKSqc18cxVQYrU9
1uVgMsWn+QFeANhH0oUa2uRIBUukNl2CB0Xk0gLI8BAd0aOY2F+fUrmvr1Z148HB
vgbYufKE5HGttnqCv1uSAtYTCoxomXBA6ynCMbjswBZhlGR+PeWRDX3YH3uzJFaY
6dTjNxR/d5IH5l9MOjqqNEiMcnSRVw0WWg/U/auAiyjgoDPKoJ51QXjhsXA62bYL
4woOdIbO/9DsTrQTjl8VymJhXLtrPOn3dPbwI01qJ928G1Eqe3Tqk7JaAB3H3YB2
MyOJfRgZ2ZxcQZfIssQIcwBxux86QOcOze5jSGDpFkv7eDuwI+JNMVdArWxr8BHC
8NNEQhrA9v70dCKPuSm088voo0iHMGN6ZuoT1366FB+JupjwAL2KhLOUh9HWxBDC
w04dDxxz1QjA8O5t4tS0CeGvQuWzKKJrUvRxuSLDDRzHMdy34MJt+Lthwft0NOJR
zUixnhhFT/z/KFq+pakI/XntiDGeUpnegy/mwzF2wTStWePmWOPdv/NN4jcFMaIY
PNUfh7yNCT2TcuQDgtMvCaKjXnXDP1T9iQG4fzzDJWJ7cvRBjyXoGNkUN8XV2Bg4
ukmWDjpKCgp607tgPOIS3C2PgUeCvGvDfCSikI6R63rAfJjKTUDjSd1RNeLpucry
Np8xT7d2owWgeCiDtq0mADGKd8h7DE92vK1qnrGwQBLLiZCdjb2cSTNwMqrpH8dz
Zt8OQlNYuvlz6pKErXSzEcFL6vP6qtUos53ZwEkR3/pwtvVCEsjZKmZibaacceob
ljfoePcMpDlmWAEkbJTuA4wZPZlwbF00s3rS+AKrlEqtEGLPd3B5OKizn9wHSPKu
QkTLq7z3HgJSHVj4kawgBbKbTfzB8YJCl+XUErgNLTecdmyGjXzDdcRlvUpSsETN
mpiF2+eSrm0sDP1IiU7Q0x2eo1xwMLvsQybtOJDLr3716H+l9KokjCi3TNCPHuXJ
RXYtpu2hmphEWUKx6papRvk8PgzMfxo263i5+LmnZtI1icp6Jf+U7sXQ8t/on01K
BLsYVDYpPdzFMp3kd8f4RtWHZFBT7gy8vAvmSCEWqVgNLs/08UIVzsT+bqfu44xw
reWwZxNxEK2wJ97yPiFzAUZtgIPEZINfzs4XjUUUXYdcS0tX2llpBKhExcMKbqi6
l+oIVXiD0eBeqIgHJTK05Foz5xh2B5n/0Zaki+FbaoKFMmN36RMCj17vJwQc9dqo
I3kyslbUeKO4msaYCsPbQ6qLWJmsCrLBj0fxLovdPh2DRLU4Ec70y+TejQSODs4x
FGadiEI4ry2cudhWUv6BSZ0j5E/ogJNIa7UdGvHtMVKsZK/JD4lpaE/JMi5v7HJl
fV+vaUpHq4Gn739NEqBHYAc0nQo89r4XOXknM6mFTkfrjL2PIMdpDC/EIPYLasdt
Qt0drYnMRbUyX59H2glG0eD4aBVo/sHiDpQgnYRuOTKm47PtvW8fHHacgvz5iEDF
cFTFROPjQI6ayQA5v3OWKTD3LosS0fO9DxHoaTq5JqJbp6LjFDKIFz1C6M1cEG7v
bmouiEbiuliwn8kmju4PVCLzRvbkUmVKFNNW7A3k2t17PJL0o+8+e7Cm77Dit9iR
2iZdlT8aK4JTp5ZavxZJKyVKjNvTYJ/KqsKT0VNLcz8I3zYWCaGfPvauzsrv5bC1
S64+O4gDGjrZLGBJsCJ8GKU5sJD7DYc+UMlVTcC/uW7dtWt1Md9xpMuZEe9OFugo
1XgxX+lWscpPTirRQZxYRpHqmumLeTsCjjBuifmxhnCxZZZ1KSGv9sLm/Ay8mCEG
At3agDrqNcq8wB9VEqNVftpDD2kj9ksCZ08FwAT1YEO5jJw6u1SSh2Ssh2fyooAf
V67Emmj4FGs/QoKaBAVhexj24orTsDPQzR6Vz2Od728u9hHZQJ1xgj2Cqr6J5BK6
+vUAaiM3rQo9OkunBHMm6eJkf6rIlWt0XnMsks8BB1u+yD8a4Lc/mkNcYvscS3Pw
jLGOA/wxHoKedCzNQINvK7WlIQm5d+EnZG36aTn3q2VtgZm1BVD9gJrNZb2V/GOW
x3cBLX30++8fBF/9kBKaJqzAPMdkgMjo2EQKUqxg1c4ieVuQu9oPuGRsA5VhxsDQ
COPXxjIOvJ5DRIgtTUpRwQZXbKxo0raF/BnxUahMv36cGMkWLWzB8WQeqqlfux+i
4TwlqhoimLTdUo2kwYiTVxSi7N4XIW/lg2WDsziRegZvOv7eOxzc3MvPaG5upX6T
+LXTfwYurLWd1O3z09ueyJfhxENIZnagSkzyUWW8uuiirBL9qkI+OVBQDhEmC9cn
JkFs97tA+X06WY7rjt4H8xy32ddWfo3cQ1+eaW38hHpWoHh7ccFHv6M+3Sf654GT
KEL2yazalWLWvK9c8oML9RCh+V1/8Q/sl8yzOKWui6dGn+/d1XYs7evxF4yWJtod
C+tw6f3vQ3fQWXbMK/4sSuyshkYY0IR2bY9/0GyMSyk3uqioUFV/DvuZCSNNXjay
yx9f7fzbXv7kDQmFBmOFjYNPnz++kFKCwwog1dpxwiiuKYM05oR0XRPZUAd7OdDW
cYBprHHtBokgQna7PC4yIBh59QflEyb/8s0K99LbL4r3sbM/M+Bdn2OMD/CIfGgx
Cfv8Xu2xOb2PRt+9r5/+gpeHBNPTc8/Ku1C4x5R6n05fsBBLEMMPe5igVkj2iwZh
ew3xRlSuGP7aN4AYTps1Kj8WYx+aXuEzOAJqy76wWCKiWb3RN+DdgswxFI7Y+f3E
UrCLYpdQBnlicXkCOqEbnCtGOIUDo9ed9XGWbo5unVTq862VXXEzmIsI6ut4o0Wy
brAMWHDcthO/Kmrfi4FaoGQEUY0EIbSaFAIQvsl5c6iqLADamMEGdZ2JxNKBG/LK
Sp9mA5A8AaPKeOmvUtj5EFuIFpUtfgR+cAJurb7AlvcY16OOolLnvlMaaO2Vmd/C
RYiFdBUd0R7GNNLB88Z+hdByXuLT9yoO336GDwkATd38MWqEIWsJcSa6DORqJZCm
tTapxCHr3qGJgJWA3ZFk8rz9dH8V3dMdFA5hRf4TGwxIDmu+B73PR5UebB9pWWVP
S90lREQcTTHH8imB5o7/vH/hEgX/qaR1hySsS6iKQaZKirg90WB8kQWYhRU0ceUA
BGyHOXLvucrtHH3A0VwRcwwHe7CW8ZmQM3s8b0A0mJc7NuLkWd2JlOTRmE0Dq1/+
pHGUOT0bvxS5QdOKSUkfYui5JMh+psvisxCPu/Mz5Mmk3rMj0UkfyGhYPtQJ2ASB
7Geevaei/OpMJlLdfpNm9KiUUWc7F/Ddg/EDNcbo9zhOk9sLtrPFlUv0Z0zWlwmp
lJ0aYtZol7AeVoUWWrJsxEaigBj8tkQe8jgnnXuZLvjCgidrbsJZ6Hs7M2IfLEwA
fxrsbNr+6j+xi6Vs2OIrCHMPpzN891tyZuTCLTxGqHNuEvI6+PIMhaGuRphtzfy2
53zRR11AxAPVdSvGx/e0Er/DogJgSj6GMA96AuVJm9iXxBAl66OSBsHr257MojaZ
F4BFyNQRjYMzFTpSiWrljEfy3hrhZ2aEBwmS6ZA56enA5voRBgRmDdgrGGbRtK9T
/QOfm3Kd+GXfeLxSA2YazxHdmUNs5GvAC8xVUWwJGsgDZo2W9bb00VgmtiIGqv9F
GR25bVsBcaq2FpaB1FrTJhqAdAzcAejzHpkzS1rCXBNTdmHi5SniVW1gHQ6bXnap
6Gy3ZpogeLFmBBJubN6eOCeClpAIZ5xWhE2gpaVtLhzIL8G1+mUqAvdQ3S5cH0rB
AKbkrRJer/3YDGV1SFK+L1sVYS5X6o38uJB9th9Ohhh3bkvdp+WGxHZ/P9QumEDm
fx3THlD0p8lgUoJkDnI4u4YBR2qv+gqJ7utR09ZBYOzSy48DcxHghx6KjgamrcAp
uudlTFD0Yxbn48iDmE0ew9+24OLTF6BDLUqj3r5C9KjjneqxSNclH6oYlxyoAu+4
1JVwqSyJRePAiIaujDJhS1Y5bNOT5DqrnqeHWG4vKxQ9bRbavHjc9MZZFkJIHHkl
3kIdbvdYISG7N03LErIIVvb9ZhwfBJ86Xt7XYkuspnI5jKwUTCr32XWqNkosJZsk
qXHlJ63Dwfs5DSdwRbPRDGfaenLZCtgtD4/hK11AcsMA/xeKKkKVKzgSRSxjgs1i
5d5csr+OYNo4xBR3UUtw0VzAa/xGRQ66ehyHE0Cy6uKb0/+SYLA5CSBbyO4Hq1yP
cGu9JChWqPONUFO6nOSO9boDwPkCptITF8AdxU3W9BSbuLU4UqYYe75MclQ6USO6
vwK4pJ9KSvF0/JZvOyPxdqsbiSnUdRMWG4p445wt/tkUnmCah8BT4Qf+JvzhhUEH
yfPPneFsEFyU14K57gfyxyGBgCSdeu0P+2RT/H1C2xDlRFGCv+lbKWcHkimZ1pPA
LBc+nnjsU866YHS75wBOJHOp2uLdf/7swsR48Jhxkz5sY+Pr8grXW/qz4H2+GI03
Z7e44ZHXYJPoh9K5Hf78r63cPO5Ci+/8I6WkeCGMs84snCzxMGwlxvmxh9PQdKh7
0t7ikB2NQJdTgTT79tbrV9k9Vm1fER3hMIRYAbCkGCdgpAxZY/AQxCijdI2n6UBX
2EUX3lCmRliFpWV+7Jtdf/qrFRvoPB5i41TIcTtIJ3k9IFtbqNweBsiulGqnQEgE
+myylkTjyXT6uevojWzzjN1Z4wZAFudG5ttb5xgIpINGwUl2gpZs4d+J7gwVEz7h
LbbztRAVkmW5KNM116dUDgLe4eNGCixXHWxY12RJWIuL99ZiBncJquNmOGn1PnIi
+emdJDmvrrUkPjIu0zGcsjWdDJ4KKSAcRnq9CZWuZkc35novCc5tJ7mkExAyVUHg
ghLXyEjtcMi6Zzp/d+AhOhSVLMq96Gejj5nl2JzvCSnNYbrfuVDyCd0CMFZ9Tnvo
QBwFxNhoxCG+marCIYrrYqtZE3GjUiGynpndc192d594Jk1UYXFbou9Pmo/IWL9N
8/MdOLFIw33fBhvuss6+StAu4f+xjKVGs5xY19Kr16FBOJiHgmpUe5QRht3Y9aQG
/YzXIZ6sasFAdsAB6J6E5UlGkyGu2acA9CKXKiHsMM4DHALkj1KslMSlUEIoVIvw
iSC7AmLjpAAZkU9f5ojAOAAhh5fsA7/qikCbyEHWgtCzSkY7T0DTGaVb41rBkq62
b+F+wWchRg6U6rYIEOLtqXXJScDm1EQ19EoYk6nXNwB6eqWzPe+NqxNR45/hOzyl
mik6G3tH4qDUCiMilxkSqFVnAspUEdbndI9DTzViXIC+bShV3h3K7PUAHYCgCbWn
qhxBhSZh7SLpK8ImHzHtRUO4NmMCL24y4CTR1SOT28Yp5LLxK9p3VPz5U+JlbJBe
RFkj7dOPabpG7kjSVKtJ8u9YPSgkayLhFsMTnbNNU7hBDFMVMJliGjdEzDzla6i9
ffSUDlI10BXdzG2EJN+HpoK8NTb8X1YvQaPyup823l+0Qanfg8lnf4phvTgOJlUC
K4sLOcFGVF+Nq48md5rVEOq3fNwO3C+XuEaiPqdjutABra7PYLFBGV+FFkjVXDxW
4f570GCPQbmkiFAWOGGwCDKJvhwi2Ih6nEfjIHPHqYxlTL5SKpWGF0XG4W/bbAGT
eu0iX/eiOxTViZmcx5YvkR0eg/bmV1xPnk6oLloIdqpGh4vUtzpqaESxfAvaz7r1
taMRt5BLvJ88mLYHYhcPJfJgh5E9fVwRe0/KzbBzV5seWE3qyIKZRK8rNTviq0wR
0akgv74u0+558Iiu39R3fXnarrDCithZBqhWFtUWeW0INvU9h+tOjfRmgSV63kDs
JOX0WDdn7TIgoSi5ChAJAMsgvct0XACAQW4M+ZAUug0f12I00RatmX6fc7AF+fSa
ybeUy6D1zDVHvwgj8FAC/aBZcwNs7v5RMoCaaLrSAlLRt8TwglA67JoCdHfcgVGK
hdqkMSW42gv9kLQpswOoRPWXmMFM7tCbAfNMcB+tfFOeH1eV48KdNnDsdaMw+33O
MJN7XWbN7cbXgCadH5fPKdkTSmWm1/vsUW8pmRMMtge0vc71PIH61JZfy/owwFQQ
1lCFngGgV7o0kkMyUy01atwLPNLy0v0RdxGkw5c3bV9+QweEinsKFArIBYIJAgiC
LYLYOEp/ANDJbW9Gl4BDeLbD+Ytb3aj7SYRxqC2CWORFzS83m315Y5n5/oPbFPOU
FBhE4bAOfJuQo6GEyEcGgrwl7tezAWsT1p9z9mANP+j9JnFed5/2CQUeNp9QHgD+
A6M8LEdcOPdmvsQg1n/aFiU02QeM0tmi9ccOGa4cs3TpezTqeBcInjsFuhZ6gC3T
ZmdyWST2MB2vuyZ3l/zroYTv0QDiUMK8ODML2S/oXSr2MG6QhJQjPp35U3GnBF3w
Qx6Dbouwr11H9kh57WChodhzI/lmG87Dx4W9dvE8iReLlmQiEEaLOBBy+tRT6xjM
QnJEHFrrO+bqRNAr4shvbj+glazPLTy6+n/tVTggeUrYCfxjrn20iljs5JW2z45R
SpvtWQIPor2J2oejOOLLi5DD1q8pmCsm/qniUF0TgLJH8ID7zPMbwePbvwE+I1ga
Rz9lVclDD33HF/s6HGuaZz+m+ExwAi3DsTu4YuDzWK2ObhzIhK5KjEsebMJ0oW6R
LpQrmiHhX2IaFos7z7aBIZzA9+6jT70hdZ8PAPSPM1T/JsF+HDD1mOCbhdJb1p3W
JlIu8zRvA+RKNTYxDIH80uZEpR3IzHhdv2e7bhHFrScGQrWx41zkS66tDx3TWZKK
YsFtkwKZCpEopPo/YbVwqq8Lwuo3jTsr0xXnjMoGqsf8rxUMtERBizwbad+a+PCa
gD91sW5ehxoDqRN3gr7GBto+WDTkyCQwWq8ByRrcSlHNMsqSxNtGgMhNvSSDFKYQ
qeMMSJ03CarN2nLh7Z9OTcDysYoPX1RJiV1qMAtI6YnVVqoZ2xr7eEkECHgcW+Qh
/xGSSGzimjKNg5CHPOcBK0rK4QI3sPb3PtbMWkW/nWXXTNLlOISjI3+wy0IDeXMj
pdw6V4nty/KWug/1/oNMwLLGDLGFn+ffV8vNe0tdZ2hVQep+vyB0qIpRSFxLk76t
FvzeZWdWOvS0LnAwNGx6u4/siUGJ09TaO01HzVKSwRq4kSdmo0XNTtdU+8tdCaPW
vwN+ApwubooxTS9gpK2yH1WrGHqzVNZF0rA8ImJR81cbNKWcZF/kJWRbDYdiHnn2
oVFFlUy70Vfy4vVIOlMBVfaXzoc5K9p7nrdN2IOqlKAkYKg9xh0NHoVSQlMevrls
8QozdXCUhKytvKGzJ3Iw59YfiORUHmOcM+Fi5f1DrZMdzKuO862RJxrWWhFge7Zl
UfUsOSLXGpHxgyIx4HwpKKsA9IrBKUx2eUUIyE2qV3EBl5Shyd8pMUW6X62l1efm
hZ+7fS3wUgZd+twG3fN6Di9NsjADqh7r5TNAyolKTTj8Rd4N6EIcyxJ/wsMtZiwQ
EqPVhHbxtfZ2Qa7VNrr+b46OGk4qP+iQXtSgD8HmhnI1eWxFyozCIcEpzvxLycPv
b2vFuUVl471QWE6YnLdH/3EBrTNg8KJKNcWxl2eM7SMlxSX0hdOz/LA8pRz1dIKi
hDIDXEVfnZIVeW339+QxkThTDt1QBz12hujGNNMy3naiU+ShAP6aZFhZNKJ/Wzrx
mfrrUFH1ImnCbJNYbexEyDLG8kRcr0Y0ygDxVyEfvntUQu2vZrAktIKP65+u9ZmH
OsGL7qjx8flMak+ILdcNLaWgbFl3hOSfESSCwI6fTEppHJ0xANdsNny+Aa3tpVeT
i5ckpZXVffuwgrWXhLzGghkvLghKPvgj0S66RZQ9lBIt+TcIU8eAsFlXCRdQBstc
WJh26U3q8ZNmwLycFQ1lroCb7gLp22L9vlTzL3NjI2bwZWesp2k0+WCiy5FEpDiZ
kE5hGGSP4enhvBXWkovkEB595WPGWUUaTg/KEgTtpGFByfyjoM5PNCJeo8ivyvuY
KyoVpH+Eg71JUcWbjy/mtcIZUv5ZkZ2/dJcoroTuE+x7bTllrPM65DI/dKrvTXqT
Q9MuFN9voCQC40DNnKKTBsg2/WmCR2wdnBKGheB90V6QOhdF2Y45Iym9gbT+ijBj
Wtjd4sP5uP+0KEmTExZuIY5J3U5jPW0pZ16ysrpZ0eMvI7EeRc3qRKyAkmRVv9y7
Ce4dAR7X2oQrxz2kgaEIrTAUkjzjG9wQlH5SWQjI21wo3+suRAbR5iFnde3cznao
JN5+kps7BngTgA4rvbHPOd2thWqM/0Dp19IxzGAeXDeYHIzFRYvyNbLTjrQQLB/g
3rAa+Om5FXmNUTfpKIKEX8XbAYX5mhmbByEndukZaCbHmAS67vNZ7pSwck20PmDi
+pFuQ6RT0K060Hyo091ShDnI7qzvNzuIV3iGwtYo88jtH6CbqyBmprou+Jm3XqP4
Y06gVKZDWx+zayF6F3RDKXvTKK4FfUP7sVwQR13EMwNWR/xw7cqfwMEQj//YxbOA
kSTxcMdAepAZ82TW00PuN5+OCK3Ami6UfM8kOee+b1tFqm5vNgjY35RdGPCqB7Jb
Gyiady0oUb6ip7AZF6NT+B+0HyCmXl8C4TJ+de64b4NxArIVEXr4W96JbfyPbs+I
3mDyfDlCKvB0Pqliaqd6Sgsti8nTwc/pDPrRpMebkD8ckqVywv2npy4WvSQpvn18
dpiz6ZppqjWeDDD8G+TdX/y0SvCCFIChk8djYq9GuYHZCY1No8hLLCJT1AzIyR89
Xl1LwF154EpmdCkf+ebPQlcMPa3UGw0FPRWeLH+dhqwtFbZYO/v7DxRerOvQX1iH
J/F0Ijl/8OR4pivBNmICq9JW59gZIELf5yO/Z8BbZqZMLken/aUAOLVAod4coyvz
1FPjFg7A9B05rP1p4k+zJh8wr1pPcS907m4iA6r6iEl31uXiOEw9CoHPxBpqFqLb
mLv/01zjn0EPTrVDpmKWpbllRL9za5dFqex01I368xIqLVFlPrQ6O1hSzuBdyxT7
Kb3MF1up2/FJXpLQN6oy/W1l46sOtrNFeruop/lkCMFXNlIdEFVAOSPj1BsZkhXn
vCoeRABn1UR9O5MFcxRIEcCD26xvjaY6FEnQFUTHp4RjViEyrOUWev/x7qBZy1qo
FwM9LspC0Ri/gf8YX44neKR8GVuMtcvwCALFLPlsqo3GA0CfPPD/JgGgsjt7Qb54
TPBxCXw+xJVG48aD3vKG5jP8o71wehCRuMfteJdCGgmnAXH+g19U8WnGf0QaMgXK
qm16CAgdS3wEyO56+v9LGfIOludrReu8AA/sFiU4WTkNlKhgivEQNeqEkxMHy5X8
knaBCFRUoNceyjFAALMND6/mupXP8FyqRUclwD6Ni8QNgzAS6tdG0dBZpGQgGy/V
3jjPGBL8LIVpu+1dW5d4x+ciaHTutTt0klSws9UBXqF1UB7BZbi0/43ztajjWPgW
rzSwq2NXmIul909Qrz6wws0sC3ee8k5fV5vEyBHedIWWhxrFNWmFHY9yxtfEx9xJ
fDhuyURU5yg5RTyuKE1JtHF1sx/GTQX/0be6tGd9vuT3Xu311WIQRxAD9D1ntfMf
V+WiMly1AyqrQZLm2iuihY/Gd3qU44sN+FZNcmstQRKhcQil9Vb1X0CgB3WUcijr
Jbw9TwLhT6v0D2nWt98MD6xEXD0IbK494WQqLL01NRXtCGzyyOiZGrNhoucNyCbA
H/m4NsZa9WapYjdDpxeSnulzF72vm0fw1niOdJUzjoc07rl47RANkCwSzleamjum
a5d5e0485yzzbILuBROJZ7rAMW2WIFTy1rPBcVkrfoNgOmN0fCRiyuN/BjOrPtBs
IrrYJ8UKItfdIoHBpA/SfnWa1Rdsx7tldzqYfKeEcktfYlc3xVlEBpKZTRsK/+3v
wP7fokh/CtmtkPVoT55b/TjiYhfQx1wQDhG0C6r3lb/OLo+i8EwUX40y+JUjoRfQ
SYZ6jfQ0ppK2kknNWkQf4L2NySsqJ/XYIkPFgn+U6xGPCFhzkWZ8cfPtGXETUfhG
r40XJ4Mcz/ba6FvGEEhhuuULIyAyrFMuGwYAr34roQOMdRwPAif646IMDS7Z7Rv8
ZnN8Ir7j0kAnwWt8+0EiGRMBDNfrCVzYBG3nteAfUUjUXqml7+xrjcBVQUrasfRl
3ft1dSvhujTMel3B8kHLu21kyXDZsUBmlfD0c19veLjZh+G3dt2PQhMzbXG9hF0B
TSprO+5skyo5OCtBXi5ZeQN/ZLI1577q1+C+8i5mLe6RS1BPZ+tIHLJmZ2sTT4Mu
MXrdnMr2MxqYuRqJ+fBsILmc1itLyP1L+9MSYnxa23ttyX50HNHm9K3Nz362U7u8
EX72FHaPON9ouEzR/1Ri9LIdhEg8s7jry9HyJkxvMxnXE/OJ6LvkHdvNw8eMjKet
3FNwpvX+cGcNChYpdOrPPiPbXU+7g7K778UnUJKNm3h2WZdM7g31m8qJQuz6aR8n
HLlJ8JHV2/MayyeRFQBBbT8Q2fUD2cHYLIc62n31AHnPsRAGD55YdTtn2EgTMF48
SqmKVhzMpF1vraovsic7kC3Sk950RP9rEwJsxEgI+r2OdQC35eSudG8TSYkvkfaN
JyzAT717JEIF9tP4g/JsqPLr4UBXnt4Ls27xV8IPufp9nzNqEF0Ma8L9cTVxeAfh
/tfYhz31NyuXzwqF4i+L3NSxPsswzAtFAfc6vnmuLcFkExego4GT0MhSpxerWeEa
rm3bf/Ga0mVMurWseLDwpL8kF5K/uGlQgzYdp9o0ARhG9Xewt4lLoUJ4FsoHPza/
udj/I4vpdYSj7VNFtoQifCNJsM1MO6OjwpPT286x2h52E+ty1w2H3+iSfcM5cjWv
AtRGbMYbYNDK4wdZexmcgboXH8CS5ZBlne3RJo+KElaEzu8ur35rebXjrqUZYtA6
FtLNsyKEC67mRww8YSdn2F1AWgR2SmA6GG+mO+t1gY4yFJHuh+Fa23ozPNXTPQ6+
IlRDOwnrmY5M7uCEI8HcpvXkaJRmLwyLAMSH5qZ7Bd0XTv8iayniKpZYrj5oJZ/z
eRim9KZdM8uo8wRC93yHC07/0stVXWLEQKlYPSPvqntre4FcVrmU025OS+Gs0j/A
3XsW58cuanef1V17Kbc46+A81IMH5+kaDzfbBrgUU4gyy3HOLhgMh9iEFre1gL89
azNA3VvoGnTZdQ6rxLztcMem1m7D6yDm8/TWWvdzucn4AGRxhIkrkdPb2BmS9R7B
DIQNDUFlFUVEqscKjFz0ydFEw8xUW/oLFQvODjlUdy/rKKObZ/1Qm91ub2GJ5GQz
y+nbE/MYP9cQo5HVV1u2ivkZaA48x6XGnXNnc4syAojJCJtlM1XPZOMB5VNtwH5O
E1dX3gt/uu1+weSc0KCKe62kUGExzkoUsDFJzzZzeQe8LdIVs1R/p0aFDPcRMOfV
MVSy7krHNSev0YIogQAYQXCujGRdAseBuE2+ln+CUyZYB0IbLymYuJ2YKNt40tfr
qQ9fPTHBjcUOEu1GWA8CPqhx5cXtqJ3oY5ZdZQA3IFJhV8u7I9QuZ5rVRjj7wqqF
gdS0R59MAjaPq8neU3CYbR4BRz60aONdFrZGlK4886iEKR+uPWS6FZfmccvLcq6e
U9RCoQBdLhbr/vXeGo+tz39ba083RMxfled+qPVrztXI0wfXRHl9zmiMf9OGWyvA
iVdNefEUsHF9Q2MbqMrBxkGIwpm1WZsE3fVQTeNCHftvMK4pEC0/0Gyx6+ZpS1x9
sOrjyHUpjE9XKCaJ8NK4ujC14GqA/XCIEHSNycy7SJ3SnTFcIJhCNc3LtXipPkAb
Itmn4Ape76hSrYnCe0c/95CQpH3cVn0WE1jAkjPthOEIrQs0rfSX1++lihiYP3I0
oqWo2TUoPFJYAb1CsbxK8cLkTmmYk/7hhvD7zUXEbmZlGhwwKv4eou+Pc2LMNGB3
udheBbNjOgv2vc7V28bbPkEhMszv2mNEhY5Rxp4wjU9TS2T0dhzPEo49KoawWGZ+
e26zhdlOwhO9O/HzbV6ZQPGW8x0mNn9T2q0QbcdIqu6Yj6fGigqWeFAGRhVP73KP
OgKrV9yegW72YJWX4sooDGGsYhiQvWjRhwTO9/Gadeh1ouQqXzdg8wvDFughkiBj
Zbzcqashy6fvUQdtwHqzvWtv6HAY0jN1ynjjduo1W/kEPAL/d54dQY2xpDba0ueQ
yoMEogTOFmmxaizevwD2sbtUKTHq9QDcq2FTyWZxbRGvtYrPIla4zyBpCrJsWANl
c3TwrA4bTgV/QoCqFPTC/88YOppWkATVrLqPSqq4EGfxT+xudDGrbizBzoiJRDyb
mwngRi5KGtLPH6Egqi92Hr9dMKu+abMj4TkuT13FHDOGJJ5Slbik8apM8C02tzZP
5yo7yTMuAySWwLf6uEB+SD3mKhEEcqABFZInIzT+zmcOAiU1SPpXyi5+iXvFzDiE
l0kXA2yiYuXvUl8AS050z2XaHUdXc5FlaZi6dlzb8XthQ9BBPzaO6bjABAQ8spvh
CjdBq+pmtsQp5Sx4iBma7HcPis/IzzDYl243wtaBPjPeLzNR57AqnIuLfL/5q+uu
uYyxnrnsH/hqMkQhIi7pwi52R3Dx/3wGjokSs3kpA2V9nHgSCuM3qZiW1hU5hbp4
8nkNo1r2vRkiFzxA8qaZtlL2wka1474PAQZGEcu9tRLPV1t578jiRdqepPDq5bv6
pQwwn7GL9l8MDgPqjuS/KRFQwKP5IPxI3yU1ojBybySphTJV4a6TSJOxuY5ECijh
xk9ts4Y9HfMXKsAMSezReY/AagO2ss5JxMtPCHoaQgIAMrIKyZf6Fe2s+Ur4WTdG
G27aZGN0pCjD1G8XtoVYn9h92js2zmlWC1c8ymsputIoNSBjA0iBYbzS6fDDd80N
PsxeQGQx8kNdtWiKD4KlFJB3KChIyD1jTJic1qHfyUUPWBh7Vw6xtH7BwCcxwkku
5AhFKVD8ifUXmxj3qaJghWWi/hzOdm6BlV7T9jG3nQkV/GjT8ubLzVg2DezVmEIf
3NVZ8/VR9onoW0zPoYw5DiPqWYwawIxrVZgw9E5cfoVsIltwm5Z9jUGYYyBp9tpR
D2YElx7ITKkb4A6HlTNPEkEoyGXOrzTmEWAY8dhyDb5vkXfuwznGlsgNCkPsQItZ
WKBfV/hOItXxkNOn2cTe/Sd2UDGVvr3ol4l0SM5+2ndB3yERAfZd3NGn93rWMVoO
nHrlyPtdF12FMa2gBHrdEEQlJllHAtlkIVjukycxLmKwSy4l9ulraiJqD7WVm6q9
rK3hOf2W3FqQrwnyqoPZ5/FFTukm3MLz/ItscReCNO9S9Eg/PB5kx6WdGBE5adqH
m77shZ/pUtW6aDwirKuaiXtpjNJR21cn+JxwuK3wnCbImneX/KO6YHNZ/b2jMSvf
oyXgyeXMGEXKVas8H2CAahrG8sH+mgly+LVWA3r8ttQsongFiFq0DpFbizari6cn
mgMiTVHJNsV51xoe8ky/xWAuYAw3znUiXU1dFY7XS0bgIfxEEnqcO5xfhtuieq/Q
xYvtalG3agCGwB7p59oqJFcaD8aePA5nn/CKrFnH9OUmQ4ueO4gbMsxI8N+jfQwl
sJvMtRQLTeQhkE3OSg4webYvCkpdh+xp1HM+EY0/q5+DpuX3MTCs1eDnkuHatTBc
5FutSIvboVFy1wVjbqtO1c6PAajRpl1COZsJCZzSd4t3AmdE+ypYqsBVPfydomC5
3pzhkzbLPoIivJ4Cn1HOW82V6lPEvtF8Gl9GhnrHgaFmP960RGWX6nwRmAYvhMnu
cJqsbgLDHRWtvYHLCfi2ljNB29UnVm1PmG7V3wI60cTYmYsgvwdovTylSz2oGzHZ
R05bvUj/znGvPLp1EaM/u9rTsug8rITLUyiuYy9dJmlrSzGL5r+guGmR1MzaiSWE
4qUnF7qApE4SB320CsdzTZ3Gg4pXdd2iLe5EmHOFblj60X4Cp3MQKnI0KhFuU+pF
5UCRMV2ki+zvtco2JztOnDfThppQU8beOlQHET/H+sDb6AUxktgVGWszvt2OJVgn
HM/jFy36ess0IWZlhzCj80yJFh5QwnZPT8Fo1WywaaWYGnV9bJYhhGzaIvEg9cPB
D51d0bH8lKM2sc5sMSz9nPJ717IILrb0HsZvVn1GoGG4GZVVWE0BjUE3qZhYFqaS
ngk3i12fwQiK/gNBkw9NqBKjVY2YC1LQucRrvC7KMe+z5wqOwuQ7K95GXFkYYwVN
itYwYi17VMDfPTxFlptKHKv7t3B7nG3x1Lvpu9ctC9JiE0YmqQX0S3ZZsuYOeu+i
qBQJPQv/0UD7W5aGIDU/IxlG/XOMBFEXF/8MeuuJAQ69eFPqIcNpO7Tw5oCnaO8x
ishM3xRAeI1V0Y+tEaRIkq0flCbAPvIuFWljqkc6apAuUEy/sb9b9LSvf4WL29EH
PKMNpfBKX21J2Y+p2/gX62PKpbnLDd7vAs07iJPEIrtopcT0qjO1xn+tDtpyey73
mDmZobnypwu8hWWqqg+U/ssTZKgamEWoc8bR5p9BNCFhDPXoXQR2SLqtQAO3e7J/
zE+TPYPxMJClWnB0uRYfsRjqEwfugNpCIPbSSyEzvIAGWPpMQfF/uMRsF7gGwBRA
UysKlBYUUkSIkRMjoF0w9Pem1W69HwFok+ZmMxabGqmCQ3bqZB4aDwQlH6DDGVge
DmgYruFKJzxT4UpoNgzymjzMD2aGn6+x5gQKsRa3T9bDQJtk5+bPXRXFGH7iyB6J
O1L2TeK1hRd4pHsZeG9AobHAJOqjb/49UXulQO3Dobh3Yu2K7rCAEGLU1Xrt6why
sUC8BtT3h0/DxwZAuv+xQT61xFrIO4cG2KbN2QoVimCXc4rkrVBSVTHBLZHDibdX
6uN/6+uTAKwZ7yfE/5x2EmXpxRLMbci5Sft3nuI3iOnXV7luQXhqrrX7gL+rGTpC
aWbCy3jb9a23fi2h+Idxz13OSiXucVxoifw26I6oQpAtOD913JqLsc+1oFB9oZvn
ss5MFVIyEXf23aui7ROTDLdntnSrl1qNmoJmmF6Aymu53tmEtBtZexCByGNvqZt+
2Jap6VlJVxc1Yatzhj7ePBRWgDFLcaWD7MxQcxmbWEo0LX0Tm6uN12mbHIWmdBzh
xnantSmD9SlhLfL64w/NvGyUxT/STGgnS/HWS5qgdVU/0V4rf88r/wJHSqIJNaoA
Wf/2MhUwC+o7+7QJpz5TSNB+LWT8o2lpi/kh9FhJKziEx62uGRX1CQ9YUpzW+R6o
NKxCYGJSnhpJWcELEBIxQQgNLRNIH/39PxjYgP8BTDEWs9jWH4JU5iXZvnNCXrla
b8tgxsfr16u6DIv3EoKq+RTZi+NKHdnkhOO6kGIf9P9OYBPchj6niBU7HsjbTBCM
SOucN77ILuAf/A1vfEay4c1IoBOcpPBeSth77yZU+sQaegt6enNoQ+O0NVZ9a719
pdzR9mYULa5yg8M11wyvS9tGZ0XaeOR3SIFdhie6TANpKcJb4hzZEjM53SBEl9Ew
xuq40/tAaDUrUPiauBb59ZJA3LFVYkFSj2fU4ujjQqnm9T4yWzA0G/mL2XPEyhe2
sDyf6fmVGGO1wg8dHmmFnZjTRupP39E3IdAzDayDapxtoWUlclrU957U6LJVjTj4
gXeifMyAZHTmfsm2C9yj/dl1cxCXf4Tv7XxF/4t1nBUzBAXbSdnhssga3y8V7hYA
sQfThUr44Aqo0sb7Vw0VXEZiWnslWya7Mugs8jPP8fKTGS/3fxbZY4iDvoIeQFOE
W5Ld2PKFYCjQtdbDqFk2JeHKKN3R+8rvAAkKAyE7gIzP9GhSBQF1ytLC6kRs0qfY
y+tquQWqzF+I77XzBGzwFU3AhW66vNOoJblKiEmBrwsCvex3u9nVYeBJ5Bs1brD3
ev3U6sa636nlzIXTiQd4WeHyNb5mXO8IxhEtm5+ASqPL5mARWg4lIcsnCIqPy25T
o8BejUvxEhvZAVxgFdmNHARQI0ws/pmq/7zRggCIF8MZaoiGajz95jX9d53FIlZo
l+XRb++ud+ezXFRiKMvmc2Ieczp3s1BbjEu5hHHAMrdCpYDWKg1gErD8QH6jWsPH
QHm+P8yysbqst8fGUDdH4mEruupJjAkMPzXopePy30xvhE8TDmDdFSZNtIDqEGr7
R3PhbFRUGppSwSI5gtaWi1Ru/UzBJ+xzkUxotn/h3ipAF3ExRCulS2ZMp0dY4LAf
tBT6/TAm/wBdFCN137TPvUc+Bt/Fr6nLFJVAnvfuFveJvrVODtwN2lLW6wc+fyqd
dBVaNFvvjEo9LuDhOHYtgGLK1OLjNaED8lslm1e4BQJFlKD8BpzFhbo8F2dREofr
VTjLD7i5Jo1Al8Yvf7KKDU9mQtMx76O3ghnqBlfyIeZg+WNVtTIgGF+dJS0tlLQ3
Viyhwy1ATv1sSi4f3O7aM/fWZGAuJoUJ+d+92tkrBg/8rPz+VSz8ySvXKjiL2eSs
7MwF2Rc1N4hazjUQocch9FNnBGVP/6SEwGSZIAbco6sZQjhnI8moejWj5btEjVii
yywLuxwNWQm7zn2oFZPJbLl9JYYYkvnzdwHKwGS/WBaTDftnt7rdX590DLNT5Myf
VGkeTTqYoSqhEtBXaqoey0mV8Wp7TQpx79dexcXzjXT9mioDsa+gSZvXeeL6GJCU
VM86C5FcY0AHIsLBuYc2uYhLLZsOaxcBV0LjKtkjPU0fvQTgl2Ki3v4tXv18Tthe
6jQqwRmbqiU5dtZN/e/ar91sDuIpXFwXA4Mj4ZWA/cEMimoYUP/CzBf2iuAuPSrt
xu0neA3BA8a5wvGaEzhkKgbsSGHiruIeHd/uIX53/tnsAXHaRmNHZ+6Zj3p4Hu3y
k0n+jwCH7JGGZE3O+tIov1VPKOxKK5NotKzPcJvDy/MFlXX6FpRxkevO+PLo83Yh
yUOG3cu9co/8kQ/4sEfmYin9lxsHbBz8XPyAPWpj36WQPGHoDHU43VHvxgu/xc8t
2bxkh3GvRYd8Prk9EQhnsG9GMFkduBgmAR6qA3OcPxn2h2vcHhiezgL6VGbAV4Ef
FtoQTYxrEUM7iKKDavzgSLFOx1K7pAezwwPxSGrvuUQM/YbXci74JNcefJnRxHcF
NCY1gbGfX4TCL1QB85Kq1MzX5CE0GsqZQHHxNX95zlvoroAZ4Ey6G6rf4nKGODDR
Y/4Gp5gf5hpyUmX9URR3hs2Zc8favXhDjg6f1trILYHSOH1LRzDoeRcCM46c1We8
Dzns27GSdC6ZFQukie6yUdqJDKjvw9y5ny7Jiws0SMvAMJvmt0FtYPweyVb2F2R/
CJmrHPGNnolRNOnKDhEWiVD7pDFx1zUnB7ESi5cYz01C0s/yDDEp/jjsgwPC5DDm
gpzOJWHBTUZYnExiYL7wKwvnZcXefF/lPNXlXyq0w/SQBGPgUTmL3OK0R9966BqC
PXc1E2YY2ZQmx48pjElChFN6DkxbEjKZ0s698KHw3Gp1yqb1kMq699bcmwbj79FS
/TsO2X1X8IfbVhxWUbqgF9KlbUYUnNWvjtaYiLJR8bWbhrB1WPnw6FUucnnwt7SS
M6CQ1FxxlvM2vFVppZs/zMnIosKrcgi//0w0ikR2DDTj90UI3StUS063LaFiXM1a
n6wgnKWR8pPo6O1C+1VLh4KF3ImkPmEjmTEWKx8D5W7NYQok5iF0ocx6w0n6y/a1
LKVktMt3jKBCh/ljFEVpZw9HUicrdaHKVyaL4NXWvYnu6nfV+FCwLO1ZSMRaGn3A
2HGNim5TkLeV8twUX2GSWVGARZU6+qeubIQPEt4/6f8Xk3ljVJAWVtLWy/BdgrbY
hWvGNE+ELeByC1+ZelBoCSfxyY18Do0saCGHlkI10JPR1KgoDCC7Ruwid6GPZ88F
XbjbTeKd8s1WjHfIVdqQh5nYk4TNIZ4lfAxp/dMEZUBdb775jwlMroPHXlRtiBp1
JLlGmbw2xpIJzh0qV5Sy0GHQ5WAhVRdIiDf9gzK1ZdoJEOmocPLScm/3uuEjHqfq
5R5l85JoHBjOZFAYAB9vRuhF2yMGBkoQf21TcMMCMnKjhDV2jnutb7kamsNUnBQf
OZsQ2wiUWffVVap22GGcrClrgNBKoddf/iFbWGw1C2F4BJoCKq1xFbxkM7VgSKd/
2f3WibR9bhX4ejMH3g4BGJXSNw58wBHqGV2cXSJggyWC4+FtiOzfOELlPJDyN2M1
z5R36lRFeiDwNw6cW2JaldaTP/xblZuAVw/1aEBxxtQF/fh1eZPC0oDyvqtL7pqP
1if685m2ULpnvGhpSEF9+3+qgJJDOhc4WOVl51y5AbN2IR1uRn47KDa5Xq5pcPUW
sB8lk//wnjUV551MbrkDksgClP6UbgcEinI8X035cZdpdQ6KA/sSLHDtBw2mi75c
ZH5rRfUWg6pDQpqiSnbHAzg0ZNDgDquPcOz357IQc0Njq3ciKhXq5bA+qSxEa6mA
Z8+XC6W4TshooXw6jp/4K3Pz9/Zdhz9ps3eQa0scYtq6kuMiXguHQtcysP2XATX1
9GZOnza18S7NjfTcZqc9wbKqK/yHcp79mGcwZ9MEt6PZMfykuhQqV2D9Ym6PRg2m
C6NVB0Z8hTkUfaUHXhqIoBoqy0h0tjOVQoxnQWubbC/avUVvys/MZ6LxO89Q5YPQ
5jHqzJ20UIQ8P/58OjcC6BFUjuICDrEKu/Jmb79V6fouBjl3KzwbIW9+UmjWu11s
y0sMygThnkMoR/bysltDXmY/DfmrswtbvJsGiom4YSBZ/sn8eLrwBUlCvKcO6THS
uD/2AVou8mOI+f1x857PfaqJYTtbzDvh48bXCfEBivH46iwOiL46WJFMlIMEZtOF
ghDxPXWm+woFXzLJhHyz7kXOqhLZ6LUnTmvotNS+VKZphDcClz4JnJGC8ViZd9WP
p4kJZJi7DXm9Y6mXl7C0s2OxoQdW2dpIKwk42jjHr1Vsij6Qk6k4CG9WZJ3kk1GY
zbM+OFNeGqkxph1dyzjwOOjuVsWRoDBevYNBXD4ky62HP2LV2Fxr65ivimpkTOJH
ARnXuyGJbDa4tOF4NXdKE6QCJ3iJ8ZxBqv699H6tvYbHXszr6tWsuSetEVX+5yWe
fzhSy5ehFJ4tnieKuD/ruTecQ6/NAVfIAcyYT9Bt9hPOG9YTLfEs6rLORbDzl5rH
bGLHwgX/zL+34H7rNO9IzoZnnf10siI0c7gjsrgPfVaLH+XPMmLtsnPMhX1xrhci
wTIKhmYqijTF2q55R5TzS6x3JU/gk8vOiz6kd/v0O/19a3Mn4AvoW+3Ku5hlDdiu
Wmk9ReiylbhXtg6L3gRnp3fFsfWR1zNzgZYeWQ0xDoe1wcpm+K2LcQGIOHgmzy+h
HexqX1XaoVTtBLKFJJUkmImQhgtB7m2rdjOmDTeYWPHci3ZbE9HD4uXuZaqhRvLt
oV60hxxDZlfY6h1DiBjfbLh1TYKHGrncMMrBfHYSjAQsEF91rUz1uuPvc9px9spG
X5B/7Rk+8x+oeJZMDXHRgLPd5rPfNJg7QDy4Zp3lJUtrKL2Wo9R8/LMfwCMsNCO2
i7ZRIYKA9kFkGi1Pluc5AKOUr2nloLeG+k+O6iIelQ0PxNd6xRtAFu6tAjY7rI2D
1YFuSjZagxGzDx+cEwLvv3a159zaQd20hctqZ4PFgdLm4PRh5XGuWvuApxpODugS
zcduE7D2H6n4munUMl8X9Tzkk3PH4MQpDBs6qkW3/nROKIUAt1Ug/bj5sWq/b5k4
dLLBJ+G1LpJxBITMQgTtgOJn30c43V7LdtHtsSx8ae5kRUpZafukMHGkiMXpbZn5
UG/YdtyjsMJGKGH/BHbzcrhpE8uKIiI2V68/4MstGVTS7niCd5qdbwa5VLUtvotE
XLQhv8epy+kmnKb4UatjoczsroEU6JrjwRfW/WJu5vNLQifj1M78DKzPRyYMoxXQ
QbTfWDh35HQcGlNsMq/Zpn3ESUU8uY6n5YiwUbctLVV7z8jeR3zjJkcg2EeGfsmB
WRag1tWvKu4mPqLHAa9M1HQBXL8z08ZDqdMXothtm36Gi/yom8HPvlAAh7Nrc3Co
AIBcqv8mTQhoOl+xo5m41cdoFxAu54fQAErx/HHUaeJfJltTuubeO5q/h2ESsFkE
EWSSNT48mHFgq4dAEayvM1GFQRQt0pH1/ifGLYha1SVh6jeSk/XuK5ztHN6N9yzz
KDDz4M7VvZwe3arlAuFpVWsQVRgMRYQ+pwwpxc9PniFaYdsHLNSvyFcUzH3F25KO
uLNxM9YWAfl+APpbSr9CxmCUuzIWAIjw364pBXZbbLRcd7eZEAC1dfeoEyBR7dOa
tSHStCIOQ8wbPjXXd2HfY3My2iZZvd/O5/q6+kaiqYLmzzvLcnC4GPBVcVCbj3XI
u3AXUMrvDB3fAUWFW0slaU37CzGZpY2k3t1Bt1b6TJwZawDAPNAfpglEvOsz6kf4
/ACsCJIkzCaUz95j9CC7tqJxHqn8Bs+KuPPi7yOb5H51dZIK/dZ38RKK7Ka6+H/3
Xm9DSfQjnwLyj1kVpxyVTPr+0DKOXljBjRd5Ef5E84Ih1T5UxLSsNn0UQaPxgRgJ
9kMngU/jHsuaYTpUSDuh1pPxnvyGjVm8md5Z6qdCQK/0amqa1287gXw13W3Za5Ug
UMelwqtaIiBkbIBMw3gbDCJvCTc0GTrcdVYdsiEP7ppNUpAcJKKM8+jVLHp+akCa
vj/dcLhiTTB1BChf8FjamQSQ/JNf17X9ZBdgdcHljvT2bnKAc7P6DzQK7OBk0w64
h7jvRKymnOlCtGGeGywhc6Nt8xZFJwo6f6TISdHJXRHwnkBlV4VFn3kGSYvv7HP7
vE2NQyqG3FzigIP7ZHP5pbxx76ondXPhtzxlEgkpYfJrgWOM2/lKxJImb2l3N6ma
ilfmb7tND7kDLbTwvfNmEA9EDQQeMRlyuqaiCXimIcR4TBdrxNgI72IxbTauidFL
sE2r32rJCvIzge4m4HL/Hxnk+l0N1GUISLf5O/f4rZWt/Mov+EUxRI1RSSbXd6s8
35OVopunnR1uj0eUV7GyCaZCDbEyThLFmj/acCgolNAUCqyexa0qSPfI4NWbqqq4
eSAs6swdLjcSOczwVnEYn8VojeDL8/eL/cVZt+sKk718wXi/UmyyFtrHihGBZTlS
yeEzHyrFA5w2jnD67DXLuEbCXvWRFWNVi7/emWG5+NIh/oPx071ikdVDZVWos3ya
lJ3Ew3/+ccbicSXv7J6M2rebt6dejXmKp7s8+ffmQWQkQwXlA2BD50bQXXa8gfdz
Uo0fk3dLMya355PcovOUQ5g1iPLCUp/3HCFHXnQBvFUNQd2mw7bvYMzHwU/wIGID
t0R96cv/CHaI+YhpzTuPQ5pqa1V6IVu9pDcv5LzTF8YGSzC+k4q5VhYngaJUvLV7
oKhxEm2/J5QzGJ7jhM0Io8IqcwEBstce4dXkibjD9igPNCzOZD0iW1B/rNMzH0Vm
tDsuNRB1CO+/9yY+U2yHtbLtziP7lDpeTWCc7CWWDpzzXGXUctbRc+kwUBawUvuL
0miX6ZXzmI2Cxf3c4a0JUPuo5HyBm6JFjPqI1QWZT8hfsstC1L2mgiKcCHo2vTvp
aEpUoVAvc+MZb/3f08lN8rxy52MuSVDRvKuOn0kyKl3vPUmzTfSMYQOOE0bBILhP
lDzGxdepLpK7PpaMhXr19BhJYd5OjnQE6+/McUbQfFy17CjC8zX9KSpg7J5jSkTc
I/0L9G/jPyYl1pbkjiDW+lc4zuZN6KDxigLP2Ybmu8WmQHuZ1fzZi+rfQslzoF1g
qu1tMO/gLhYy8ViFQV3mXiwzcbdN09/Cf2WhuIgoCJiDOWqb5985VyiJAEf5odOQ
U5bS1qHW646kMYLRdWDy9siFY0UCk+Agma/6Ip0v6S1dkqC48MyagMw5HuoyADT2
oK/u4YmfMIHxlpYkiUSPeav4E6a/jWACOX3zDAiZAbiex1AruVD+O3w/89EhzUhn
fxtH7UL2FT52B7d9AjbTKYf6YERo7BII5VZrfRAO+rR4WFR2+xb6rnwRLm5oGjBK
gAWJnJNa7Auu8SBNiZza0+OzlCVpGnF5+tNcdm/nKnGST8YZL4CwRTklLfovR5vZ
Rp5t5j1Ksxs9nWl0OWeSuBPK4AnEHeCxg6IYpVAR57uAeVQjI93sllIMfIFRqV8h
QeyxZlmPKikJIa+AMfC4zsI+VPtngenMkKA6Q/uJTJ6WVeXv8US1wsAkM4Km4Int
Dil9f018GxGSCQ01pbV8XFfmQb294dyd50yyORn8GtWZ2OYOd5578AYNlC/5D80u
C6ii+pDriFg2AudWjaim7ctC4KEPlGz+i7qaLQ5l8W1T7IrGsJUMBEPLEiJQmWhI
tQv4RbX7l3Z6/fwt5J7Y9vwB6aaT+q/2X31/ETlk+D0Ojp5cQ6f/gyu17BirlMxk
Np1nYcjCoXgCJ/vlIRYnKl+QGqubytAbY0F/v6R2HD4SFzpEqMvQOF/a+t7vgn00
JaV++ZHWsJBS9OrN8d06S2UvaTou/VhUudF85rGrUqgI2cDI9PxGj9LMvk71w9ve
X+kYGBrgwwnpX/PFvErHIqqyaeeDElk/bPWtuj3zWS1WinKDq0HDfpEnAiD1xU94
6WP37iVfJLYoWBEn/ZSHukjr/Sek+2OrPjp7nCGBOUIH6lnx2LF3YkwOSQXRHrqu
8QDJ1ImuxDIIPmtCDsokJNPVw1HzaXhMe26YI2XxcsBCHwkIKwfxl+OZqQfQaJbN
5eCR9pYX7f+sLAHMCkShvnJjr5P/bSWroyiJjpWgI4LkoMPtN8gL39QAKLx4MKvZ
jgopdoJQEOTPDwnrjNHcgChRMErDF30g37Yvd48gYYDkyf/+di5TnfPUFR0cqsH2
PlrKOkNOLBUqZ+dp6dfioHmaYO/o+Mg3QHXy5DnIezHGpIt3yVZCGNpXpjOV0sxg
kyBmrLRUdX0nILjUAP13L54SccVuwLrWsZTUhCrzR+5ESBYn4E5cg9rfSKsvKE3E
WPqq1IV02s2jG0k0kAYuhgOI1O8tWQvzgL3Z9KxXfTOw6llYn0gZ13+dusa8Bo63
xiaEI6VKXbypN/T20E5iqtNZm+F36vQtc/DtEehFFDPstMVgqucG08DORI9Bqpys
R5qKOuXL5iCtxZxgnYG3YeIe4aMgSD06gAaxvMZHLfoCIC17bTSMh1bM0Rvqfobt
5HfbwjzteI2DrjVgHJj2sJA4WhQGXwkm765GqjliDSIrvgC/E4Q8yZ5gUsV3EQog
fWPip/y+T4LtGXIVLJOOZn7cHsLFBfkc784gco2dh1GJkL52i4JIWEir/FPHlvje
05nS+AJb0rN9PEcsd1vlFV08nC98IVikI9NIlj7n9EjMQe9Lo00+UhJoyyfKJAXK
ayRb2hbK+FDmhcCOXtkSLCXt66CmgHxYYGNrTKcF3ajvXMIsQBTqhHXe80EoSGzl
y7nJPHsy+8Vf4VqyDUYeZZ9MXAx9rR8/60cz8udmnQ3GgcRrDjiA1zB5fSP9dChA
lIe1114p8sEg+ZKmJyEsZztqkATEx4vsBOqmngqVPcObMt/TEWAKlWamU81huN5Q
v18i3fc+W4hFRQBOYYQWsnvojBmUW2of3oUk3rm63vKUCAFoMksWU7mn3Ssjavv2
OQCaclcH1+h83V+vgnAokRsP0CDafBNRWkfkmtX3RP4ImjZya6gqypdunxTFd1+A
srdTZDyiNNNyVXcMYtUhaphJknW0EOoNS1cF2wqoEhHbzqGUBeqKWy7hRDGaJLo+
WGAxyU+RQomcczDdAdVgL1/0TlDLb9zCQ5zk+MOYuCPGR6+r2V4JNSVmnnpYd7ZN
y2ExmjCfOb+9NrbQXSJsUkIy2vx6t8+LlRtfgTHsPgznmScRN7DrEKTkc/1dU46b
gOYXe3SuyBMezLvjnanQEAmA9SqsLLdGxzuAnH3zWC8XujoMPf6fGoNgmsB+/VmP
la96j80oG1ze/3R0onZOgMJyi37k/sOPs7+QmQuAcUjSSITr20yuc14iZZVjVO06
cZ0t5Dmc0TfNU/alUlZtrIh29gKkkCjQ4unnXgj3t+J5C6l37IVdmdetBle6eeED
CnkZKeGI50NuS8K57Jiwnz806fB96jgtKoV3IcIP9Usj5ifCHOXqwac4k/U0H232
KTJXqgrhtfYFhjGzbjJUHrOIbjEwqiwrK5m/3/9sX9WpQT0/T++iayMHbAWKFaR/
lvxBiteudLmkTuU2//slZ3+n3sC75uhEWQOk3E6yCGudpZ7jliuJO8KYSNU9+bjn
/Y+GqX9XYBXitNruk1QnwF2b847fJRNbTvVI6+Kp/pucNya+YoiPGOvQ1K7Uze9T
G9GSLKWgmBQUGv6CHWPzHYVW1OC8tgvOBvGio2jxuTdoEJtjKxtCOGhSz3D6iaS6
x8chHz5FNV3U6gW+tAsnnlru8ZBMh8yrH+K/aeIOQUPppPdUtnv/b/bKqwPQZWyj
wOl8BwWa2YGUQgnTaXw7kx3YeMUGYoX2tLb23gOvULCQ12ee2yJulokoLQBi3G71
Xje+XKuHf67CYXOfmWApTtxk+BP0epZLCLRrnNQ57J1aa5AGqKvtQpIsUdiofhmM
PVk7DZcYsz8lKDHJApSQ/KZEjFOHcVnuLodx08p+M0jrxe3+ewGC2VKqLYk5F8pr
AMpRYaUAuv7ZuOmHjB+EId59Oawwq+KQt9TaUosl0JqzV/XbqcQCxhTsHgkIemjD
pmrVP8IjcfSPmhqi0FuD/6L4AtDpwsKcDFDwzfxEZCU/X8skwAebplh+vCCbx8jA
kqR77uj8ypSfwOdJ8rlZ81Uxk04k8GA4FeqWYQ+D73W2bHTW/VePYKPjLJzcZe/L
CrABKBJLZgvnXu2WpyRKKQSqMa2vX8EeUbdsznD2mHUQPVI0RgD5NZQG2MbGqtf5
JuEVn2JVgg61KGI+VXU6Kvbzw4AadI3UPJjaXxg8ArHLhsBygGjbiex9fl8+IgY8
eAi0XFc498/thEK1UaqEpxtsTlxFMkU4ZPoQ/zeGzFgQUbdvE3cXmwC1/27uHazm
cVFawcsFRFr3UoXt/Ec/uUynmNMcnyM0CFnz9XvUV/46ez/MPmdTUB2FMG7KVJ19
S6lpkiv1WvoSc4A10mAtEY+NyFio9j1VZ54B3n8n9+/tcHu92xCdb8QsQ6k2TWu7
CHMf/Ic+DTi06O4osZSgaaB88aQll+jN0o2r8iVrJHnT9sxqi43JOQH1nN1C0+f3
TSYJyQtnmW8cK0zAXZI7VMt468RTCF/mb6ksO39SUK6PcaGzqzQMEQ6QgL9tc1mj
AVz7QLHdB5YwEIHnRkl91HgW9Ud0S6c5R7Scpi9Q68UmFWTir/uiU0bh+eNwlSCD
ecoEgM+VKaZTT6YTsGiZ/NDyuL6MQLcVAyrSgHmGJCbchi2P/I9OpcfW0FO879Wd
+GXaJYIUUGSroXSAhq71WHhOlKg3axnzWjXijGSofcnYn/t13kykUoH9h4X5JT/c
9ZtvtMihKEH7qfX1nFOMd3bv6eYZRJxqne0r2+MOTKz6uHtGUMtoPadEeMVtBhxS
c/ZQZfIpxsSQQ+YDNLN5yMrPJeS+OYOfRjIz2vB6X7D6gJ7ScUEZ8w7niLrWx28o
zLg2Mt4gR7i2iVe3UMbHVD/J/kQ1wI7bx/Dq+1L/btzPA8Q4xwTXJx6JC6YIiw7U
D3lkNWKGoxc60Ji3XTTOEg8UuEp9BfqchcoBa/1BF5rqABTMd4CXzTSC/Bte8gX/
CHHaG5aPrK9EMzX1Ms/AveOxO1kI8dwaNGRTZWA3qU1Vjv3i+UbG/n0u+NZ7qyB4
+f2FGBTD9TW4Guw2jVWYsFXkv1MphKGCHTZuk4FyyYzxcyoahizvY0/abZy4dLyI
v22RlyWLc7sTJd265DAzqT9QcsyNShdkiwc4fbFylttaexisqVPZmThU6io/Q8nu
3h7oKhuhdPT9j+QHw9Pxf/xbHKjHyywbR/fMsvtKzTyjj1VmYVi/jMW9mw4St8/k
w80caz/3coY8frVQ5KD+Q1xPmDUfEgHnH1nJTANZNf+jpfYbxI7hOIA1Ib8hEuZQ
nm74aYsHRTv94uivi9g/AwOve+jEVIjSqwfjCMqaTu/gS0TPYgAK+vdM9OpuvjiS
f1jwMH+mm3sNr4pL/Upft1TM+P4MpdcL4mUxu6XsQ6XHMdNs+kOJTYbkeR9A93q3
a8e2Mxj1yiSSziLGBCqjBFAEbLEl11pA3uKYF0AldGIyGdJkFSOk3f+F+hkFGOQZ
qW9JYYv7p9Ez7+0zNhphQzfF8HMdQM4zV6roUKNh2+phnbixh22hxgOcTPWQhzz+
YtXkIZQE6gBYLKovQKg8PfoNypBlvyuuxZRkqnA4DP+yBxn50l+JZ3t5xc36bOjI
vxK8cdZ/cBwiIlw8LCkI9Z2csk4z+zTwV6sL+wXD/nzfFYiGhLctpgnMPEGKN6Az
I57nmd328lB+hAhcGY/EIgnxc8YjIURIe195VechbubfkXB4qA8KGhVYcxK5U5ml
gWRpset4gceCpYD+SGG9XMVStzP6MHY76KLp01xLOJavy+u3UW6zjK1UmX106w7A
Mbd6XDsqZK1izW3GiPPOs1/IumwnCeC6ryuY/D2iMT8GHuNqrb3eFC78xThEI/L6
Y3gvHhk55I6IIn6zdjjx8VDinw3McmBAlWaUkkVOXe+CJC7I93Or4kEeL11xXBng
EDUdW4Elh/SjXoQrSR6EX/fkABRQG6q5DvXM/ob3wTXXvPNWwGJ2OVv8pq7rjEpj
42Ulwf/lPn/vO5CcFLPpiMoYKCOL4smiXxfI+kGUOcoqgfHfxNkWNlLtjye2Uwg0
fxWpAfvsRw95gaXDK4vg1X1yk+XoXBatUyKzjDKFJaRcw3tFKccEdBR3ElfztU+a
hMfAF2PIuR9FJcA5rQEs0tAs0W+XzVpRBte5rdQriy0F0Sl6D52LRfBHPaj/I/qv
hz/Ybru6zx1p01Plg4WQ6F1Fqvs1pMvVt8SPKf2CBfqGRdi5oDVC3p4Vf1AkKPVw
SD+lfNHHqVbazJupv9/z6Uw6wCWmBNHJYCHnQGD7ci84gF+qL0Kf6Qh9QSjy+Z8J
QKqI/WDd9Frhqj6jQKsYQi+l2RfCGzJfvdJZVwnbgVOYjCZR5X5CiCUtGSuYQaAE
6dx3ojr66KFRH9+L8dfHASh86J2v9WgY5vzfWq7RDhygWl2HDtlq9ZgXeVw0ZPGk
56aVvDirvFu4HxJM3zFFp/qYIPWPKmAee3wjOn8x2kz+MCqg6oK/5+hz1FysMMkp
27A78yI0vsYrCy1dETO0xrXagU/1c5402JHZo4hR5mCzhz/nPIN8IpG4nu7+syeh
eD6T52rkbqdYdje17gdl6zr7ciEz6EMc6C02d8xmX2lWeTXRt8W0U79HDmXt+OGA
4oH0ajsehgn+nOHdr/1ubWWoOnGlXS2onZTjRai8q0DHh5ExxND1Xet+rfuy73t1
T3rVxc5o/Tele69EP5cupY3Uc0xM+w2dyEmTCgYHcUNdqZj+QC4t8hLhiU6fGH9B
bfp+bq8uNLWL28y+FNWUSCki38g6ysltE/70rhHkpLjUE463yEOXMWASuAES1ura
isHb+ZNHsblVluEWh6vL5uZcQYonfvTE/CfaL9kjS5Oj+A/gYpKQ0lFhilMIQL/S
wV7n5wBTvlag5X3elOsPdG5aaouqX+7hRnwKuQN683aJXbdPWcySAS9PQrSQR6Zs
d+tj7cvx81FyzZt1hNtbTt70PJMA4E2dtPvht4yP8gWyRuRF7ehz1Wmn00gVuabR
2zvn+Zc9/mZsv1bjeyBit6xCAgUfjp0LszLSCb6eXmTAdCI7dcxcTUxjdi5yPkbF
K0Ln5o1zYmQ7SvV5tlTSX7HvXMNuLW63uLkik7H3Qc530XSmrKCabCmc164Uh3Pj
0ussBsmkOxM3Yuq0XR6z/e100VGAXKFtCJJehGFdsPVa/x6BwNI2mlUHEYQTvjKO
ldrVkzJuOm24D1pHNjg1Myud76QfoiHth/SGqgwGzsU7Tn7ZAz5UVZQwTFG/EYF/
tx85Upu+maG1ZKmAO/uNoiYoKMn5ORaPqA3KuoAt3PPPRcV0PxMj8iJq2tOD6moi
GT+/TcWIz+z+YZLzIM7wuqB0hGDkK+/sfkpBpfP40LJuQ/IqvZXrzoqN7tElQ7Hv
HvRm0S3BPdgOftlFmsN0mcfu1hVjlPMYHlJoDLvW9bzOqO7gqb+DrqtMeTM5tFfW
y+lzsPpSY8mO4krowTwNOMqvxQLGS1vxVFdBBO2EfTzGzQEjjg9eyVX8y6HHm7SW
+QQy9xy+we4F+tXJY8IVfEzUtHAalBA/h0Zi0ZBpPTRpD3w3tNoF1cA3OGCHDgwI
WgFEms7jPUvXtJXyxUdbQMHJWLnBm4ZqOsbfib6frtq8UjFJXctCHDGaM5t4UvIh
cI0nu57r/cBPi/x0zxYp6l/uYbUiwZrVfPph1uypH1Kr+Ijk4xnxAatFP28YLjc0
eg5+LTR3kj9q5YQYf9QF5OkxtXPWoEFzf0ALhKHk5gkTF6zFIp3qSFrMhF36mMHM
zNhqz4gMr2ejwLGn5QlaA8+WDbIkn6rdRSbvxmyclJ9hCnx8EtHJqia86PhTyG62
m/5tRYdtSEKXo9rbGpiDBi/qenUiDSRym0v2khD+XybWz8/z3uHc/06iuTTCtLv7
+q6413+jqJvLwH/p9f3Ho557FKb+mOr0Un7Uqew41xkIMmXYizVMNnc4SCuo3hD0
Lds71/Urnaty5y0eelooSYvj6iFGxHUPKkGF2iXHufcBK3Afl8v0I5jwE7bm8v2c
ZtknwiZC6tZixeV7hVP0w3BsT+6zA6xYGPa2IxsYpOnOGd6NWJs208qrmsnGh0E2
HUesFYO+fABEz44sEi1bqGgu8C9DMiBtRzuOI+JkmATykM0qbsvS1c4ee5eZ9rLw
TP9hNlRmvofwSp4np1EQaS3J4mNu942pHoLq5hneVmhaGG+hNLVZDYT9Boe9hIaA
n8isKMQ59gWimIyJSAbKCwTqCtUgcNI+848dKaeadHv7tb9v0lY30brDMZ4OU72V
2eV5rverrybENKPQUKPiwUSWF7dp354MTwu74yxLmtuWRlq9qQDbkEP9v1eGKqJ1
3ozOidagT6N6fPuPQBALKv4bQC/o4BadrzYUynql13u2Hymib0neCfAJvh46GaOu
zLWuGFi1Y19PYIxwy6mbJOCkVFtmG+x6XUkhv6w4b6hhB2SzU7HzHsvJ7mNTti/4
e1nHZA9F26zEIZ+EW3cFGfpq+nJiXKhoCLJcA6wdjhtcsTffAncbnS6HDcXwJh+V
zC5UzveBabP2MMDSsfEPgxOE2Jpk75MZ85eWzCp/82f3ar7Sq3LmWwmCLGnX8AEr
KSFP8NM0LRsHALOTtZxZEd8A3h3IPqwgoXLI1Yp9AW1nldUHNQzkxpnrCg0Xrpgb
tC4SRWykjkGU6CmZp1j5hX4JvRvVz5UDU7Ei9LnNMLGJUYyIBpwz3aR29QWBEy3e
G5bX3uPEcfC1Sk9KM4A91X+bN8RdCI5jgU1OqMMVbdTNw+Nzf0RGBMqGeRDb6Hm+
jcDcGrjKVEk8ewi5qJFsoySgAbtR+4iCkq94RouuvMefNkXjSykOzsm4Li2K6sal
bO74BLjDIGYJSDyO2nQ7me3TB/Js97iLvSCeqHkFunjxv/n5J8CjY9XhFdMIR6K9
V7IIj2KaaPz+UFQ7zBV9qSgGwDz4CWdY3q2Ui2y0mNaSdcJNPgVP4LAv3vVNV4Wi
weoPJtKY28Hw7C+JS8vsir0H2tSra5OON3JtxWaApRShclvVRjN0uD5eLuNEG3ni
vfi0l5qKXSysg+M6VnycXm99wESXzhuobKdrX8FyPi5kog1jNY/gmqp2ow35zQRa
YZMtCpzglCpFPTKtrzb+pPQa1pPrZh3jnx/u7urYjzalW9Dqh8o9k7MnFS6FNSRI
o3Fk68fDsrPQiKIaPj3SC7LE/W9wIyYVDjPCmt+0hNjrodjyvTlezuRNHzjZyj4f
0HMVjV1455K/4beIgUVFHpjpL1SHBNxMa1/qO8UATJXW78MtrpwNwFj7sYagUSku
N/XuLWkM6UhXdjdwLeL0ODiVMlYW+famViTAWZwXQ/B695nmArEu3b0Z4pv9edkg
3+FVcmaOgUoOGKI89m4rsd4W/VWJDEQrLJWHY4hHZhldm6OcOi0Y2TY/hrvXpXx5
tiFI1bKmhXEQvrz60SNGnPnOeGFwtVnbLX4zqeYbHpMr3w2WdBEdAhdyJxKxER7C
d/u2yTnCI8/0unA3JZblQ717DZfQameWo5ao45wf4Y9VBNH4ILSisr0LtEpEbOYW
wSG8j7HAcFzmwCXJqntf7Roq+AypvCHsS4Qw9iWN7NqmkFy0/UquZhTVW9Wp7UIM
8f+MNQza6fzWc3F/xkh/ZCEEfgJbMKZcvKtmrhXW/rGo7M1D/EwWLwqACI4yoj3Y
Zmw2funB1dxApLstiTCEiv9PFz/fLnbGPxpZP7zibnkXHasz/sYSqBZZxRiuA42I
94M/QnWYhLau7R/srBWcog68M6j9bRm6Ga3vp8dS998mUBablFPkIFrO1hnk7jtC
HM8SPxE01LE6WLNyrCE70vJmB0IL0JbEe8mQK4UvJaJkEbqgx03pkYrBUwNPKUXK
AjxbaO97LMCidukNUN58wTVwa2iFWm7OmDiEtCqNTgicNOGsM1smJ2LIzj762XtI
ywi4VXFvaivu0PG8On1DJtNYE9OJBf4yjG1onoE+f76KkfwVJHh2xLNVqgQlmeGQ
vJFb6ouYJ5ZIFOP5SIBr5dY/Pvj/Vx7Smw14Kk5ssB5KJ17tSCVWLXx20RrAEyrA
vemiCCv7WMhJhGkLpknbHayO+LkMKkw5Nhc2RbXNagrImPkxo0zptG2co5c7f5Vh
g7b2gnuVeQyt0Fwip1avoLP3iyQFJ+aziMwTmmYpz1DF+uxMRu0EkQ13LSFBYCYv
INnqcNdcKK/x6uuuF3VZ407TjCVbxc7PcZnSgsCZh93MsQA0R2DxxxM0wg5L8CKV
iEeevfXsSQ+kPMCEAsJbSQ2bj+MUazO7NeQ1Ia+GGJ/gTQ24coh6xR5TkRRRnzSL
ZQgAu1YJ9+TdaVWOrIwUnaSVhjFM7mVYAJArO+u0Vc5HujgoMLLcGfPuGS/wCMRg
y+Mu77yHQMRyiQpF1BmeV3QT58WY8P3OfRH4qQEyWn29NawOrdKWx5VzXX4dhgfg
4yIW4WzV7GDXghewdG+EmwLimrK3DFvPawT/nb6USqIj7OQOeAxOVkXMVhcuSmv7
VY0EwN9S9p05JNV6yJQf2BwTjgna0IGkKrSqFkU5cFxbL76M6VQ5/g2L4RfR83oN
8N4+4mOkLNkvaEx8KE56xh7zOetsTk+mVP/fQuvcZnhuRQbIjpLFLNGGs0vmlDDN
lFP8Bd0uO+jH9N8TOqfmngYgQqhyC6QVmfj+add9mdb6M26GYnRUcLFIC6X+MrCe
GgHdztFIcrfkt+y1IUn1AV8L3hHze7XjVES7auQ85NDLDK65WnrOFhm3DCkJqJ9Z
NS/S2P5rZ/pi2+oa+OIItC8bgHOzxH5W0yDBTQzdMWli8t0GK/xCnzapVH8fGDKl
qDUAlpUHTVPd0sWqQn45xSj0pVhYCyk/yZgQJd9agRoJmsQ8Zjm9sPWxhY33vB0a
+b3JkqMUlNGgrtsezoCGaSkfYYTvkhfCv7+9moM+TOOZ8WJFb8RNuqD50zFsyT40
QuITRvZnJqSdGNwaFALuu7S9z7z6+gsP7jNAqSLuIyPpwZG+PnRzyKWL/I0X8BV1
EgzmGvbBxEJtgtv/RA36spytmT57l8wnqM2R3i9trB/qrEpTRQlu7GrOV59Pbr5N
JfKXJcQaOcs+Mcmj70+nsrTxE9/hCW4qXtmgPd9jB5Hx1kYyKRthpDKZjgAOsuH/
aSYPEBPKPM4o8ZIS/8VklyjXKSxjz3/VmFaBuYLy8bhz1g+waMT4m7MlVTCzpMGt
sBdJlNrQr+nNoxRW2s3/7UTsDw2VKcGY3S8bG+l8r+7hymmr5wLOK+b8C7de7c9+
DurUrH9Dk5TxoI4ZPDIY5NHpABalGpqxAfL5o27cwzf2Dv+k6hrr2w9j6JDsMUFk
LHxgjdJ3PoeEeFNG3B1bR41INOQ+fifV6LuigFLQ3BVIONE1FM4FgSeNAS8rTi2z
fuAfjDzPlYqDHvWOQScwxcqOu/Xaqfz/JV2LFEIx0ovcLE/oidiOf3SYxh2/cnyR
+hxHvajpiWJ9NuV0wZZLFXyB6YEgMmquflvJA/CGg9oWT3QmN2+I2rZW+UdBgNNf
YKrdmMvbDWdT2OodzMuBSwTAbnEkTOKm0uV21YPo4jwbO7VVYeZoWoP26VMRT9UL
JLLdOxJwh48TB8+oB8sHm49Jbhz7T7+e6QsmLVDRh3337sUjPNo7VK8Hx/PWLe0d
flsRwd+d/ScNcz5dCJ/8iExXdOPcV/lyqiEVYWbEvZjSN+tOmS4L2VtmeOI7upLu
RrjWhqhrJ4KnQceDakJYBFHtQO8qsuIa4Ib+/RNmyE82vgYMwOafzCWbmJ8av1mn
sX7K6QtSlZJPPOOUcHvWU5KMtrVyP58QZSjwpGbJubDlVF1CwZuzf2QevBQIXZcT
3ttLmOPteBaERvoR2IUAgrZjURQrFJaNq3fv7ZsGIocdXoFiZCQLq/47DnpnVAKl
Jzw/x9wJWVJELrxzk8gpeeopUo5GGwj+ZnPJOWqzlsXZ5mtHNqPeynxrP/2oWMm7
dQ8oQK4vkdQJiewfBTwDJIQWYQ8Fgf43mC2OMfgaNUCybqPKaQHCimNBxvC4yg0E
5P7JdLJNIHjdVX7nNadeqFnEtOzQvRDlsULW6X7iM5adZSFatUYdABxA8adVGgpD
AbkEN0LchGgSbR+CKfjoE5NHQ++GgboAFsdlvIvEBF7ARpvHu3UXghjBizEz6Xme
ScO1HLgdGSZnK4vQxbNu/8lQ1knx7cWo6CKUZQm0/7zgRgoSe/z8GiKdubw5hpcG
gGyl4XIEJQUHEmaNLr1CzrXUICTJ1sNRrh8Izn1WvWOzHnUiLHCaiuSgTbXv/UCG
d79yiGU6bgFasDun0r91eIVXHMeouITQiT9kOifJHJcJFav1J8vZJH86N2nk+WvM
wie3PZgBktA2+09uO+/yWqWcEgPex+iNDlQEA8xEBDHjTk78xFA820cbsHu5tFG6
ql1YEEetVQhoqdFMaBBOIAPY15F6GepKFjpE9zhSvZLrVhvMc+mhpwWjPzuMq+2d
VFMPdFalpMSfg6D+rmn3mpWnIUNmuZbEmE9zJaJ+KqMguK55aleYA+0hDYYNLJnd
6wY1eNVEUmzN052la05iQb4lXfOdOPwnuXf8DgziZtXdFXvrUB/V7qIOWBbak4Nh
Ox7jGbPQcbxOAcLRnU+zzmJx0+SRyfWwsORKJ2ql+px52L8kGBRbfseFVs9yN0b/
VkA6mTDvVPnZbx/fVk8eYrDAEhQucuJn1cx73hocZxELFsqMwPQof34pHxEPhOfv
dk+hrA8AfAV9LZdMDlC+DRf2xADGCz44VaU5Cnc47g4shmlq7NWc+QtQC3nw5/pZ
9ihiDc9QbtD+2rJ54LETsHUPAO63nJFj4tpvD9KQCIu5ooUu93j7otZ61cRolNso
JBJOxpyKkwpM5Kl815xuq9WnBkc/DuLg81D54H6l8tJogRGmhscOZqK4ibQDWT/y
g3Hy2F5+m61/UqWgNeGUvCCquCGBgDvEV5Onq9UwOVm464O1f99hwrp+IrJifN9h
kdseLEOslHRY9TwZkZFwPlCJvCdUFF1B6bI940fGIVeVlwp2ggIBUWqrGR2H7GfC
hIbkGazKHBg8DxIiTXbWK7oyS51xRDVOTin4OrqXOYnKzZnHps0pbKLC5yyb84HQ
wmGfbqgGlH/kG3ULFZKRzJSBQhh2AxnSNCNmrzNOHtImXA9vgPynWdUAWztqk/kF
/E69xPoOuQlnqP5g6TLn01ThYuVFOa+aQxAJTdM+5+V/i7n+tmoCgOeTrMn77pYy
9Nupuys2bbjatw/+nW+aAIXevCPZy0j3G9iW1XdSGLXoBwWytyHd7gJcwcLkABPg
wD/uxiaU8QTP94xj5rbXeQrZUNA5ZLbaibhVKznPConJ3LZSMsEtpND3hBMUuSet
C5hjAzEuB3/jdSMG6kldGYDuY9BK6pp8IIYh6zN1OT3gcqBaIes7KoovQQHWyHvp
KLvWzund4s8aMA3M2U5hZKTguTTtqGN3VbTltPViHWA5ro/2Izhcve+NsndEqi9I
GAa9mqv/gFuQ3RqKfimgge/MFv/E9uwVS0/CPA55Q+/P2ZxxXnoGvysatkmnUckn
qLvLq24O3aZCYVQzOQh5VTc66em5XFme90yvGBfYBLfT6hsoeZwD3a6iwdXrz35v
LR0WLUl0AZsd7xP9zDXQfrl2Ul5R7ubPv4eCioK8fEYnvQtTr20fzRP5VIwl5fZC
PF5NxduqCoaAG/ULiA2MH3hqwzNceIpvSm4h52Xydu4rnuNFKg059EvZxuRyPagX
78iktdoAWK5cMCQCPmTN+sHEsDMXUFIFl/W7lFobwxC27eVfcThwfd9JlzX6gjCx
OJISTsaE65lTwbt2rfzEbH6KsbPf8Q186YysCGKZQKNd2Gfm+8fw1MAKyRsjjE6B
cQjXwAJ80pWmtZbYndxaLacvWePX3rAps30XVhWx6uO3fMptdueHnfEZigGRm7pX
HvUlrDZBXrN37GEPhbRBYmebHErQ29oX3pxKDcCy4Eqt5Lch3Eoz8jyy4psgNO3U
ZVf7IrctuaL4eWcxmru/XRUX8yyzCTfbsnyczjQG76BzPrYONMMGkqiSw1v4le5x
DMhTm6ztlfDCnhzHhmt7Ft+URynxTyRhQEzaMhhcoM3Li31KU0A0HFtjjW0BG7QY
vijRqbwwUYf2vqhEYHVAzo90lHunk25Kj/yieefWRFikkTMpCJf6rRjeyen3kjCp
c7gTqQMrVo7IuhV1jXnU56yVVL8c1lTjgyGyA4ArDhpq0tFcu4iPBXLcs9UqMCHK
RmClVhjyYESBm6TU+Lohs4QOeKpjConKN4aKFB0E2ud0pu7dpvYfveYYuME84CIM
lQvsu3vS0KD6FiZ9A7awp6YAGKAipHQ3FS+W+tqPUqU6jP7owDjKSapVKwT+SvPs
SBzoovH7K9YWojzZ91tYGZ3Jc1eUhK3FGGkDuxdrPdqYwqBwAPVNmUDwYbp43m8j
ebaz/oc6rh/7WfwVl9yJnxLrdfqQFz8ztEYmnUaZdmSbYZkK2qgW6esKrh8myQWx
b+ywAUvlLZdVR2t2MDfYyxC8p+0on+24sEhDHOI/hrXwOi32hvZXruiK81xOAiJk
kEaGaXP7BQ00vef2gKEfb0UlnZ6V1IgBRIPf88gihTX/odjLyxL0Mt78RO8omHSz
qzfUSSqoahVAdwo1mhMRCpcvfDzuYVFX7PwWjxu5HRWKuORwPTEACDEijlEC92J+
4IlOs66YrIYYLICXur8Il260v8ZJfezDeNoAXfxvbM6rCcDB325cgjNwG5oz3BpF
WPlhDdsKHELc6OBMkESIOcszJqYucUGQm/o1LGQs1zFOdEiYzxBKz3ci4WnJWQnS
VciRj1TwlsLyWjHv3ky//SL5G5y+Upc1uQgOGFRshetZNG5kWyiBTPWg/uA+SOQb
uU4u7WEXV7Hy2Vs381yo3RuTzc/sWemKHWa7I3q3TBD4xp/MZFBErxrhs/mRgCkR
CPPWo7JIPJvKKUYJvrrCrvS8mdehAPL6PYripj/Fi+O6xSO8u1O/TtMPyTwFh7Rh
xlva7gZfFyByMrSVzUxX6drcbnRWr691YI1segGZSigFcgOdY1tc6oHJisCcoIvV
tpbYJB8/9QlQ6dXQ1cac4SDSwO5O4ln3rX4dBTGwInwLL9y2VmjG3ojgLUgR8Avm
fTvW5q8FNlFVkBRAmTTIDv+XoNDiWKbvhc6n+Q7xNJ0DGnmrJU/1Sn386ia56wtW
/n1lkjb8EVKMVw5Tz76hxoZyuEaUB9T7V8qmEFZBRjfYV52TYMsrAU6tbqM8PIuV
fTj8NOZuvUsgbwDs3W4m8Zq9DJLTIBlW8th0m8qlhp3cyDOL/0juOlK5+N+YP8Ir
cFLoZN/l2kt8EVLbFJexaxBC2nM9E6BUvUldNFA1Wa3QV+Pes9GBqc2SB9ekAEfW
ZxDbua7wVLpdy9fAdMFxeutBp8p1q3J+Kg4vqxKnJXnr5ZRZ/ktD/iK0IxKlGuOP
en98J9MA+Pg+/a37p07EUD6to9Bii1DgXDsxl6MRnGqbbCb2pxMNukA+Kw6gjsTm
1eisL+RP6MDOnxjRcMbJi2ZedqA0uuO3+5edllxlsKTNFl7dvfb1Xx3/3zqYYtqP
2UcxsZ7yxA6fB7Llg4vWvywV5bNYBXgcHPKjceZxKPlx9sHZgHCyrwXXggen3UBu
ROYeB1DySqiW0c7nu5hmvPz2BTV8y4ARSMltLjF7HNZqJ1wGePPrcKXQeknmPlAz
9sXospcPjthSbRFfIdnRDkQ0dQWUNwqekO8qzRfTvBxwv8NMSxCSUVqdNLVN54vU
+La3mYpFIb3cRrqfee8X/Jhk6iLIoJY8dJdyncEg748MBgbmgF71tqQb5JstdxDz
GW5wGFHbt6wEm07aqDKqFghNyEuRllGGBhLd2VfXoDWeO/3WHHnksR7ZCJGw4wmT
lQ6SBlgzbKy5mctJWf/1D5tTJlPYbmznsnjktjaXMxFjbMAmPAqA4+R4BLBw28pX
pnTNa45aCwN6QqNLv/EkNAowkN1es7SWX5arQcx6IPbc7EeXc3KS8YQI1ddqwg+e
v68jjiH1fATXy4exmioSuD+ndUojkw1c1PsQEIVkVRaXXltS68q+Mxh8n0ZsHIEA
DUExizMnzRXk1Is+U6C+VMa4j5fsN8HZ4jE7A4PpdoQJkLsl1RNE9/YFqD22P5m1
Y9G+8DwIQej1CJlSaXOH1ZaxGBdLV5k0Jl11CPmENZrA7antbrAyn1hyqgSyREzK
eFoHanRqU/GssvY78a4qyim8MYfOXuvsizG1X50tQEl/8yqkgh5pit/3YQ9/AlAg
2LbE2YZXim3fM+EXGOhSSzifJDI3NM63/dgFrXMBQRCt9bXnyFMTEiUTvfjRPcSJ
JfVr+xHX++Ik15+y+zNTskzpJTGNs63ILWyN+c2sY3oFV/VPZouFl3JYfKvT/Q3Z
8Artagj9jZH06Y848uA/0vnesmblX4JJoMDbYf+40cxZqR5OqP00+DPGcXpJKZpM
9QmHG7NnMI/6ZY6sxZ0euz8gna15XRPXY9e7EWieRa0fXKu7sQudZSGN1P9sXhcJ
08MgAaoObNoBVEOEYJIMDH77VBUr4B61keYaKfv/TBxS4e8hwZpRbqVjo0aABgou
bv6/MvpzegumoAcM40S1j8IJwPyOwqEZjBjJby+jql3kYEeAov5QtrWt3MmywVA4
PVmmHcKJJy6Fp0qpqwGnhw3BPUi2Gt2RhjERrOl1G/021mLvFNDa6CL89aVrnpU/
DTfuIm3w+57TyfqDFezbgI9AWVKXQSnK3kYG5r9JlDtIHpVKIJcApDMclEH8e2/F
SS0GK9kJx7pOo3bvdfTnJmsEf33HChTRB1JBVK7vCgpems4p8y+sgPcEdedK68Lo
kn2ljOPLqa3uFeYkpJo/RKMu0MXBUD4OwTuKJG8WSIFA28c1TJ+nUjk+ANB5Tjkg
mYmkPFmBKw3jNr0Fl2d+bz4LmDJwHF/ATnLxwTO1jSMFwYagCImd1wG3OviRq0a4
EjBrpnWGmQjlNZ8J6HfpJXAnZjYCEiRzQ3HLGEt4YIlgwfRCSNkZ9u56eBDLlZKT
ffmBviiYIs+uyn/unqW+9TmRZjxyPBcy481vhmaO7NWcs5A/VNvRfDZkwPrXH4E1
VJ4FLQAlsUL8jb0qOPWJSSXFwG27D/LOP2EVsUZNuWuuEJetI5QZBluTG4ZBKEv7
k4FkKhT3HEXilPAOthmYyeZDRg5Ff7zbLGJdXFMlzEjW8Cy3kaxHjqfoOOqipIA/
H/vekCsAST1RhY+kDvp7i/7YYBaXuTSIMdmOZn6ABGUV8SbdHDmH3SJoBlZQPyUU
ugiPFxaEdURsZhsD+gVBG8vXJ3gXzWNQVOTPAURRf+BvuqQ93Yt51zlk4AAezPcW
ZfYHK8txnJhwd2gsTHJEBKFdtuN7GyuyFel26YLhiW1BF9KUNamiVYmzGHV2TzlM
UnybkYJi0NyXmmGaR0Ym3SsjNubEeWf7G8am+zVewOtlezp8rcW523gXzPOLnKK0
ydK/dTIFv3plXxf5vc6VVwpGEka/EAAUOIUJKo/BASZmvO+clBeNNnMcuATsHg4+
ZdUPrLUZFHXWb6mvdTCqyjMhdbl0YYmgopSrTuvM9IbgPUkjdElJcwfLADwc5KPE
iTes20EsQSZEXL4Rdd/xQwwFBRxthmjfAEGBM8FQJ5nGZWRqOGbT1YJNUdot5g6G
woJs+M73SNvQIAQMHvYCxyb02UzpDM0Zl5UlUhx84dxM/LuQooI1FvzgAJjzpsDB
uy0UTNH03ZOPi2EE7LOfC3KqCqiZ98bcJnXpYIuVNRKF+aBPNNbRJSemHrKj7Bq1
EoC++SOlZgPc3PIj/DjiaAHQ0ELvCSYrIwhfWj3HDIjIe+lZWSISWC+aOkEYATUB
k0QjsGzUyIXig/GpGmBPlNdHtg6FN4gxPvJvw08ySsFnd9Y4Ob9ADb5cOMvmNshh
1DTKzkBN+v/c1hDwcpZWhAQBfC1dB0GTyuv88MAyRdm7mb9TWx/kkwRX685HTph9
y4g0vvqCmp5lqff7oQC+2aZFuZK77KYh8oIYuloKRe+ZzKHaLLZnlke60Kpt/uEZ
DMf6Br0fTIIQ+GM0Gr9w5Q5NNkr7wgZpg/r+qLlGA1gLveX7FmkZK/Z2h6Jct/rU
IOUwOjf5XAfYgJlbnKWrnOBThrthotTwK6/uSazZSMQ9Loj27i7+wPHNGM2l5W2+
5j8OIFdqZPAIlkrFAprjNFaXjjK2oDdebSxl4gkByWpkUH9YyQvnkp41iY6MkJ52
kIcoerogFKjMSUoOcsLe5mnaSoTjNgfPkFw+CQgJdY4Yz/Unc/2MG4rV2GJ5TCSm
xjHiz2ydos2h3yTDzLvdCnqGGkuqR7BojvKEnruPbXj6qSdpfHMQOZa4YAaYUuAA
ElOaRWhPSw5WZklGdgE9JexyOTOx8lejujO+vf/1qk0yCaTRGzlBHg5mH+Cgjw2U
tvMoQP51WtW0AmQ2HSIJzRBa9lkMIetdya6Rg7nF0bzTpY+bM1H4K0G4hkneNHJQ
vA3QP6c/ELCcGTU9GXG60ZhX9ahRHHv2Wxww0DrBBN6w4giL1Wy81JUOt6uKHq2l
gS4stJs6yLzwdbpznFrnnk2BD/HUZ5s9Hr55PO0Y/Ex+93k/kcufzlOvVOJTqusq
GGUmZEhqfpAv8N6XnkT7ZXVeaI6umk43A4WFgcEV3X7HY5Oaa9zaqrPjz6a0mDk1
TIvX+xYSLavYWAZ/6Aznfxcxl+NMcwyggeIhgw5DS6JXBA6S/rKeQFFcaRSp165j
7h3FY4maOpsw4yvUZ17PK5wi1bRmvBDRzz2vFVdBH68lTv5kUSkBTVYBlWyE3+YN
jRDrNrRWMg3FbZzFCH7V3xJa6zLSlTH+KealzPquldLqR6HRi1jC1Qi39byyac6j
Yh9akQ4jZrq8bkbCl5a5vPwVtZ+LfqpeX3fTTNjqtfUTEu/gk21jsrkqt4fUKK7R
6ONdOVPkYWy0++/myB53y8h1AIC6xlMUm0rncluBEqsSvSYCnUThq64L9uL2+Cw7
KkVY6zhSg62u1gTq88qDSwnI+14LTLy8eK8Ej1A9xGxzYmLEaB79ejTYmzB/bY3x
TZcQp1DBcApBqSj/QPLAHvLV9KTbQNAdZ3GZ7QNTI4XK4au0zHDO9vzsT32b0Bo1
mianxhoZ+yyFlny7DUwTAdPanbJa1CPLGdNrQojuQ8od6+r/OrjTPSWxnx857uV0
Frz4LMqF4kxSBsjC5cOmNt072UaWB8KcyLd+9Xtj7nPk8nzyiR6LftEw9Lk90FGT
Jhs/LSH3/rbxxIJCv+1QJ5EVZqgsrAi0Oai+oN674rDdE67dXzjgRI7JOmqV/UKi
q5pUA6uy3H7JtQCa4BEO+nWwSQi8DvbFM/T0utCIFVBsgIY9TSXqDGLy7g9cPLTh
YP/PX2zWVHWNWbn/ZfeyglWT9Gc0k1ivjz9JkbYGs79W+xnSggi20TJ+yBQzCzwf
smHNXi5M315iR6T9U9Guh7QShAG6SE+/ZEvYlXKrg6laxjc/hcxzoRXxov7qaJak
bU5+zqjQGjWbEY6cMrul8Vdgif3goQ92f2yl0pzxaCeNBHKpYojl6q8AnuVwiPU2
TRX3L6KkbLch7baeArqko3JKhNVoPIhx0rw5KTRJqY1sm0YfrzMjv9kw5/7qT/MP
oGbk1mRP7dk6K1pbKX+p+wMg3zqfFByROl9QZVvXjmJUFlWiJ8VBkHH96NitODr/
BC3gS7UGgbmc10qNaew/ZYZWohVKl6lFVGLRJZ7MaxNA3l1FoR20f5k+Xn7M2aQw
+c6iiNDqZ5dmhXTnsW8loP4dPyeIT2Qk+m+kgAbNGYRPKe9vRqdRqoGgJJV2On5O
01en8Sv0R3Xx8LSZDW1EM/YG0T6KxiD5SkElWc7K4por1XXArAU0N7191MFI/rF+
up/TxT6Qr+G1FR1DELHQhWt2HynjfDzGjxNtk5hrV8R/jlleQXTpYQiGStSNILel
LadTi4TpEncc2+FrheQ1LY6QyT5Sy3M/c1i2KLY2jwRP4Xz0BxesTi15pJwNACsm
cL3Xc49j1lCXKQrjDIIIeo61Fy2vYl3/Css1Bnm9zBpW0vP8O08oIaM5945DcVv1
JUls6F82E5Hk5Q8q48KAGH0kJEkFtXHqOVeQ++OcHukApI6P1eirotEirYRGGCRc
NyiExpiXlTymFSV4W2oMGi/Pwm33qCcfV+ekI8vGhOd7MV79qGfF1F/RRLqFrvCV
2Crgt/AljehdPmOAxJnwRVUWLq45FJ9/IJ87bJFQkC8cOUbk0PiWM5acMTIc5NQd
X0+nEZ2An9nNg9eDka4EO9xNYMeAQNAJnyZ78Li1hzR+ey8xRV5wCvqpvtLghFiO
P1r4f80RxkcLVMz8oQdA+o8Sk3MOK6PBjKkHKBpubu6LX9ErKLfim8Pqd/xYwX3s
lKsAZBp3XydhvxKV1ACYjyctxr8rqcthMMR3mNYG0xdVagXC1pXxoQf4ECnnSUAT
/7/yiGeeCk5Yf3ZAxe2v13fQHFKtcgsSLIA9BtxCV48Oc9jB0mMkw2eLsgx05mZ1
Mb+2wpyGMoszNAH/8PJv14TP3aXONGNs2UHBk+ZXqG+RvpIPvJSRi2XIJKyeS7yj
WeF4aSEKfoOxametSXiz0ZTHc3juRQ2oK0lljfmsdUjEgyIvQuDu2zlN/YEkjIRf
j4vbRdYkli5UYs46ONN/BH2pyBzM3LYUMPtRmMCq8ycGdrXwUYvm3QDaMXhCnJ/W
Fp9YHf2ngbFybhZIGK9NWsspCWnrVf+66cLSV32DQ6nyUHaLoqzVR0iM7NWOFEXa
lP+cBUQ9pN5Px0Obi8CTtlpdgrgkXSALjrbvbKragapX9Tt38WmDaytSqfAb5gt/
NzCaSXTX5HhBXpoH2QAjSh2veaS6D68Xxv9YWf6QRPNIoVtQfhTSc8MgByPwyI3s
LQ98z762mFJ8eo0w2A/alt4QjBsagQ9VvzZY2edBiJ6RtaBEC30Zk+AV/Ljd/fHm
HC2nodHDSa6ZgRHc9qHbpiUkgbqI8NrR1XfzswmlOFten5RphNqk1yZLqfEYgAG6
oX7/xVKtJdI8ml6wc+QpvGlyF8s15dhr2D8cHb1aVV59GzQA4aVP6F05gAcPSQVY
xAF5S/uao6rGJVU0g4UW5rtPXMV6h33Rp3ySMrFeW3v6gHsMxs4Jw7JrZAolSlc/
hiZ0VlEVQI9rG3JQeIkmweWpjv3P9GQhUHKSXK4RzVVdb75SaFxIke4SxYygdSrx
JnKZ1eRvLbHfk1ojovbJzcQH2XZoydsGnwwb6AT0lMgPITe/Dsa0Ou1NdrdZ6wPS
spBlgPDpPUYXxI+RG4yZmoJqn4AXsXoMXU6T0dJkU4AKUd+YbtJ41L3WTFFmZilI
GgATI5eGUH7V/nivtcwEO+upY10HUMDloVmEb8IY28M5SRqKadZrHI98k1t/LC4m
RhBFhtAWWT9zHj7t89/LbyiXn67z+6rGiCfHWRKuqQosU46Aqgax737a3ztmls8r
4VJMA/9gVof9rStahX7tgMIApHKu7KxTKyYhpjQS2oeU2+323409nS2XCb5VSUke
EpVT/SxQydDd2cmBFkeBZXvJgwetBttRs4JFydDILmyT2sZBjAsjZrG2isM/M6k1
iw+NOQ0dTv9bGlIfdKH3f9j5E7g0T/MicjoC8Rs6Ox/m19ZgAVrA7Rn4JZJBTQ5o
TDIOQ3rFLL+3codZFP6Gi7vj99M6exl4fHUMBjRVE9VC/Xh/tSYx+yCadWov+MBi
15vbOLwbNLFPqEHdXtH8E8pRBgVIMXQ6vb3OlMPNwoSFJzAMBhedeoCrxaLFpJn3
v/p9mZbuhoVLiJPf07indrUywrcZ2G465LACaOaMjX6x93d7xfI3b2N5R4Qmz5k4
USeEz+PwvCcthNFd4l2EkpO5WsvkJLzohk2/DsiTWd2dJk4Bs2g/WP2VfqwmHxQj
X5Ts6fu51TWP/txkAoHFlTYmAQgB+nWIOkalEBokkD+gFVi4sIsmanCsa6OFg140
pcJJEIl4EPTGUOlnUNL4Yibgfykyzt79SuCpdIn9cXrFswn5zkAavDTttXszYFdB
shjwIanC4iOrWt/6cW7nUtA4kgDoFgUI9ZkGvEkdjWqVrxYzZf3r1qERGo5hByol
TWvX4QFH/B3LBSWp09qLqCYkaq9yYCxCYC6AFigRX+3R5PSsRMh6R6gexFfaldua
XWQvuzAa83NKusXi4ox45x/D+s5mHcT/NobIIK1pEDLFC8GvcPOll3uxh11H2GPQ
twSCmDZdkLGylaAfxr14ymxpATorxIAaOED5u/bd87XjWhWWe+TkLvL6nRY1xZW3
UrSfefBGhoTzlt4QhOtLQJO/Ko/XzYKFaAGdH8pqVrKfx6ZsCAM2aP7tX+dCM70u
rnmU/wu5mNdkeSbNE2UDHLonq5gsagPHhhvTlqMcTJP4Cpdclwn1gxujoiO5PeO4
oHw1s0Ob1Sq+Qcyf2KVKfN/BSEYqR/wLlu/ZprjDbLGZYnKqtnX+pogaphWu8euw
Mf5w+aKXQ20092xYHLo7VeIQ3jASZeKwrIOJcPnISHyS91gVEvrOVF8GqytkCkkp
AFr2qrKgw0pEVfLuq/K1d9wszK+WW2LqyxzTGSHT6HfeoT0Yn4iX2ruIoLNw7SJR
q+yp+82HFrjio1BiTPQKjLUB7tqHE4qebPkk84+iV269syItGiJtx6bL+D4VUJ/H
ghEJ3Awf7ix00M6st2HDlrnV2ugbQAvaSip0kP8jPNRl5/S0lcfMS0AsfTkkw5ED
LumGgePfUJ1X6PDrmnNpwIAvqdv1Dj+cXYtKB2jSR9uep9qjH5+Q7cvkAvle6+jl
Cnq1jQ6U5qLtodqXAKIIwOzPy1OaL3GsfDBCkDwG4adKlTDzMH62T18ErrUgRC88
5AT4eUClHGcjnJlUVCGHFGU6ueFlMbTs+5XdqRX3R1PQJOVWTJbAOvy0x0Rn3jUI
Q8IGZ6QbaG4xHxWyvVOA3GJ5pedFXXqeO+I6FPklhpKru3svDx9d+MKSmv781lkJ
5JJfkWzUFr4byYaPY6XZ9kP6CYNMV34tRYDMNJY35yFEi2ed+ZJyz75HsmTCNXJd
EfPdewjhPuj6uwdqxyaOcbBduoRatNxpqmQ2qYIEOWtc+Sw42Q/VpD5cb1Dvll89
SVP+k9uey2FLMrUTGuQdonlZaNHP+n4T08u1Ebvhn6RBGgIcauPU0flOemm2Zyc7
YEXcEUwZ/sJrLuSwTrXVZgIbsTOFNE4ltxQ55yCQtNk7EYRHF2UvulDN4D2xMG7P
yAfeopkZ/9Y94i0S3X/D57EwUK7msqrRyA2edwqMmCTFyaXR+VSmFO50CfJ/NTDz
dLCd7wOdeiv8K+mc1hgkCs6qihl6anMQ1g42wl7kSLXrP7M36reOwmr9K15bVLpF
MkIu46iMq+IfWfbQmrEbMjDjvfRqml4GRVGuTNdLkKpoz/QtR+esjxIfUrUcIpKF
nzDpCXt9ugeyJvlKKmjq+l+Epq/dvzSUIy769y12+JhWfuxoE+EEPHOOOnhyBjFe
zBy/i81dMlXrl7s1FAcIWB5IJzFRxObAJkKKNTbw6C5/xWvpj+G1mOEER7spuDbi
9FpkRgIjShQmvxtRFpEW8iyhLD0fh0gWjMMZ0ZyX+sxLjuJ3buH41VsH4MXy0kb1
/XwLori42acA39ohKRwpIo+8Wwt3HR18l5FRJp9AY1dic7bXrgx/ryotiCcRrVUw
77YlO/mIEEyBql6pdOCL3yDNLWK9Sjxx+vnL6x6hEbHhMqGep0yP16wX3Uqgrxux
R8DHn7eWA9B/UkmEx070e/5FAIlba96fvc983iIvbJ5alZugkbhm4NX8dEHOK1yu
ByHZatkHoFqnHQ9cKC2JC47L/k9/fKHW0V72b2jhLoF6Oj0aRwGmJzU1wmCbQDVd
mynGX4iV6M4nqKZzENLcQLi2wqYTK0lGldcz3HQHm98Br6KkWwGUIrnb32N4pOmG
qYhvSZk5m27wMONpSsGh36sEvwUzG2A1WqGQIS9LGFYWRaYOheRa1bXmsuHtxwfx
UftyDsnBG0VJNmCLI4EdCGwjwmdL8CsLV6p1RafMy2+1KocJiiuwXkdUkp0JItjC
tciC1zBVP9iKao+MPBuWf+9hPLRtU8lb0+YI0mcG/91OZ81MK7U3Yvbw8cO2qCxg
eB06zM3Fab/bZbKzEKrdN1noG/x8ao0TuJQcRLRksWgDNc33yOZYezhCuq9A2h4x
CSXhyRBOar8cN0YJUzFKf19opK0Itst2mTTl/TO/ahG5jPoIjhB/9eGpmO75nZuv
033jxLQMHSeW+adOJIn/5w8l4iAIE5cglprp3wt94G70kDY2XLQjsUAM85iJIV4J
fA7VNpo3I6WCMPy3YlOrQULTpjnr3cNdwkEU1PjMMG0ckT15lR54GD7/gyY2yvXR
WddnU8r5Tr2CfyLHX5S8clC1qI8wmEKL3Yua+H8mEaKQp0zjzBKk2gzdEXT/zM4U
JiWBJ3K6Z5m57P1zzmmwO8l9iekOLM53szUHIpSGGER0xJG8czq3vGGRhcFnJ/il
B42x2rfFsS8Cz+twDuooLLhwONun0CtFpZL4rv/q4h3kXFYgW9snPnDCYf64IuBP
I9P88Hva/MADn17Ib5Y3uPkWUcH9ib9HKf6Sm/QF0AsqCYv9tQtBsMFCVyO7nd0X
47Z3ps07RjRFbleE9qKMxDMEPJru6jXACHEtDWuCLcVUNbTMHK+EQCe0DFmzvFir
KdADnh/38Q+L1xfKgKQRSnRmGF52C1fGFEPuid0HMElKgqbw0gHfWG69+89UpaSS
L80XTeABfUBY7DlkeIwE0BwHkB19UDisusgC498lu2CMUFLqtEEP8PeY68oOPbkH
mGtlBlgJLjxRs9LrXVvMMeCgUpe1lMRt9u2DF6Oh7oa47fn/jMuwcgZODQ0BiOET
HRIt5nYTgv7EEbodaGsJRdtcAZW+XNiEkjXZSk2icr7QnsEQ4FY5YS10G8zMlFGT
UbrnzpZcCwbQti71L7SMcvqQ5rNcGw80ctUct6GsScN0ozQB8nworXwevJtBeYNb
tcnbXMC3W/YQU3bh+7pIONpypCxYpyxhV72P1S5RDQEXslfUDb9dyRAiTXmiX+p4
8rKLjm+nIPfFY+uPNTmqC1zMV7dPbL7ZZgkb5D9VmHlEV50Hf6bdcGtiI/ZK4932
Ca9Ov5g4/dB5+XAs7p1HR875cOLqR/AeeysxoPqRkDYgp3O1LvaD3I9cy+EMsYIg
wz27grKfdW6zrpkY3cCzrHS25VEEucmkDbznd0I0f5NJ9isSk4BwP1+AjeBXhDVG
u/ida/dllLtnKYK/2537JtCFfOQDX4zmETW1fhMgz9GUHBi+mbFKZUZTgBmiRTeb
AszdVMTo1QvNAnYgWthy9T2sxcFo/PxHv4GNQnm1JbnKevmo+b3v/AZ38QOdEIEF
bIELtfUHeOuzYeNuUU2q+U9UpLREFHDiUKVZf4d0uOAR+2eejHUGZu3Hk6A7a1X2
9qcY6ObdD8co6tViGZn8zueJjAjUx0Kl6nwcoSUnji/G2epKdlTZlZ+yW6WgbVHc
lWzw6uF5R4LyCVJdumJ7ZCAHZdXBFrr9PSsUPxj3NNogX+uIoqN2WBN92aI7ZoV6
DF/YiVNWGPV/2dNEAaPkREWFT1YwaAXYacHIn3JmeVXidEakc1z8cr8/4/bwNp2j
bG65bFjsS6Ft649LfqSQ7QhJcmOhy4hY8Df90qbU+nBHnwNMn7nTFIVLKlXZTjWj
9FKM+hkD7Mnir8gJmEfgkeqdCeFwoGkXjazI/sNyCy/adW60S15geqq95MApTTpu
uM0/IUXJdNaoXa8GevJgWGyHQnA5PgTNSUJV+9aij/uXqf+zJlO0T0eg0m0ThX+F
xYPL7mhg6L97w4SljIA/xJzWNN7zwwIhP0jB9bp3AKRPbfoRCqX8vk+6wt4SVgq7
av1ANUTiVZt+dvVvHbPvYs5WkE6xQTlTphJGMrq9mTUg7gVi3lN/zbU7fnaZACEG
LdohSoHgQbnO2rZ7zG2B4zJC0dCv4CdpVvnIc26D9jvmrFCda2oSkGkMKib4cyc4
9GsS98yERVYYTFdb1HhSGWKqctz6UCCEUgttmrWKrso8CON7ZW0sbTWySYG/L4uW
XW/32HTyB06l5BSBSQkAVTV4XA7pdz0k2TWnEp7kN6Am4JpxZLoRqrGHmavpklqp
R9fa6XryUnCiAMhpjHvtws2raEerIVgXS9nyHRuqKp0zixYLcf/ovgZVFWuf2vLC
+ZST6+tW3Vjypd9kxQjhuGwsJUDJLGiGTG3Uf/6DEAoMr+1symmXrxWVabvwG1Xt
vwYyzo+zRUfU9+Cyo6aTAJvEYyewp2035hwZ3o/M8selbM5XYpGGcpBg+Ax9KuH3
9HN1fME1cE2+cMbIiD0iayMUpkpN5wO+5xqZM0BS00y6J6XB8krem/2NIizfVRSF
EWYe4hMTtBrEKrNarflMpZN6dwfS7EbzY4eNepXlAdB1SNAWMgs5Mu/KkuSEmWrz
6mAR7Q6Gr/w95AruceS32r8YV0foubazRRdJIBx+EiXMAQQuu7i4BH7eqdPRU2Pl
6mMNT23BMlx1w7WLA7/Gq90fFxmkgDYgc8OM/M47E/8kioBRuoqCtmvyo9CIcqWX
1JcqKYogyzNpPwBS5c2RXreKvYWvR7QhE4v/3yFgpHJqaxvdG0zJqoRW2W9zbnZU
9SThWjaV1vj/4wd8FXhHjd1h46UDmUNUmLnubwQCQAt+usT801a3x57dHtqZ+uoA
i9Jv1rbD8ZzvlnsZrKNi3NkNao4+uLcIxL0GgJcDQnkeIcJpe+UIZ+/9g1StnF5k
TWvyilpMkascPZ3nodluIvu1i8mNfOcsnPrX6KpCX1flr4l3BT9Q64am4X93vhWe
BiemSVtPZxHs2xl3T3BcgvcRxCZXRX6BMtvqvukUg3fsao4SnybxtrltUEVnP0qr
JghSBc4MbeIgFvTY6ktagi7o/fBStflbjZqhq4+Ela2nW843eHM8W8bGuv/xV9El
EDQqqAOUTmVC5o47Mru9HWm//obQ41Z0yQcgyW1TQnfsN/bmA9715qLQqhOEUxpE
S3bJNPw06XR72HEIOEVbYYM+FsYpZddZnOeUknhXzerAh8IEoYAZ6aZJ6j5MJzeS
Kbb/rQNkUttM2RSBvwm3v3s/buyRAkpPqd6q9NrZKd2mjRhWyEFOrharI62RrCjO
vaZFAmumlNl/P41/Z0juJ160NKFOcbLyjpb5VZ/eL/E13pDqZIKoj50P/jaMz5Ru
3HU77kaHqZlpca9DNGOCadt9Ky5kia/ad+4t+3EgqrnK9xapsEfdRkHK6o9NNv21
o+1bIYRd+TjdHom/Ju41FRvsq1hgyQxqMaZrVJULmvS7Vx5kK+CkoAR8b5wQ4Jy8
Sq8c19datnpEI/KwUdu1G73kDd32CLMLhLNHEyG5L43SzxSMaf4fCa5Be/utKhLp
IbQR0gi6Rs1gaUpP3sQneFNTaZAOvutL8TuGiYoXb5Z5o6yLQn/ZbF+n16T5+qRT
NosoihhO3AyK5pToptFWzg9HwATWhdFel0v3bkiAP3cCnldRuiwzpybStQbk9Kgn
GmkmS0GAExF16PaQhXUUiZq7CHpIp3KYLiurtWDNpdxWIyKjsai+GMe1MCmnWzkS
sijjEeS+dlf8qe5uDfmVizhylHr6UM76URxESaAyKrq41psiNRDomYpXpI8Vghvx
ixo/nsTecIsoLmxg/d6/Ob92p7xL3Cjw158kzrZlrWMmdWc43HHk6Qszy0Guxog9
Ba0UFJV2ntHQ7JSEfs3h7s+gl+zLI5JvnAbZyLrT3fRbzqZ/rjUMntjzNft712t3
iwqqVoTfEfLVFZg3yd3Q+f8kbqW8deJXPyxl4eFYw+zyv/PQBX+VbQd33UffWpID
nNaMUntFngbfxQqiAYoslNEW6u40IZ7Rw6CjlWQTU52RHvOVrKDvvUDePEqiEnui
9DPi8DE4DAJSAtr241086D8jb/kYnf4d1AgJE/MuNJ5Ssfpw85IGjOEQNII3AAB+
hXMX/Bad3QikBd+FFAXXn6EZPcgr6JcDjHHQuxIOWgDm1VgTTB983UrMopnYaXy6
Ss3ZeR17mr3mb0Ka0HlNoJL47bGs5Dm8AYmUsIOH4az5I8lP2WcX7q4wfX3t4wvb
LRccYWxDgmpFmklub3I02W7kYogdMvUfkrE29M6hBPQ/O/tgW26QCsrRfdWU2js2
s9NH3dNnkd9pS4VM8mbTmO5KzDZ4QpXJfzOpHQWubeZbhz409D2YRSULwjbakocZ
mVknce0GCbtArJqn0/iXclzt0V/e0/cdMddLz1WM1mGuq1JqiZEQIqVfSWYAorgg
r5LH/L/Vx0Cj7NgoyeVHQr8Yl0CKd/zXdbjp37TDIisdC2hc0ELhAw9S+fBJJh4q
TGX9aomeScTLi260HkS6kTIQB3Fu91fkKjUOx7E3DbQ+bUvSGEjl2YhYa2gjsYJL
jp32Qk8/Kasdn0kMdhzlVk5jKROj3FqUp8gRyj1PmhZRJh7jzCsWjsJqN3FHcG4z
QHPOBxdxHXNvnolMkuP9i4h4NTdmmooIigOATQ1sGH5aiVcxcEWk2bHV7gKu26ez
nzv0KGcJcOtGKrR6adXseN5FwUf10cRwqJZrwE9zcEJQmOvmdGpunidpuFP53Ekz
QVDj2xHyTmCfUFhxJPMoUyq0/yD3bg3gK3sS/EBv9W2Su5PpvHBWO/6+ZRfRAqZH
bGMk3w0z4rLuVxhUYQmFOD9K6HvSE2TyTB79UUfwio5pf2btS/voZwSQoCO+97jF
I6mQc55VCPH3/PDeAFg689tsXmDPqS8iq568/WS19TXiHqw1PGUmrfGBLMAIOvah
TpYVdsa62Bz6KMK2rb4a/nMUT8/sbPKtRTOrhr3kTbU7IadBLiuO/OsrW3boqEgn
7HnXFjtCKBC0pDcVaHG3Ub5q8ewCQ9np8pN3EvHk5unJnsP96LE/XPgZC/itZF3S
VwsAi9pnB/s33dKNxoIqgLFOaTZ0LqR+ESdgnZE8JKrMqgBEJD5fvLOCkDyscHeb
w9iCz85BnUfeLgkWLG5r3QvfGnVPhg2hjrzh6XNYUJlZUlmDGnywp2iAB43c4YVr
8vhp+lUlVf6rr/xdLTkmpJ59QH98k+ktCMhCRBJoBl8XMMv9vamUGE3fT5/saHon
sUtXaFRUbr29JFab+NVMz4ALJtypG+yarX+f7V/dqzxoYD7Psg9l3mq0hNyWQjd1
ucFuFmCWEDfwzdwaumRTfvTjHtomHvb7nUEpW0+ClIhO5PrelaV3fQdP7UT/ctK/
86jMOctYkTUvTxhbn28ek9KGZZFOlKYkVLgjlB5cICULn5yMgT/ZZfwdBI/m6Gqg
B+c4Xn/PbCubjU2yBrU3PJ4SvpC3kADrkJKR9EmY5baXcys025NlITTPZU3LeyAz
Vf5g89eNq6AUmeEyxI8kX2dh1gdzFL5auGssup2Iohp9sVwZwoNsxiEC1DNc3TAA
YUg51eA8VJQZaywLD8ILNuB4ykEXg3wMDYHs2sMtNvSMlvOZGidHyRAv9bDnAooT
UMpUDU0ZT0+4gQEB9sPiVZimjaeKGUQ7D15AUgu6o80WZUKtlcagjK+BP5jRQ5UP
amAdEtL9oWdG00mHQDin40H40p+YwMvHVd/lALQpu9eZ63RlD/7dEqZvxp9hPmsE
TXnVGqyuepasdp21ZNgzjScmlHy5zSFdYSHtnHR388qpvdW/ztCxAAeHsufRqave
+FGDoca9DXt/vmQc/l09/wMnbSuJOU6fUxZShiUeoZ8D362RS8ejcb72JDJqNOU0
bbrkpgM6iZNDAT/2TgVQYIRh+Mc+4eBuj2v4FxK9w0OY9+3W6Bf9Ww2Hh4JTZ3Ny
qZEpHk/5XsqdKjlDun8kyilYnjRlF1l+x/Rn9TTO+NBt31E2pTyQybgNdq2od+8l
ZxRs+5BQXynKepKd9ugqzo9wKXLkzuB3c8vWjLQ9Jd2OFNDlY/1j2xsuiZs6U1eb
L2ou6L0gKua1qiqMVkEdR142WB4FCl6u3KnFU5YdGzhJS6g/pFH5x0jp4k41R6nN
YjK2IwfcZyMvDwRhIrgXvIi5ihLQmVe65Pc9PV/aForUWHjKNx5arTKUEIszhUd+
jxR6yyvM2J4ofdj/DciP8/EVjvFb/vWW6ykfWPlXmit5WYfv5i9TOCXUmLa6C32S
IEqOB1XjHtbGTmkGWixPCJlOB3J18MCIQojEODcske1o2kC8lqYMoC9dL/BROG/n
DfZ50wzFidH/zf5f1ehXG1NyPgUxMkT0feGl8ZrIed2n8Zl5M+WxBU1HIf87GllH
iKn35bVLq01oETHlzpPH70gknz0B3qHxBscndMwE7sG5m2XGIIKi3a8VyV2hSJ0M
qMvr2MPTRVqvz1l9ddbbaZNDzUzAbjLAf5xP4T0vVHobWs6jFXjtf2+zJa4g27Cj
KA397I+nDyAP+zMUw9O7eJ1NxtEgi9rDkM42LHN3u2Rla69h4gF2tr/Sp4LYiniI
DtOkV9SZV0w3JQpFSn0HJNG6KKfaWvPVAmRfuAwcGm4Tir3tjq1toHXp50uAe6Am
zeOWlUfl8aHFxKZKula3+UpR0/Vw/D+iCNlLuqHCAmMYGMzgjks2mtkskjI+3GwG
93F8Ep4MNxqaX8hOIH7aR3AGBvU8EmLhfU1xAOJLRv1dnmxneatC1XHv+XQ8pymh
Ze4sjkxM3qIWB3EUMeDTZfSZp+NZ6/Kncz4CGfyA5CADczs6UIHwKEAZmj4AyeZQ
PPJqp6NNr6B7eV1NgH9PhCWUtLWAAf8rvaOtetsPWi8rX3+noTdd+O/1W5lQfyRe
j7CyzI2JzIFolkRoOGf/tlCcygwGN5BK2sdDWfvMbSOlv8bhwP+aKQ5EF+BVkDvi
99Tpghk6zp78ccJivGBwByyz3EjTnawsXiUfnje2Xd2ZObhte+fuVfKYNTrvbh18
elqA0X759tDJ7PCQC/mM6bB/4Mw7yYJ8WQ44ZGeCTq6dt3eOvM9VBLWPKHK6MLSb
AO5zICMw3wzuN6yTNzPSIgsqtI4H0uHR4RXw8heDQTVc5IhMG9RW+8/UMhsH7wQ8
EFesFkCIamZU3HjfcTtrkJJLQX1pR2FXQhChjrs7SSrhBONi9P8qLf57aBHJQjId
LQBQw9an8SqF1CE6xDRh1tgh71oHLgUhyavMPF1MrlOW9u577XTHGFgy8UiV8+qf
d9OZwpLLJINxkxF8jwCQX80ZDZQHVwJEaqxeJpFVtN+V854TgIzr1RCMRKs/BIq3
PCC7uQj6FgbJQlNcFIhDnOyp0Cuina4Oyqn2JnPl6gKAI1BsV4iTYXnisTfb0y19
hrKFN7bAI74qnRgcbTJBbqOZIQJc9wxqWlW9WHQj26ek0H3CypSM85bmpxfg8NN3
atQ+bJvJ11h55QkJOOBnZHtJ93+nkyiKwvv6ym+in5kckUH7130aKH5t6rzR51/9
1b+mJ/ZHossFj+/r1FhwQjQvxgQSGKJifWDMGl/UTnyZtMJmBks/0fO+/GEyuMJx
cYGI093gyHFshRMrYIFbkkM6jwfAYtkhEV7oldGr/7xiLQKpi8ku6QajepA1z9pV
nMNAeH1OCVymlczMeRYYteUpfDEO8iAvzX8KKeye1KYOQ/CBs3GtLLzT8LKpnFwV
oRFtK7MHsYVY11Cbi8rbkNv5+NLcvIBOJ3jpdxGqmCCj9GHTf2KDcJE768F1l8Vp
vcvDXUmAGQhJfOF3lT7N80Q+eCgszMDbfRX2FrH8SL+2Msad97haG1xYFvIO/xdw
ibJdQ5HNZLlfLv/0Ee8MX6K2rIwa5jIUf7Iib3Ku2+z22w0Mec1m9ue7MniqfAu8
ClOhVq+ehI5opyix5K65JjTZhDXWMHaajHhN5ni06b2vVn3ch2TADRUJ6MDXl1Jd
9GX3On7H+1I33i5bdQj+qMIZ3umlvFqxmXxcL1unijTzsctxja3nBIDWJiBmJpIx
16bEWcANvAXEdt9ONL/6E1nUln+zRXUYd9nFYOjivpLbkv/dFt5YllM4yoehxoeW
fxQUSZwQnE6oQilJV+ReedoHBDL940u2BiwxLhta4HKTEv2wtqBl1u6o57C0UCv4
SANGqOsxkawyidz/oKeby3d/+28oD0L4hjYbEW0DINPspak4Bx7NL6GTti7K30LH
/lqFfmj2YZy+LbDTQSHdKOt59loGWBkijaEMcfK/Y45B2PixMjvXFRt3uK+Ulciq
IUPAtKMnP83s0GU//my9ZzdCqp7U1wMwhiseEOvCensgyQFgs2Br8EOpAlvFcG6O
EQZIKhsqRJSJIFNgnFEBn/KAUwzJhUvwBS6IQbovXNqjOj6dWvi0dKXyRAINzcNQ
j79UBpCClFWNsWHXOrsRZHQi5hM2Jbz9rjg/4IuNJ6T+ib+a02vNdlzIaAUkOhn2
5KuiUEAKclXYbOIQqJbTcDP6SitInYiQK47ggR9NpUTdpt5uRLnYOP0Yp/ddJk1I
RMyZ1t/Sx9PKGQeJy0U7MtO+UFTp1Rvf8TWEGk0bnvi/aDD9pNC6uHIhFAb9m5c4
dhjApufkYeNZvktdJrptHyCOf0W1p12Ct0Pd4rh3w9ldxHrVncsij9Etd723mXvK
YMwirfQsisEikF8g7ttpyzacRIBh2yg8Df5kd6wOo3zbVQsfkFVm4gWXmYOEOy48
dKNh49wT0o1TLUB5w6w0Hc7mUGnoC6YYuVddE5LPekqbD3m6d+T5YJ2h3Y9Jtj7x
qW5U4Fw0jtq5Q+zOz2IVLj26NKykHcibtYu/pt7eXzahjw6vloAvUuSQr1dWLosd
9Xl3TxG7JV0CRy5JwZH9DjPJmlsnbpRLfdSFP2Z36F2in+l7Gai11H/QGl80g91g
h3s11mg+xiRqz/fjVODn50CwNPVw1Q+hJRXJNefzFSY9i8qmwSvHmp8f0T1WR2yf
7EA3ZhI4sJjDC9a60RdHWFG9cjthX+nxXBbeGZVYeLpMi2vwPtrsXHQUjOJ6h3PH
sobZ5ohelNoN2fuZEkv1WI00yDnLeGXUQpAh3UTJlRI8wu6Jpoy6qBSQ1j1AHT2h
YYwfp7u2/ODFkmuepZVvw3TiHiA7m6wOA/ekKu1ERuX+lT/RLR/OF/fuK3Pp9ibc
RLR6ahkebkIKMBpVijfSQtWJhxlTU8ScRIh62efGEeOsucFweDCgGOCdcTIh7L8x
Jh5r+iWhhONL+6qBTmgjE36DpDe+d7vADR5qArkjAeFgI6X3Cv81u0+IoJXcH4PC
LY45zBI94SmOCHZfgNldj5nyEzlEXQ2aIxx6rfKPqrE0d7omXnJ/8BqdK/4rvo+J
0AWURTBz6ywLTIFaozygVbeAvKub7u7+Bf+c8fZ5mg1z99UfYs60xuB3zJKTXURz
jddwHAWgVyO1z3zk1JGcSTNck8FtTkJezE6AvIdAtrw216oqgY7RYrg1dHfGkvoq
9SBzNTD1JSq6X1N6DdWFEMJJHr5z6/9Q8KlkRUNOB+7KpysfKDEHTGTRHUWXGH/l
1FoUjOKztWFz3FwtwVWhSjeiY9DMetMqy+HjpkvsmlG2BTF6eM0LFjSuIAmhla27
9//PuC2M4R6UBZRvYKUQpqpzhAM/cDl37UC2/UBKgLUEcUw16pVYUBu1DDAM153t
xWCgoyQHGK0owsaIQTsI5Jn6GuvdZlZZkNJzKe7+Rf3vyKzWXJXgpnHoe4U20kmC
ESEuR8++PO+nrdkfYe6uYnLvm8See4S7EkpmG1VDXgkWel7a+sjHrdehJ2rdOZ/R
k67sDbtD61tpySwM5cbBoO3DAK7Y2iygZxw9YOvPBqKvbgyEzPWSxu9PYmfSayml
olgib7dyPoQtSCCj7BuFAQrye7cgOPUGts2wX8MWenRFHC71TeVZGAQN9nlN36js
VVfnVFNllsfefl85C5TU4IL6vAplsL1wH/rlvuWgmWz40MQrRsSji6SinJI5yfft
B9ki2tPG/WxTeDo8svdVys4OXGqMtsy+q+oVB+1/z9ztxXHQLkQem1qWrCyzG6uJ
N5dOG5dWh3BZsVOv/9f45a7C5GQk4eWd00+tG9f3Ms+fnIj64bq7sqIcqQv8adBG
E+3+pgvz3vM21W2UJhv7JXyxzlyC7UuZ6OrXPtLD8F+K157+Vy2/TCIZFGmCQT0H
h2b/lOeUioRmGl3h8BJxU6IN+bhF01tNVVRTtGsgdDPEVe2KmR5D2RVAySH7lq7g
KyyS+yZJ4iQZrpbxHQekvCA4rOsgzajI8qqh1FWWraYxaCU6H68YjU/g7043liVE
7ipNSExWoy86qjsIJ7i6XmknRTMFTd0arS0zkImrWNbON45T7z4BG1gO407C33R+
xfpRnZUR0n6zSdXwJKOjnAPfzi0skmOEoHWlSN72/tmPa3whMMUSZm++Cd3lRye4
pa7bwBsWGMrzzAJ8BhzgAszKSnMBefDzb/QtYCQYK9zhJF93PZHLaiVJw/+7ZkSE
fyZ1kVCdOE4G7RB7PVRrQrqK5+pqImicCd7oW4+QqjO8fO3OUN/rbDr6ZYenylKY
NwH+hMax+SiuhgnUVMCife3sXFYQCdCZeJOCG/LRGt9akL0TNGG+hVywQ91TIWKv
cYFe9NTAVuBQQ1MniqkwIPaLM61J54wKH+LohXy4a0edFo9WN/1sK3kaHwhCSFuZ
EE7PuB+pbK9fXQPhocNCX0jglj3uCcakC37YBU/Mo7nPc1pEY7cpTY+wpSHxpB4M
DDDAFWp7HdbThiVTRkgEYVzlyySTjESzSziQM371hTA3sBW9PXFkU3FbZf3O9vAw
xjamaLy58T6g3rR/0c5cukDQOOBBQ72fE9ktRjsVsDTI7M6N7TqD6yF4roaovs8K
8JqMNDwpyiFFOqPHcx+Jnx4c5OzFIeMn/KOQJ4umpOVqqspgod0I+9J4R3NuV1NH
m2fm+QlV1n3ku0Jk7W3PfyiQLwYjPfdq5VgvArhuYVI9MRPHpWyoU6A+CcoAn360
pcoE1FvJETiUkURsy9awEq0zaGPQRcHKqcdH2rWt+Z2Z3LeD38kqHEoz50/LsLJi
o8SagVVnr/AuZyEy2BDHTkhGg1flgebfHOH1NywWErJIhkClPMKbchMg9kRZe7YW
GZKFePXvod85Yea9wY8MqlRuxTfSpA7oALIaQOxqOKuYtsghqSznvzP+pDAR8yVI
mM6G6NbBSm4CyQ8nt6f9butz2t5GBVAX8uryaCTMSJS3XhhnLojzqNOvEsbl1BoT
TIExda5ylmzHmYQfEJ8Hdphb7ZVcgUitcD6so0Rs8osYoCPMpzxAMQ2vNNWAkYWZ
h8Q+G96LTxxxa2DU7FIv9QGQvHKOFmXy2HhfM315XfTrpTzB+ua/J8VUjIu7XYXL
VtWAnX8tjQUKCjwxo1MVFFS/kTIhYqvNHc04W++5GpdD6Cz5MGALFb1stFLEwIum
w12erF8AcqstcpVZAIWDR1XClFRI76AiyH+GPqU4PUUpCCfHm0jlg7SiuBgLpqBf
3HJLZE/BSNYfiL5RcIsRD08srrZ/k4TNA1Py1BhQ0sZLY1b5OY6mYI3R+i6QSiBs
eUZyvOWzn8fH7ITrsM0IQwdLNJtnfFBgfi1Gv4CgxOpJ8hRBvdBKwKaeSfItDqJZ
IT4FYboCMPiOEAxuRykIrRN51yCiKSiCLQBdvTReeJAjpbWL53n6oisLi8R2s/B7
efY4A+aw1lBKiQ8C5istveEMUqxHb2nU+n9LDStG7nmteVsh40kCJjQtol6ZeE0Q
DZ4UjbjfSieEfSkCPPl+nbh9AOqBLzINCyltt33I9Twe6uw8u03UPf0qYI01x+NN
Ob/DjhC1czUiYGOS7HZz0lFmFl31Qc1uSoY8ZGxPoLYlcA2l5u+rYdoby3+IqtIa
vae/oTP4uJko47lo2x/tbgqr/IY9+mQqfyoGaW10T6sUzgAVj4nFYtUxB1aNCVot
4r9q0cbYLVe2O4A9RTBxw0SAdDFdXTdhb1xuioZ0jRk3qApp0mQxlhJlYnrNa6Cm
ail1qPYI2HiOh50ulma0FriYW+q55x3nWlb6OkOg4B9v+l+/e+vCs8ptt1KFlNnA
q4LoyAAs4wqdF7oYRPtDIFt3MnVVVRdUMlXcj0PRgQXVXMyvTWA+yPVy5X6PTAac
UpReZ8LmrspDCLhtZaIoygnXY01r5yCNTU2S3wZJ0xG1/jqgSQeKnteDhWFa+XsW
ZN6tQVmwwDBEQU1QAtGZWi/rCWkO4WriB2BqODb1JpOV08cVYW7lOJN9mboNLp/1
vWruchwrpDOdgVbUOLVoUQmPzDlMhhBX9RJh6AxsbaqJ0hhzN83CVA59WJxSakR6
mVYzjviJXIiJ7IdolA8SwFv97MNDbcncfSb8inVj2REo4+dm4lxMabI0RqhEFF3A
Jc2dlLBe2puuYYhG3wIrNoeEo/O5q8ow/2+D8oNpIh+1aAV2ELgNg/FUrYYl6Jrn
fK4NnD+pNBFok0g14CEDuT1MFiaiHN4OCT2W7lrkJXJERWOMFsxH5JFkkf1ppJbY
8g0Wz6AEZZ9tbnk3EadqmeKeioRH9WfGxiMrW3Dw3IZq51AqlqNVSANSk+zCKYc8
c5+5j5jKzD1AGVjWj1SyFpAwo038sc2S0+/MOAXd1pqgv8fnAspzYvy0PcxsXANB
GNih1uUwmvrW5FoQ/O95S/hyS1+9vFvgufVGTqbFHy24sKr2/WwJ0QajVW6CmIfU
vLuL77kkhZfEHQ/Tf42fpd1WSY8wB1Xpddt3fwo80CKJEDH3fJ6pZD7na3irNf2d
aLu2htyeSgGGKoCZ2kySpSy5n3t+bg2vAJ5cplaKuhsnUvPxJ1fDvK48qtWUH/1X
Z1vg/Ygr5pPTTw6rGAwF1v3QDNoGOE6ACHkN/YasWKygr99PHDbPtVTZ/dCVgSRr
8Srj9VDpIYC2wLHKqyeJgBEM+3WcDnWsklHcSMoFWzkqvWfB2uZNXVEzespXrGEM
O6cE5NQAJZOcFaQxB/zqH520U3Y/l2EN7cdBywntUj+ta/54T/rzqM1G7YYtnRzv
QLAYG65l+U8DSaLl7h+YGQx6GtEA7bE0ACvHyEhFPYdAQjLUipA1Cd7xfjLqRD4P
H5spjRerJdfcqOLD62o+zPDQeWQgDcPH8eHWjhCiL9xqoDNOwGNB05WEmqHbO9G+
auDxiU6r1cYLKMNx0l2T6rYBKvetzAktdJ2Dz2PMx5pYTOhznyO/VG39Uq1Sa0Mo
AMoM8pkzwLfIDoLHO3LoRsa0caV9iKFZXANTI7Ij4XB2w2nTjQ1PWSYOURhC9JlI
BEo39z5OYRLt/UgG/gtD4XG7dTCDxhyydmsDS04Ix4rj91eXPnhqpdw5CkJdGEYz
7s31/X6J+qq70mvRLAn7VIK1kIVm5ZtWYQS6RkOesBq2pVoWSJuXRcVOKcASl2wt
a7iLlnMMTm2JYF62bv4pDXZk6i+PYAf/NnE+y/T7pIVsOEv8OotjXbRuocmCgi7l
dvqldeLgXGXDGGqqDjvsCuK3vpC1/Od2oqlGQmJuy69m/r2dXtBx5Pv5CGhZvJZG
WBmnp0h9IuvzihNliWGrAU2uS72ep3ZJa7ixKeH9bIMsqfx66RuyFmTz68H6ZZGw
5E+kl+swTOZAWVI5aV321hXQ9arvoNKAUFnptZNItv17NPxHbB7gCWYXmw+UrAMJ
vVSmO8uGnS/0WYPkG9oEfVghDrYpbYIy5OQgafMWt1w1lT7VYsVOIVZX5hXfTolU
/yrnU42Gkb2gcsZeiJjEspu60Jhhpq7u4sftk9IngSyKD1D9X3PyB4AgqNL86qUo
8OxAzY1TodDB8vHoDBrDU/74Y2mBvzp7bC8CAkxZRWRpxOzltzCptVl5nTzF0gex
bT7PbylBQiU2HHaJ55m1EhAA8uELKonNdkrz/jLGHy0zGO86B3auuPRRoYgPUwVi
+zOJ6qoEdvGfMnLbqBzg6D2rbXTrhqvwBoFObENbLTlsyA2f9aFbkj4J5bAggRCe
bfUIbD5O1Wi5cKq8HXlPZphrJB4H8HTes2KmvZsrsFvyNKlgieovs2Ejl9/qRtv5
BWdcsnqXlJVQSciuHZVyYGQwfz6B0xHy2ZrHzw9M22pKlBTndlwmV5gNhBLW8qGf
34sfx/DJCbA9+IteAeM9cWKFfKrbH6KxibCLtfNJWCRMven74wqJbIFDJpIeS55w
UZWjwHyXrJPWC2dToOnsenyYOL0sAfpj2GhtIS+tsVBFSs36EMrQgaGPOylR07tG
KPqsIUrWlseevybUNMaebA5E1iN/rLeofcGs8cfBRZIguLB/46/D0ExYUZsGmUNr
t3g+TzLoJ1JsSymhcBusA7GiagEdGcA9e+gVbZ6tXtvqmNUiJ5HFjU20MfSzmVK/
bvEI0zryWJxBYwddTPuCDWsEXuAvA6UaBexDG2iPg4PgFkKQRmvSX5oukFt6l/Hs
tEpVutJ1USNeA8rUZv5+dsP5dND/88FDHUKjGLG1X3EwWzwJeQ8b5BYyzJjXU3gy
ooT4Z+Xytt6u/JwnIcBZJWXTzj4jp1jtyHTl4Hfoj73dzK2k3TatUX0qCnTYSP/s
LNTUn/mQbRBcRmJyRDALfwDpHDSqvWakljXcGFYKHUgqu0NmvQNKli/D3sL1i4b7
r1l3xnAcvIhOMv/RuKLJd6IomNx6PYZW7HvHWommsGXBc7Bs7JK09UFJRIXlFzIJ
UmRkIFDxRaVFHi328Bv3T6QuT7bOwA5xcxgO4zuX4eoaN2NhjK8NoMWLl+dfkajQ
o2Sx+pco5hUnOWZ59IoNiG34bo98h7BJPFJccG+CAkW/u5smnXRzPoqQVMBJi3dv
h/iqVulfMDrE57HwjNgs/GP0KFRG1o72uFhKkoNfT/w+ZdIy60DADk1atHGTc/9t
R6YY/PiGCx4dK1Z+8HwH/IQVjgA3tllmwNr6/J8mhtGa1fAWz0azHEEDJ5YRGEVd
q4BOY+OoemV7ulBlj5YVIPTN3XW+XhK2b33AtxlxRSKztMZcdFwp3WiLI9DVUkAd
KnPzHasyPCbop8m6MNixuduGP8Ha4UlYdqguhJgmkO2CnxPUCyb6+I9+jwTlj1Be
P6xb+C6x9vZsC93VR+wP4Wd6ZWyWVS5n7T01oDtpKe/uLye2GogQE1SRzelOhS5x
dJHku6wBI/xnC+RREdMYR5SVbRi7sBFZ3rKVaJzb+JQWGrxEEt7eC8omja6E7i0D
447+59qqqmMysKIKzm8G+YZvw/5QpA1UgstUC+n0xkDbW5+06QBLYkwuzuhqGEuH
tHlqew/echq2U64QYBPX0nddyKyZtbg+7/5iB2+uYACxOKd2lvYKfpL1Z8vyCpTc
KvmB8pgaKtHP6kwNYqQHJ9bg+RoGBKjHYdnGvjaEasvZxNT1Rn/zGu8N+1zky1TV
W3yRD7ZJZwN7c7OoYxODfx32m5ZX/EX+eGV4RHnTSw27CdDHH7rby2uYPSMZId1K
C79Y2UGfhLpASGUvLUYBw9Br1RzxdWv6BwmoeuUXSpWUtr1Dj4hRWVftWcbBUHKm
71Oaf3PgCGuzp9UFusb/vL9Utc021MZ5/yefY7/fZc/DoZLJYwHoJ3ITPhBfHfSW
5VZtQ0MGGVNuVajZk8E9ZhUi4PrmpowGlRnsNz/7npCmfXHd1ys6UdrNOqzwk6WK
qtGrkOWUkY/UosnV7pPI+dmBJynk9oUQ/zfvSW2QERl+0xyqzlQGnV1YC4LzHdF4
HNsl2NtdglCAkcP3sr8gghk4/T9jL9JD9T/MJrZdIbVvWU1wfq46ZIWJxhSnS4hT
bp4Mwa/1pDYfP/WT9BJK1AiXcEFOuq4loBLdgS6VpfpAzcQkVeC+6lR4zt8zCjLS
Zl15xSI6HPfGpXcW8pELiYFddJySaw9LvQss2VkDpXVtmJpzuRg/JAJiAf8gsNqO
lYJZTsN6PDIMKo+pE+i7LafIN3Pwa+auM1CPML5Cq+JRcPVDJ7cUEPA+ADpR9waL
86Txq8Eb5svdv2TBd1OCwCFAUJ4BL6Vsw0hZflQNeOi50SijJaKQwxN/GsnFK2t/
s9jtS6S8FZk+ENcRdoX8e8vSgMWqTrX8W9LOwYKzZWceYD9rHzQoCbmBnWy6xBCu
BVVGxL3bSO1RFnvCdG24wYnVPAEU5pHf/x/DzOgaJjed1d9VGX61tkctIn1JQYlC
5Km8x6/n2xhYo+JIGqpkBp5hWTOI+UOG3npFRUSRJRC7+0c5tmhVHVbyZGvuz3Xr
3ScB1J+c2n0xtfpQJTN0UnxL51i4sAwOd3BrL4+gPSB0Tk7iGL03++03qJxKasaS
mhuLebaNqO4hXVbjXRIY7Jnbbi/VxyTqlS2bo3PNC4SsI+1yZo5zaERv0W7Bswed
eymS6XQGN27am0IFdnKyWif2NgvW+nBnur9/Dahjh01XbkPoRuKyURqciMSQxhpT
FmDD0X2/1c5dD7BXbl9RWpovvrqBTbZ+z56N4GNsZFCQT6grWQ0J6f3PZAc0+C0m
lsjsDLPTGO/T6VzsYTb8ic16mQBqOYW96YwN2STYORbTPWMp3f8S1aRl8qw5j/WQ
GQ8y0IjQERlO6s9jIfiIW3skCTvc1Xe5V7eWT1KdK57WrTzHSJ1c3yekD7EGpZmw
/sGB+upr+Q8BJcSHasL95KVUw+al1lpigyIyRXB92DtcN6DenoC/aWtDt5UEDaZA
iVPpIqPKDMSTo2Z1sLdTynn0QMeiHO9ss+gAAmb2zUDedYr2X4wEe7LpPSEAlz5h
bz9XjBuiTMKb+7la0T8HLiEiLjX5byTRCiK+Hqm6uFrSVRr56Y7yEwwMCGsNO7Ta
RZqsTqQI4cpTpQWfMZ69L/6leoVFumiF8xsL3a7NQcwnGl3lFFRW6kRwFutbqEMS
qbcT704Gn2XCU2WJ1eTUC+niqEUArsI8fE8PBWMNzgRmcGlIrgiUlM4d28dg87dP
FTKfK5Sy+UdPinFmlQFkYdbVY3RT5JmeJX+afxW7wLfqCeWv+hQCvTcy4lhcwG7L
nJL/MzPsN5WcBc/mz4bLZD1cy3cyIwFzxp9UXMijigJI+0erCeaOJ/T84uqH9syg
NRRviKN1YGXurHYIMft/fyRvLyggVwVbQPv7m1TLLor4fbWK1ElmuQc2sTXR0PX1
ez8MZQL3uxC6sblN+6a0JIogbfHD2aXGm8l0H9dY5EpZKmDb0p4G1sUlL6T85z3V
y35tdvIRqxzIEtvNE4HtMOj2V9iaPCNQjr7NTjFpqWe47HzrKzWf1SX5XfStIW6R
Ca6mMiPhbez8Cfv4M45FCDTtS+EQ9HhUxmYkf3qU6z6d7I51sXxZBDlprxSm5suU
CiglgUFVOg6y/IuxuvxTlriQm4tyTVd6US7PEUyHIvVeuS7puvCFNpkSRAojHUlC
VYiBdPO/fuUHlwYCvrBPxIq9oK9D4va67IK9f0qZ5tKraX/V0UoMZkG7KRHFUrcL
s4X2Sq8E4wCGWN673x01pPAf/xgG6M+FBDnGpjXdR16EA19w6aWQZwNDwLlRkcot
JkZabbH/sK3fqRm+s+WmS+w0kDU9A0WsJnJEIcgkc7kuB1QuBA//e8dutAtH9cjY
gwZNCPvsDHbueUG2UCiSZKaJReeASz/BiaPBb1CD3KqPNk2laqk1Cq9yGUv05fxI
0DJhyRAyUNjFu8X+JEAVl579V2Nsw/7fRJ8VWYQwnRW8ITm+/I9SNMCAMmo15n79
oExfN4SrE1uffxcV1UaJ95DMjDamaptuxNGzV1FLxbEWGUZ37j/s1NQPZMuvvszR
G/TD+fc56+VSEzSOCNcIJs2Srvz+kLkqI3ROu/cWMHXVnO9AM1l8IHViq4SLEV35
cO6266k52PJn45+L7y3rf4BVHoYxvPzFSXmm/jXJYex/4nAFxTw9nVmYNOtxaYtu
2xHCLqB+gb/3IO/ANC+LN1Pc2K8rKaFBloQbz2TM2SBv9XYyV1O73nTsgDN7MyWW
1iRgjMlXAA5uuBENFeD/0danoOCXtKI2ieEoeWIiOhQhKMxBfSBSMuQUd7dr5Vqd
ICje6IBqMVAPPiqvJfTI9fkj1sIostXrprByi+qGdI+9SDYDjSaZoaCyvhtrIcO0
4TDXBzVatd96u/uGd0rvqzgCNv+m9Tn4ipg5rJ/OxtHv1vGmHcThyk3qt1504EA9
ZIjk1GLvD1XyACEQJjyjjURWEZSj2WLKFsAPpjR4iJRGuAzc8UwBP0GzxM3NNNH1
cYoDRUXEpqPgA7E2e3OgH05jYkLrtCia6s0P2SCb+//WDGADGmyxlOe/nkQdFOnR
45kzHmPSk9N0KTt0HYt1zGpZYfGk7BMvMNBYElGpWkdVjzwcItVArFh8glfIkrV/
IF6GN/2pI9Ts/up/31tkNg9v2t2WFE+/p5QJ9g5yrllB9dp7HQ3OFh7h39zDjr0j
dVUohjtRDkOYVGADkJlwMRgp/80gcuNhlxkAOmoIRz38q2rP67yZBZD3o4a2cd+4
kngS8wXJU/wEbzC45vNrJYsmJB4N8mfnORIelSADbECwUL+VQVBzNILf0P5Eubcc
mhPJNqxyUrXbhM04ncTCLN4CtHIwrtEjfT2+cc7Dyl9iB9ubHU9G5N0Pc2Gg0u+X
d2J25hKcVhNNXHyLkGuvaoDSHX/EC4zGOOLt+HTt1QUTq0ip8C47CaEaLDKVUsGL
H9GV8IORQLm+bFxgXGPCLnCb71GUxbnWNu0rvOF1EIs75ATnawPD0Ft0JxpD8Tk8
HX2+Bgz5z7p5CT+DhjHRrK9tAfYAcpTQUPKaXeMWvQpPGldsNeNKzNOdqGEvrm8x
48YBvX6rdRSBFiXiWr/fx+3UqGFP/Dup4CvYHo1QYeM0Evoad6SleuQicwFlP/mS
DRgFcjOAc0H5MkPTd64Ct39PtKSTSxGK4xGiZYavv2hUo/BgLYJQgkSMIaPDiLfl
I6DTUcRCvqSqO5Soe1RxBjyJyT45NQYKtWLumnZeW3VCL6r40K8Y7NzNxJymvFCW
ttZA3ey4UHH9eoB6bcGmXcpjCNvn+jFSiIi6QLwup7GCepJiMCwX5pswxdFl6Hit
6tFo+9vBzQipmfIHLKi6tcCVKaFZTzZJlYi2ytg0hls9G5jX+B8lLwaN9sZsxXzG
Zd/Dm2HD54eGGqUjX6HMq44N8ih+YVnGHoWTb4B2WbSmozpKTK5l3CxxrCRk2w60
56yKr49H3Dc01hkqC09gdSsJeh0cK+udPskHPun7o8Zj3TM9J25vvTlnxDGfovE6
q6T58r0vhrNhcPCamwsRxrmxjXypHXQhZN3zzfAKqAtfycX+zb1yk9kZhtKE77sj
KLV0SSnEaflVovbJ5VjThfU+C2La7AGgOIFdUz/j2DPcC3DZ043VUPRexbmp/qQF
tfZ1TQdVgIAfT9RDpHRaWxMMB2kHIBCmBiRMOt9IGPu39rkwElB3zpB2vK5Ez/yU
cjiA4vcNuFEHswnMnkJtDnoALnD7ztaZ1vS+qJOf8BGx6LnIYTgT1K5zfn75D/AA
t9Nn9W9Ix8r2Jb975fXINn+I6OuHQGMADTC2uXlGXFEGRehD5kz0W5emE+E+HfAc
pogvbkBLRhiXMsJO0nDWOsvFA71RUUpdpm3b+hhJjzGLgF0Bt/pDC38e9p1jjOrL
kLIeSc3n7Yq8db2j/a6pArmjPrsms3xCnyP5Pv3CUaPEQavW9YMNOo1ADl8f/BBT
6x8EmLBGmPa6pMfNC8WISKOnGTImpForsoIG9rcPdr4p/Il6Xhn7wKU4B2dVR3mK
R7lb0fN1PaH1TyLsXhwH68JpJidSrOfrRqoflWApTAXDLS7WZ5ynb/mImEeLwbWQ
Vl9ZAiXj4RgUWkNBp1HVhtvDWDnd+IQ8EQR5p3dEwZUdnTp4thLGhVZvdfJJSt8b
jEt3FfFH8JpnmZ9ezOYWnBoAY9KS1bf4O8PrZO941WG5PKSxzFUYyGycuxA7S6J5
G+sEfWWjMR2M/PExvOBh4PqcJ7pKxjQW+SFUa6Iunw6jrtdxjR/YZnuWHMOhxOP3
XR669MEmEamSdl3gCezbNrItu81J1x2am/DG6TVNPYcsevPWWxphjMnWJVR+fyBd
Q22FpW/7nBUaXCkqMP53RB3251P5+NghBOADMtX69urKxeCfJHfy0YkljDp6XFuQ
p9EBpH+FUVvYwRa+ieR8jN26bMQ/Wj3gUAUXE5kiMDhBxOeVJZOwqua2NgG11NaL
2yRGKErKp0C8Du4NPwUqFGKO94dWYR6Do4Thtout0RVhnp8vQIhPVPbDEBiG+e5l
pBBZvTT/7gI46rtqyuyjxi5GlWY6r9CMf4HcQfvUtIvy0oB/njdkTK5adN95vLr3
qaaQCqDg8yqZnpcHEJte/L/OVYtHwsGE5Duoj/oFYkIBIRoUMllFGpBIXINTZCcu
KVCGyVq8MmY+FTOqHYVrrgbQ3V77Xak90ZXUJxg8kEL0rigYQGqGzaeEtwIHurHG
eVnl5H17Xv+QgE+jhIpUh4czNManUNtKyvUBFqi2x6lcJUPB37F9rzuwIgIZ4VHC
vkixxrgzdxqlD8IZigCGv+7hPU9DFodx2vnltPOdhzaXjHCfTRhR/rxpi6PEd7uE
QezU5Zv2G0veEexauvz3oNLeaQtCBHyMJ511jHmr8S9dmXRo1XJ5FFFrxdg5Hrh3
Jdjjz6bSbcNZ8YyDIVwDrQ8Qm7EM3LawAvnUurXhPkL1bViM02Q2Ds3NOCcWlV5S
3AGiVipQpEwVpQDSF1lXP3wMOVmDK03NWsgqbbHix6xs2TO9j29G8Nt1+d0Ebtp4
XsUBn9cIZYtPQZtqn0Lu4ndmNcwszKmOvnSZUuS44viStcgZT0J4c6Vc5rAhN8iP
66WBU2emIz+XydAXNznhwtb9Un8+6jwBZIZQx3DOUGgpQtN0G/ZNgSBtQCJ6yQfd
9aRXcxqI79ukLp1nljMoerNFZWcJD4kdHARGzvMc7X+NC1WbNht4KUPx34azVTOb
b7S0cUXcy3FSTWgQqDNqt4guub6RQwYFyWJH5AuTwfpyC6F1De35UcQL1Frv0Pyj
AG/4LhGuPeJc9kydgOIjHyCUoCPUR/29ZIEC0FyE/imbunn4gYWVagB/bM3ZZmBR
LYGsyqCI1z2ljzJxvCggmNe8v5D1qBOFFgcu2zntKuDB3vm6mAQnV27ZOnVZm/5M
dPLzleZMtYb6l1BwYrCmeYqxcGom2tZ/e++g/IhyyqheZhDP66pS1Fzla0Xl/+FP
Qm/KRIA5ld/gVDW2o6cVCDpeIuzSNYr9nQDrKC8Qk3jkObUCJYK+FM4y9CB8Sp36
wHMSsFthdTgheE4npVRct/bMDemSQpSSCXtDsYj+ZsY3AKS/BnjlKTMo89oE6iaA
sGQz2xSVKC6fIJWbFYkqa3PMWdDIgUb3psIJ0ZwdtHaFnOeSjshOjMPRs10NYRZo
txgBTDjslnKdcnQlS6A/NvHswVIWvS2ANfxide5YQ4TneI6WabM/ROXP/oR9c2TJ
J21d+iUHzv2dp0lMUYNn7futiHK4bHRZlnXgSEIokDqq+aOk/E1QqsvzzD0t/NUm
NxAv4mA2k49JO4YSpY8AqCiPq+UZn2MUGqRJFg9jW5/yBltmuC90hkpbc1NPQfU2
t0P9MnKBaPVKZJELGPu1S3jwgPCgezstnQ4QRiZt4WGeCLMeZVItzxGP+jHzMAAG
IlZmFPkeWyzfvUqdDluC6qrcrmpG31RN07FZFoiVS0O2E8kosh+N/feooeEIxCMz
jkMBLOArJ7fusuR/Q5tnt423WGkz2UPKT5JMxHJvOJgUCkqn6gV35FXz3ZkGjGNe
WebIdC21ZakFgXfv89Dpcn318DEeogKuYeeZxNUQ1DW+cEJt9LQ4eQ8lyBULvXaF
GQGAc6+BfXoeo/EL/QNRc/eeSAtJqATqdQF0eT3s8utmQ5jYlaGyBB9a0z9Fs9c3
2sbl6/yX50U8hRyzRImXmypgVDS8qK4oyuCipSHAlNd9cSs3UCDp+AvGugZbI7ZE
LbZTHVHoUlnwMJogaUTSp7jq4kTJaG3vHb0SvZ1HYM7q6gzlLuXoHHm8XutbCCI1
eYg7jD3U6xopFRXLfUzoVQRxeRop0/iIAfDNN0OcH2sj2FXN4geVHq7IXmI8nr4U
2wWRNNKaARl61RokFkEBxG0Dmuy3n3qEJmKQjCQzV36Ud4MqUhJFm74XIyt0Jxo8
5S03iwhFgZ3ULK6IhMeSKrAuhwjNwplDlzCUJh4DjujqMXXAexjJho1mz4PT/Rrd
CqBBMWsMQ9INU3SLHyvqJwfVOKpTVyvXlicym9c4EkIsMss8weV7TnY8FgnFJ4Be
dpxm6rnrD5vuoeWU4jPJeWlpcqUDhwHaWNXZxGiwJdGcL1FGNE3xpFqsOHdxMpTi
Xzjzhwwg8qANLZ1RXO/9Mje6xE0KabavzWkG+G/Imf6DFSIBKzetxF8H9XADaihz
tWqZTxNatlpIKJVTbDw+j05rxjkd0hMZqSi4cQKc1cur/zGV8SEWobb2SPI5Mpg8
8GMSyn1kLWXLompKBELlRJ+nfBW5wcrEUyykJvrTY5BX206KliM0dMnKFPhNTW0F
Kb2LGIG7kcDRbgSYbKUYqEgQ5QFDaDmWN/ed1XRkMM6/mb56O4WSkgsYp395t2rm
L72+utTY9zWwIaNWBqZxxsGdW9PZzW+3F1wDHg55bahp4JybV/d/FQcufaE0CsD4
9KxItpnAt6vhftdxY9dQBcFKKmmcL+yOhr39lGiyQm+hAPh6HynGpCPBCNV3BQSe
BLCnAj6wDgw9iTCs4+UHJm8qUewJiJ07EvaOtRB0fx8r/t5a9vE8kVnxPUFh0Vvh
83TISWKrl37iwNSuuABHqjI9DT+LSBVPtupHhDeknL8GIneoY+oJS/bCYpujmF99
WC/cqSuopLboFnFZ2FxcvkmgLGKZGLZBicG5blKLpERpAawtj3GiRdhQqpR6KZBD
dodHCrT2+TMaWxw/ajhp/JI1RALNvQfqCvRhCcgzKbkcdsTlUthRLtaXC9aazfvo
kY9/IeJN5ZabGKCv1qVI/zRhYI9t6rl2JT4sO8V89dL/Skm+CUggMnSWMmph/p0x
Gm3lnLfDeIki61pcm7bPlOFMPRmDijSZadtRIDTVhJqBrL7IimVvuX5hdcmcYS3Z
ukj5YKAE7BeLE/yQWmdGE4618VRP7WjpBkHwGBJ6yM90UknuFz8jn3Qu1PJ1w5+m
m+0bAjSYO0YvMIzeu5MbEwyDksHK7DWiAGlzF/0s1uWB4f8GtVWzvbv83OmXTmyl
cLoZF7elL1gegu0fcGgxv5SHzNLaDOfLAUH0/PNz4+D3LmMQOwpk1sW2l3J+5HEj
NdDV+BAv7CyHxARruWy3L+U6W9A+aZsWxETDaaTWOzQ1OKa5wcdAm43JDDq405ri
iFG2Wjb/kqVQTtPUdGmPDNO76jqmYW5XvwU/Bzw/nz3akUu7dc8AzsWkztVV/cOE
SmmVCRGoyTRercBQFq2zNO1DdCpZprYCEK4bKHU+sEqGK2IxG1RwzNGiyw9lZ97W
nCKEFLlOFpxL8/mc/ZdKMJEWyT0QDGqp3WXso/oYyn2VwnEpVJQ4UMaS7KNBnPIh
zcINt9tAF2dKlytlhyhCPZRU7b1OSmupVf43+dqxOF3A+yCbkWc6oZ8HQaNFV0pc
8GwYdtw7Ir3o/bY4tHUB3Ia8b/F1r+RaJCpXlRbdEHVXG13F7g9/bfyjLeqbS2+i
kx2Wu3W+2ylvxZvejvliErMTQ3enIRr6HyZwcNskKZnwr4EBs0ODAN1dqgcmy7Dc
erTqrgKuXf+b2l/GW13yBE6vmfXjsVroMqE3yCAqJnLDWW5bOjFASWoygNJM81fr
EbWaOMxYQ2f1NmchXu7uEiIl8KoK77ZiXLk1rTJRI5bmN++e7/swos2F24a2h9np
QPddkbp8tVg6Fo1Qpn2DCLuY027nO94oAQ4G2fJqTi7QY8DRwd0z/VlLr4bvbyg4
6EMCpXU1rVjOe4r6+8LkwT+QVl3E7qsvwsvL1tt7jdCh2jv0nAXyumBgzLmROBxW
T6b+9SbdNJ3ajo37EMlCi6+3Z5awl3ZQ8hXbRrz8fZFn4zlvdu8Wym035L7CqWRg
ET71W0BZwxd8OcVJZvkAGAZFnjeqyT56n3JAJb3dRnTrTJZdzn+DjKJsJZkLzdk6
gZlz8JBXWweKenpPlUEJ3UMnCr5mrox+ABgwSSt2eaHbcjj06EPy5F5hPF00Ioqn
xf8MFu3/IJhl3RUcrnBkAUjCsXr6T+vVm+gtNa7Lh+knGvPY2whutTyA7d3eplZE
fN6HwlQ28xO7pUDLa6ZOpq3L2wDen/nRvaYM/gwbtuZRpKTfyKHJF07LjHvM99bI
DY0+ECiPEWdYOzAYfIII+ShDy6JgcyI7YvjZPP6BTd5QkSllDYfAgwGVTsibdBKL
toc5geCQSm6C7rdXhruP98i0Rqr3h2oBwG2q1me3PDA0TiNxNRkZia/6buQCtmfS
yQ9FTW0lYzKLScI9OA4SLiPpJFkuZWInCBzyXOuGe0P09bh0X4p8VbO6ktEcrMW/
XLljIfU1j/ZOA/6ANqDqQ4rIthqKpy80PxFQQB+7eA0UF8ZB2LSfefuvJL3BO6ev
Khi+qFIytG0iYXO/9KHaoiCNLazX3zt1wtGA1vBEE3/1bIEnEq5d6qwNGbOwGVa3
jVLjHn13WZsJhDcI77OloXWR/EFtnrg8U6OFSAtChw9meQ9L7ODj17nOuePYlVN5
K1dssJseOnQCplGcwLr9V9L5O/r2+9U+rbPkIqIDxhSptou9jFauYAOJNgBCnLEP
Y0pRIfKtax+nDui12KIsEqv8xOeUnlCRbALXTphyKJ6rvXkzqVkRqI2PAgtaG/Qx
p93Y8Tp/zpjYLhkxs3L1FGN6s8NVy+xXi/CQl+KiGuWhBxxyxLf3vEOvVYsp8kHk
JbH5wG8BCLEfEnWlfXMrC9RIZvQ22NrYSKgi6XpjIcD/bUkwhILbR6A9I++7WHt8
3dlPxj2vDvobR5A6fJ9MzUg7nkny4iwKOpB5GOoVUHVsZ4/PvYRhyF7g54N2PmON
Jz0cKA2640hFF8bx1bIQfgCCt68puMXsoV4nAKSGA6GOs6uSYPO88vbyuaqRDCPI
IrncrKoYFD1pKye8qCQsa1+F95fNFmT6j3lBWUJGErVyCwVvkbDfr3G8yFMsp+jP
A/eAo7PeqLmSRZuUVyR/GwCnnSL/mu0pjF19WnXFJDYb+YHWC5+J98hAdMSm2t6K
de8PutfjWRbHmekiA+t4MO/UXDKVou54EpKdumnUYBnOkEjm2eOgtgOfSjI+UMF6
+jQ+DwDtjR/sFTdolJFwNwW8fZ3ByphlYo4GGgDSp/7yO+D6jiL2D38WJFpKAlq2
eQMyhMAPW46HUyCtKh48OYhwftjjB7uTz4q2iXa6JMq7E1uqV0JpAWV+4Mv+nwJr
vzGXkFAGyl43I7nziXsc2XPAgdSUxN2ZnBRFjQNlMhtp05xx1pQlPFJV028MqIBU
/hkV/uKOBYUxfSY/8o/Y03kTuYsq+C/dDMBOy2Sa5Qihqu3l65AlwSnXEdgZpN3k
0bpqGKPeDvNnkypVaHNWyYV/A7eCNuYcRS6Vs/zavF8U13hpheCrAkMz622xpG4Y
N3W8x71DyMypDyBlr3WFwG2iuEQvJRt61ZwXHYocJsuLosI8v0gCQ7yng6M/HMpU
oxqsMxkFttxiUWpjREWWNHKQLMw3tnla5blx91jo7ACYugh0wCnfsCO3z4Na4dYV
MFyBG/mm59yXfPUMAuM2tQakxdrJ7mtUQ13ig3og8GP7quUth++j6K9YwsM7BWoT
ZzZVALGNd3zqS/Auu4bZYk+NdH/Y+bNVaYRJ7wiaOTaMsuu6nhNrwB2AWGOfD163
UW9eTvF8sar7QvZUZ+bFothcwzBegebOoIL6zMzOpBlpU1wFmBfuoC9kchRA+Xs7
J2qGkpU/izdRDGMUCuOsDXoVXwmkggzk9AXVVWicl4rsJua07bp8zVjJ3uvoOPXU
rYDXaf8S+xKMCZVNgscDwASI/TCy4bbjVLMIEclYvYh9MKn4/d63oY8synyllhZ6
MJyQS3JNDUJjQ4Ov87A+GC18yv1Odbt30j9RM/s7+2hXniSTgwCDvPcwxlgEF2Xz
rAKLHn+CpCtfgoWgOMPPJMZhM9mf+eWA6T1ikTuyTmG+/M294QKKjuKCFPST72DC
2hIeOFaAJRL7zRSzN4dFUBWVfvxhYmZfEvfSsIqA7ow50Dc2Y+PwTiE5EykqAfd+
MU5I9EWeKcCckMOOaNMxkLGXNB3IV46L2r1Y0UXsiQYa+APKwfNSP+ozbBRXLij4
FLCKkRl21Edh3DVNBGe5q/DLtzK9sQZou3KWiDZ9b/UQfRmW0BV2sn6TCmO6MlNS
mUc9/wBzbfEq39FDW11AtSlizdYyrTrzl5cgaN8CHCHq3AAAplz1YLxu9uib8LKU
SZfwrEWLutk1jESNHEuFujTuWIJ23+Z9/OachlZDEpHtBbPKzglYj/iPPwhtv5b/
VrLH2crCEsY4tynTOY9UyVOnMryidc3jchItrHUpYEIuZlqlrf91dhMKIN9yRAy4
FY5LaK+Gzla0SXIWSLT6Oal3bWaHNgQezyHsRXZe2wHT6gBRKJFRyPR+kEnaIxcV
zN8s9qmcSE8tLHjfAcUX3Mzf3IFHnM5zzKziA/UmDMGACuAD/DwXYpMug6WjeAxf
tTZdtRjp5QufhJ2HKS6CtiOkWz1iWy3LfzQUQOjLuQuUduumewA0TVDNUajjhl03
8S3HT1VU1Apz2IvIp05TPRYwgiFSt7wlab4OtukgKdpmP2YkjIWVi7v/rYFykVi1
S93pYJWPqdhPwRz+ldxKq53xYFRVN3eE1GvQJEv1wkX/blX2mc5WDu/5+JZU8S29
dLD/ncrTC0sOVn997grlTzdByhqPHh+xGggvzWLc4TlnGwCYxIQBo0prozPBP5KY
hE5i3ZIFWin9dhW7wqSmrdZZGUuuAYWyGxVRLfYJOPOeYhaprsGu5BxnmGoFRSHD
vqFzJNOHb+CLFsMERnZlMTAE3iu6zpAUZZp6W+BZsxovIC2X2Ve2X07QE35dtWnN
P2954Ei1n6y0Ewx+WgAgvNxsBVh4n5xp+czfsI9OYnoUcoALmuylzOfav1jEVvs/
TPDUWMxSnoGnFcsVyHqI8HaMUpCSQvIzkbTm2yglUXwM1zA7ANa8yitgW+h9t681
bUeowf4bIMnkj3/y+xXBwEEwMIh+dYPLXLKYp0n2TFx5skVKMOMx1XrB0YHwKa6c
7e3/HaIPkG/72UI5Z8DgSAklcSVrGzemVBv9dRGCjBzMktF227Tp9zL4ctb7y06z
nwa5GD9Xwsa1NSWfktoGQJvGi5OfOUIUMDTTN0XiDksxHdvbprFJ0hC4I1cNgJmN
pmi5oO1Z+4Nx9F5OjBThvjC4anNB1vVJ39jdtsc6juiVSDYfhgJplJlzsT3b4Q8g
DLYp+95LDgENa51ItWp6bioVfb4tC4Y2h2M6N+BRjALyeJTEWBF+I6BKhOFDrfqC
TkzRh198Bu+kCMOJBbZKNEl/n5VSYBpqOXdX4c+64kb17C464ypaljytxzEjG8z2
V/Zy1d49IZYR4VmxeMXqLuqOuKOdzifotfIh26wBjzCSBvHuO9PZk1JXdajvctZc
3Ml7Pn5Sgvd//8DwlDkHuxCRBaD65m9f8TFhgyJFhtUCeDg9TwHbODlj7RDIyk6p
yw3CrCHe/hLuHcvdBQmC2GaiIe+TSU8xw7El0mQR3N1ARq0HUEynp/+qE15EwH7z
t24w2PYLkHD2GTEqJMnv+cgoY9JUvGFqIUiHtDfj6atk+dl9e/np3Fvsaj83kO4E
LziIntCc6sfI2H3Y+ZO3p5g7eiBujCe8qPm2xesbCDRkE/RKSbU9J2PGd4rtrIDq
v04BI/cNy+n7cceTA7gNDHI46uhOlbPWukvWWbD1ctnedgDhqoPDlNRidXOz4fEX
Fg7EI22om+BxlZe2+HEEgp/b8Gapvx9V3QVKv5WHzzcbNcElCLqqWj9xGF9/uD03
UcKmzA+gtAdho2N0TMffLLFEET2YaIs63bP4d55Tr8jUJnRZg+arSO4/ogm+oNc6
xs4nWem8FaMAONWhhHige15tuil1vnZ+eq8no6RfHX/YIxZULk22gjWU+Hw8qiv2
YwNiZBm+O7GItiV/jQU0IuGTKaeFwNIVkM+8XeQROaB70PRqofVKVyV6EQmX/Mx5
FJOnmdMksn9jAd93NkoK5B44dI7hwxPYgsqpDBuepidMHnkhP4ZC26Qr+MEzT7n6
Kb0+iWIiDYYZ1lySVYxApffzph5SsEqfxqnUjUyJiMTrhCc50uG14560xAq6hkJr
sv4P3jMHN2iyNVCrMlSLUBNR2775wLQA5Ft8O8WoKrEdA7JSrhsd9ocsFpsrsVMk
dCY1qf3LDNo9O3ge3Y/tH2YHclcI+IP33HWBdL+kwrAA2FkGv0N/cWr6MFU1Z0zG
Pvskr74Y3/PrJKAtsSGr5z9K9IFjzK2Fwvxrce92vUdU3G2ECgXsiJLbybUaYsKg
sYFmHJWxnKxIFDfe1R67ySYQa0wExX+XlY6toCDmubXMiajOgViynl2rB280XC+x
YJVw0ppMKVPH+IPALnSvUmHVotn3NYE15TKajHhMDLolgRO0qiSSuFDQZgItxq4k
38n8FJhUt2RU4X+fd+u7Vo9UWUC8K9rVH5i3McD4A7L6lJEOYYZ8QB0EhojYoiNJ
iPClwFIx4fTHaLhxR6tGA2zIsFFLXkeRwsDWLsPz5pzPh4YCoGyC+k31ZAGwCGpK
GbkVa2DoG05+A01z2VD/xJvuI9liFahv8G3SLWHC6StTmjXl1SaRksl3IjsWhBQz
G0RiAkrjW0wLuyMRVRLEpLnHOUbiOj9N7C4P5tyAFLFqpAPWG29y2mwNSiny0ZrZ
8MHKicX6840gDq4ATOjW6XkKGtTEVhGwGYAE6XK/fFIeSGXv6V50mMAvoJCc5IDr
R7+36rqmJXW9pHJ+aBiL+mR+6m60sMPeQKC2GoCHVOpwk1sigGRuymCjSMPiLac0
W+lR6aGvipOwXLxP88wu3RTvkwM5E5/IYhxMiL1sYeYoS2zavvvIkaoSULJiGf9j
reYzGOB9cX9rTBOyHlL/52AqhQYw8yjvpB5AYC94aJS4dW+JMDzEloWaW2yjO/m9
PAtWb1DDJCBW/aOxE1wUPtWUB4HpL9tdg3HtFB81RJHWTxRChCzOk58026DBzGrx
aC6pGBCWIdUG160v++HebabWL9sVF1E+037oG6lq3lraXEoO73ik6yVApgJVTKx8
EVB8dRa3knA6mNJkSXmn8XHM6teC4VXxRO0J7O7O8Ss3i976x0LdnufaetnSnbrp
OwFmGycTGe2rZ9V08FTvOES1EYbjFkLX3CIYBv8LVUTHizpLlf+BAuUcn+cZvge7
biFopgXMomggHNtwuPA/uRTgFSIcherKRe0/q94ZuhPW/rA22YnBeCwdF4Mk1tYL
+rbq6Z5UckWbdoXj1VvsIwi/twFUwXcdB2XfT2A9mYmb9T/cemmwcLebK6KQ54nX
FvFk9ZPeckGMUp7wiryB+RUcZix78nNx7K1xH3WT3DvWuAAqSiMPTtYc2Nvqxywg
EI06toeMYd4WBXKiHhCXtYPZLCWLF6zNG5Gbqw0x1YCfasAK842nuuPhe8sGUn+1
2O4sxOpEfF+ASWNjNrwYh1mFU1aSwYA+a67WXaLUDXIX5jCeSmmhYkIo/d1cuD35
qWvocPjvUSyeDWSiBMrBeh4z/psq3MQRa4CQMrKIHcDr+CwUQfAEnw/4oM5AUrzK
mNbpkB1dl2e8MWgirsoYEBGEI507Ncr11nhVM3zoUA8fg/MKlXpAoKzp1hihQaPl
+7998o91/wWFXrIdCIhGxWsOHvwektkJCo1W74LU4R5efe3giTVUx+ohYwEIrrQW
gGZwWRZMJsyzbB1qdTKyqKDPSIDgzZE6Qtq5T9ZlNZmdEK8USlBv7kQsJ2AWITKQ
wo8yYrkaZPbErxiCLIUyL+PdId1iLMjtxjhWGZDGvaEY4rlm5Ls1lRqVQZI70qSQ
0JfSWklBCI3FBQhWG7gS9CBDgBr3o+E70bOXTeQhngANFQbSyHkuyKHOW/epUAiq
uoBcfD8Mtz0g7JSaJPEEHsDG6bMroJ+uR0WusHrBLWbaM2FCUfuyxa8UDq0ibSOG
2+taZV8bTyPSyYIjbW9M3kZml9OATheF+MEfx7SGYEFtlqB059rmDq0L/egizqB1
0Pt+3r0yg97h9lCNavWYSYiAUvI8jk7CP4IuQvFdhjRxseyJs0R/8bQoe5EC90Kb
BCti5V4iBdW04rn9hTlYBY6EYm4a9kr6K0grhHMhMphVNSkT1iuEBTz7PLpDOOiB
6KZvo7EfhC+KxMSZO+lfWl4LU28HcAsrHxEZHpKLT4EGR3GyOs57oAaFRxDsj1NC
QMmAfxdVfzQr9AYqPdGGKZQO2s0M5YhXUEKTIJuKybFXaDb7lbRqreAsy5WFj4e5
iiTtFkl0iqgEcNk5/LIYa882JP+RqtVyOW5LOjDe7cPFRdNF+03ORDoOAvR668pa
89+LqZZp/jBlZzA3tP1RhqVuY+HtMfcpYfiEn5iSOK0pKt8CkIME1bjAgyaZHbaj
3Ppg2hOSIGhhcqMoYnjwtwEwpteKca6pofyEXBrBMzG1ozJGtJCn+VwloBOMgpZ7
43cpGj3Tc9iVZ0rtjvs1ZmWTPPO5pgM7He/7GYdpG+ZbRDog++QU//JdyHIIpoYH
J7rsGCTfO82csp5UzZUrngv7Cz33Pnx3GjZPeJNgAJ4pxy9gBfUIoNHZ/AstqFXK
FFQQNotOWd+6/xfIuu/H0839IkW4H2DBsfEoCms+4lkHp+9qUUNv5RSN4fJuswHx
tqcvd14+VwV6UKG5qiGvInPEXNcfll6rg13h2PZtg8O08Qyjb1jvWnMHlGEl9v9L
XmMpWuBakN4SOvoNhyrLMApK5HK6PsM9YO803nkM2bZwqMQ+3oulbR/iuSjHA/vB
45LIUL77QkBWFqIpG32CiUpYWVfDEIxZE3Mr4tDp/zhKSMspskzAQBiif3JB6uKA
ho+rRs/fxhDWbocttYOiUGCXxdJnZy+IDfbI5+x9vUDQ8bXO89W0PdgrXH/E0He9
iF6iNQ2ImphaX5k1WNmazzCdKhINsuzQm8/WvWuosPmQLh24yt6fU0vA0GJcM5GL
e2J2HCz6VOtGkmYDrB2oF2WlbQ/3N/CwyNqMCSKZbMkLTX5ARMoJYRptm1/nPSxj
R+8eVDRwsU8ZjSQY6gO6/IUrerRxtmelu8N4rqcewEHDti2H13gYW+Kho5Tf/3dB
Cum15ti0vN6Ki4M47OWInSPwMu4cUAMTvOiqRyL/AFv2GaPUbP0EozLmmTpPpUYi
qt3S4lqNgWvXoR9bW37bi9KEXd/zyKYDXOOuGmAuPO2eCAdG362TS84z5kGaSIIW
vyUfOehimUw3adPeyfUanL0mXo7dEmqNYh/+zwy+EvALg7IJ452LaRdRtlEfueW+
XG0p/7oviukAmh5ZCKsM3vyRVjHvoRrzrkNk0P5bhj5xaj3didOWlS25gjwyMyPA
i5IuFLsnaa0fZOLeX+zNjRnxCva/m/vfdYzZCMqpvJaNFwTP8HD8DRG6pJzdimdH
ACkjXrx3rkwIbYAGgSUfnjk+NnZKr/kt775obuqrjfu8zCT26ppURkkndWvQCCWt
3xSgtqPu6dLpaHvuZ1RYR21YPk+sHizn/ZHrgMrUrcrekThoCD7ilJyS/KYqCG/r
PylbABmP27HNwGHazm1xeWJWCCnxgPmuu/dlP3/GbaxPaZchu2FaVwVo1MjUIpJ8
tF9SN74GL4li8Z/X4Ky8B8yuPPtcXyrCAHu6l+LAr3arXr9aX3lE7OubOHpbop4T
KbXER2pBcySw09S7LnQSbssKuS9x707F3cko/ayvW5CvkXhZwY9rX25KBSNh+1Mv
xmvy3kVniP0/FvTsllkFGoCH18shLQixj5EKUxFfTW0dlbkd1Ybe47OPJBZHuoip
WvJUh3VGQgbeKZEdwakpk3MFFV3ZLrJMWnjbyBWMJKju9iZIAFJqjnYAqmC1gsEO
KN4N5BOL0a/6YPC9GaBMLxfqTDAH/gYpk2KETg5CwZEAYs6fI7secGQm8QLlP+mx
G8LJveE9AA4A+/B+FXJowzgO041qUTDx5qrhdSZ/3545sn4NLRvnCo9IZzZA+R+U
zsYY1gmhDJdsv+na0tbaZCaP2bML1R8os1Uc4jqI+MWerH+zvHLITFkv3oEixpH1
5UFobbUJLhFmYzyMiOCfhB+0CvpTlDlo72Uyw5Lpc4bx1WXiz/mjNhB5cOXW8HpT
SVYcsX6XHTPpquEx8Q3DQNpAJxfs01sRc6jNqtLNpwOprgFQfiaOWJCMmhJz+9Ac
szhGy/kAZi3K0jVYsWDtTm3oZi0cE38NRxFLLlwqGX/Q06hOS3wD+XGQHJVwBG1h
WgYMArxjYp5s8tFkrmj2E6I5NJxC2Y/hcUCdDXMCO/zoK3tTMlhC/oUX5oDr2Zfl
RVYCKacZVhZBtHL54vfn4TYEUgjn590oSMHK2SEN/Jr0aQ7yq2fpMlGe0NZfKVZd
BFGkhYvZLkKLO3CJZ4n7B9QKnNyFsWY8XGEmU4dwZ4C82H6SiTDEM1lfYbcxMK4v
aqfReoBEB9c/E5NE1Nd7QgpwmMKNp2gIKw6u/EX1hj+a1D123pFlq2itFiVCj/yg
TSNcYQKpaZbP7aLYiaKDQrLn1aO9D/nvIol7xbwT4eOs4jox08jBT7CMImO+mUH2
RwIPCpaJT920NdRJNsR052PUr1ns3uN5hGl6HDBM4lBE2P2KfmmNMtthoEHG2IFP
btf5ekC1C1IOvW/HpM27VJyp8Pd1ATa0Nb+X3WTkYlmvrKkDrnqIsrBPl2CVJRsF
qG+9MyfRQHdQNSYBYpHUf04zRb6y9ToWaXEIcMKzKJzKSYKOpN2pW0Ul+Bq+1jDk
Y4SrLkYfZwB/9jNmlCggX2rwmBj84O7ZSCTQZDwNrW4QXuAteSeOkzDyXl2Wvh1L
72YwhaOLufpyJ3yp4J8n4tcZg6a3qBywG2sOlG+ag0kIgmkSK1tE8KHxLp1GCJGW
eebvSnW3yl7oXytGOOhNb+gA1HbzyFWwdxNOdKyV65eczySN6YuBIjph2GEIasao
VMoVrqGjlh3wM8rJK+gbmyEypg21nXcCcHoo8u4uGhsUbggT7cK4nv1bN2F0NM4F
xsNYFJw+vMwJVSuPoQ1pEVuZ1eByjuCQelk93lKts28xIFF++KnwIt+SkOkvKGNl
QuS7UQPwy+xEBM8uYdB/y43DxgTKm6Vbz/1OJCEBgEn5y6GfhCDhXpgeeVib+2l7
HzXOfvPnEycvm4KMJXD8/KGxbkl+zWabQ3T94PCepGkBSw+cs1CDc6pKcZoTWO96
f4g5D4LPSAZ5F25Qsasetwqn9LoouZpDIczsDqwFLX5sZ9x9jVfz+ROkT7hrLSYQ
GNRuUF0MWuFEst9+EqTrsRVSqHuOaIGvY1eEM8vzXUxB01YMoGC9c0E9uBJLyCL1
BsSG/e9nKmHmJgI43f1jZMCWZgBh2PQZ2XGZA3t9JSUdzrYLEb4sMlDne1wnG6Pz
9BVYrfxaI4OACf+y3nyk0QS3jzAbMJjPiGWav3Jr+YtySHfQDkyd67ziX2xDWp/i
yTmDgN1niggl6LqJQ6sjucu9CDoVokhIKbniX0zCVsXL2nMhTevPNwe96qXaVSYy
ZwASVkoGk1ne9RlHOg5Q3Y+UeIS4sg9ujzEsWXcPAa7DFhwH+VFj+UPkcjPcdEEV
V1o/Lw2q1UWZodu9zdck5DhYBkciCSokswKZfqdmPV/Q8QqFPOi0pVIzavzbX1IW
/fosbm8Z9R7j9E6xq5E0J4wGMKq0GlVP3+Qemkdusizj9HYCG9j0ESSepl7OdX72
uJyaTklmZu7vaOKtb8QztCpfLij70klGEpraTYCj2t2Ilr6ZoSPxZGNdY4ewahg6
Ao025J5pdltTpXkNHOdAkzqgV9SOe273rioXFj9T9OvkyKpa9UU0a2qT6k5fE8cO
sQj2t75NrrrS4X7G4FMOxCf4Y256zrmJgmRCSsRIhSmeFIHllzyWZ+8eww/e/O0W
l7K0B9WI22XHY/5x4cvyH4YZkqgeIrz5uhEBsG26pLigDznVakFoAHiaXe6IY04Y
ac4ZCUoTQnjuhxK/Z8K73hTGMg52bJFclyRd/7WdqS5G0ftnvdPUhJ9I1jHPQ9DW
fXwRTcKA+tNrkjLja8pYH7GCl6iS5R2L9v61GoaCbDicbVDW7zw2bn7IdulyW4Zw
QgYhBOzfie90ME2xOy9s5hQp0pNa5afSETXjgVUv3lRBXIt0CymQmsXisYZ3iWbp
xVt2TCyCkouR6KUl/LwKV8Hg87DLwKuQceb0rrNv4tQVZJwbX86i33AmnCIJgUAt
fxxqHr0wxUwBcmhCS7rwsPZkG1bJ2cuv1cqv1yXo0V0QVpJ01srcs4hTW56cgE0U
oTkkWB7h+chwnHJ/l23I3irWMONx8v4t18kRSqJmllMlQ65L/Eu5sRUZOfoMA6M4
wqVUaP+VISjUCPsIkU88WDBmGXHdENcCV0Nhpjeh2Pf4CtOaYaW8EXZOx/hF7MZ+
kn3GbdIelKJEWXTE/rcUvmOs77jOAZogNfh7TPqqZoUQ0Eb1YkT5S0BZPBSirwZt
JVyMWONibZxchIpIWQVi9hCy5dMyZUsefcHRXIgpqx+z8pscYB2sXNkLBqQRAbD5
5ROS2OQxXn/2tZhe1PeQ0poKWvMkYGfZdbqLOpOGregrFuS+1aPTWDlBZyP8BUy/
pNTbao1q5JhUzjPo/mwF7zRWfmFgRf4ieqb5HFnu6XdyDhrOuGKT6BOoqGpcRYFu
mG01bTRYnSBOJG4DukCSINb2rC816Ylf0Tiy7GrCUHTcGrcX3fXJ0yPdM9N53prv
yrCicB1ztyK0H456FuSMFrMDfGmQErtmFMZElwVOAoT/mM3afDwjwRntgjL2/Fc7
exqUB8/uTou3B/K+bY41P9P6xEAM9buisQ/LvAGUlj9MhpWT9ikiB/ncUAvdK3v8
nbRFER4hvbMUS0OdU2I3SwaErqziCRN2K7GibkI7CLfeSMNnSaTDeTbjb6gAJVDb
crqVG4hsGUZ6o2TuIAk+JiulH4wAx9KhGHQyyCyFGAAATuadYEGbrcylGDJOQHmj
Hv3h2CQTdtIL6ZszboNhYz/uj8whQtZVCJE8zzi6h1UK7QFP/ojOJXjXUOA/j/HC
jSOB3GFKZFs0uoZj2V6y5VBQT2aeSYC2zYTXdKd5125C6GOJ75UeupO5/nW2z2OM
C2x9s584LOemv+zDEsAe3tOBAsAfh1Td38E66QUspMQVs1iPI3+7QvtRMOPsw6sp
7Y+nWKNex27TVrUob6xGKOhFXFCBiiV8TerQjk3tCf+ckVAgR7/o73PWpsYCPIjg
rC6JL5WaEA5Pn3ZEKE1usIBouo2IX8Fbx0p2rP6EqgYGq3G1IkLazu8o3LLCcjta
xgafFlyPpss/ewV7zYLfCPgCIggdIHl59hAR8lfktYK4Z48EDCr/9omxUp7nXBGU
flIVOn2WYPVUKbdRnCBSGxewdfZ/VdV6k4ZfwcmGIw7eSumVGb38CnXmGUeOw8TJ
1ZDLM7VMLkM24pmjrZMlwzT1QUPYHvYT3oTGzi+nMuqz0RuoXAPQj8MbYxAT8l5p
acA5zVwLOOmy49oa+jaKkLtS9cCg5V1dREtZr9yay3JQNJ+1ztHvhfX/v+1hJZ6t
Ob2C4Fm8eWw9fDoxczr2TqdKK9kPqLP8dz9jhjveMnOFtAyD77iQ2ZFzvHwHkfv0
ZFvAUyEv4WS/Qc+gVLPr4lECT56vqlSwv16JQLMLGaRskzJrA7bktT3d4QyohGdR
pdQJJoECEP24Z3sTv/KKRRrs6L2QV63mljZe26PWHSUTSzz/vdYN/KO5KeAOseWI
/hYCsffiAYGt0uFvPofsduKIwHSudUdkj89TzHt10Hpkfs7cjfgT5r/QsHMc9mAg
AA8QCefxZWAOXVkta2RZfdWaRJJieDUdBQTMwgaUlsnyH0WxtUiG588QGjT49kyA
5huImX+OYVs1GpejMuoOw25NS4RCcJqR9lbwUaCaIhmrA/dPdeXCIpaTLT2pKi0j
k6UhjjBn4m0vyTPSK3Gkh7dvkPnW6Eeq9NoSzSjwE3kvEHYsBdS0FSrv9NRBqgaV
D83c/AZoXpU76mgWdQT6v5z1qgSc7vqLZdrNax6vXm6HEX5Aa+UsTSM7D052/UPm
8BokOzddsY5w8xAVhTQuUDWvuDqQcMQ6HMPBkWL7l1M1qt5ogT96/C1+pOZJhoZK
78fJhOJ+K/iCJS9MPDuR0m0264t3o4Jxdfdl/nDJAV27qMTnzwVoxwoRL0p+JITD
eo3yXPHD7a6sU4U5rpavrRQ9A4Nu3bGkEZqOH3PMtEzvc9wCtqkVWISDy2F0Q/YQ
sv2Cm1s7CguhUNG8SGncznX5UOfchKPRXRKwLPTpty6NBTzJFGhfYx9yTvFChKD9
N3BW2fZnUwPBDm2U60VIKFXd60wBXWtOiFjARUlxMpiIeXNvLYflWLD1VymW5MJw
9RksIw6VfXm/uW7uFzWc+iL7r27P8sx/oVF/bF+Dmm/AggVR2PUQV/DKjBl/SGSs
Luzg96Xh+ejmRvYrwcACPm5IP1w1L8GZlB92/q0FSb7zFBifPczvK1JVKv/2Z5kx
F91MDR5G+8Ov2XPnnim65oHqHtIC0fkrZ2yuidD7yydtqJ2OZiEKHvKI+GjExTBA
BpvEDLdXsnzPsnQuuJxgl7csNKpsA3vvhhlTYLFsRmNzvoxG7QKnYHxaHPzx8f8i
s7/pUFZS6WqKGyXETN1pR+9CnWpc6ykEoKe+bi+IudN6b6+7xeAzBOHryU9lzD+S
FuZkGS78lCmzHeWcV18vp3qsHbAyoYEuiKeqTezMb/9SdWdKq5WMU448hUqSQZmM
a0TOs7wKZ6J/2VWLR0C1UdTuaclScg2xGzNC1E+YVxru+e2ou76lPSb4kup5j9vQ
T/18I/N8MQCa5KSGSn4pSby0La9wlo4O2EgkGxdHMSCQ87wmfnPtJqVOsH3cMAI6
LlvufQ9/vIljIeK4U903emdnXy7e/ziP99bqenung4wLvHYiQnb7oiU+fMPVJVqv
uK1anr39hRi2Xz2keFN3ZRmmz5gz1VmjZIJTWx0WWLm3cbEckitemyNrheCChrXU
wwNNCDSd8M7yUy87evPnI/AUeYFVXNNQb6iME6TQQLkDrndVwkzeUAw6V8QebKCH
ngQycoWiX83OJinDNu5Twk52YGuBJ9PeCGzldh2icxOUpXV+eEMEaQsA5xoL4P7z
CqPPCTB7xoQfit9kodOryQHtshdBMuW8/DH+p0NkUbcwKMW9n/8rlmTCe6egjR/j
DW4vSPtAAcB0sJE/+r6xEFkAtu5vOdttioAlasMZmwFrbo2PhS6zhdXEjJzztH3H
Gh7xPjjOB/rpghUY5vNhtOMFKlbiUxFvLLiGYVGEU5BNBok3KGGjRhI2rlAupME4
NNQOHIE7PggqQHa3IjxLQrviwfDReeZy83cY0PldXXr1/gSCI+2ggUTLr8fZs3Zu
ntV5VLnNw0JE+eiFLBEK2vPucmfZDMmO9Px46lo+6qnBa8IIRMtO5muQkpX5Hw1r
TLWMiofPdvCsC+0c8BCnqUqyhkltjsXOhJK+ojbsLZe31uJhcAptklg38phqb9oF
aI4TJVdneCNEwatpodKfd9B0QxOkQJfYQRzKYNkhznxsMdM7qHBVXTfozxSlGCZT
7xjnh6clQZ0ItS2+Rs2XZFQihr710bFvDB0ONITLLb1Pk2/KSNvJ4KFe/D5dWpua
cgCS0MpZFcvtgRoiyo4GBORWeRSFfmaMA2LsCgE9jiKdf1/HQSGWqf80rBD6esNm
U7tiI8u1gtkAm0GvTR31yciLSZId7AH9v+TO9wIV5SmZgQ5DX5sglbrupeZHX7eL
geWtoIJPD7tXrjNQs41PMdhYc6+7WX7PXI+p7eQtc3t24O4JFknRmzIRFxqNqF39
AIoUXbi7I6Y4njnhSOTws+iZOB/Y7D+9QwK+gLaFl1VN9HvIjrATgJxZCF2bG62I
MlHjUNz7L/xfARq7c0n2ZRa1+0F7XgxTbQV/UH4yhKainXDTt4E39YbSkdNUy+OL
NqoUdVJXRJbjuv52krW/g3U6yxC6LpY6MmtgTNqLR+pNoUwDELTKXI2Eke1VQzyF
h/0V9JQzyvVKKVMWK8x+EjqOzcLciiFf2XG05gKtLD1NhxAUKilxKnb33SBWgV/l
lO49VF/9O1xBfe+Upbn+Z3GXnDHisR8jNN/XAsvhXofJaEpCvx7CuDzXCqU2lVH0
XTD4aGamUFRi1t1gbiWvu79Oi7DhOndLodmRXvJpXKCkJUzlyI4cEGpmFSBDyrgk
xoLJo/zOvSOih4QHCAXu0w44tRH0YNIg6EA+l2P+HLY2qMTIVPBXZbvBfS0OQ/pm
PtwnS3DKqsFXOSEL6y7yQNvBN3DDJphtHiaMs+nUpywqA2X08WozsHAuzy3rZOmo
SwH98e5lIRWgDEjP2JjqP3kV0fSFDMhYx0IOUc32z4I/tzAywcWDoz+9YulU8nMJ
ztDBRkKL09hKQfOSnbyz/dmaNn/jKkXxKpgBmXIxxVDgb1BdkLLRHFjPW/6gkNlu
CyFKK+bDhHVrUGsAWDugN/A4vveYGuldqxCCiI6PQYzeP7MQYeT63bZ5JC8Cg5kU
37oQ8z/8rESUzUP0qFNGtDA0Z7oz9ifOb9RcpKkVj6bGV1HyTrFNQTz/cSJAMLXe
eqKqLgp8MPmVSS73aOxKgnFGG04lrEyqq5uS5z7XH44lqoUXtgWhlaI00O4kxsjb
cpJfrRLwcWq3Hbnf+vaHGfREjMWjq371giPLZcGwhJQ3Pa+fMg44vOTa/8Ve5x4L
3yjiJGxpItan+nFFWD4ycHKVmyvaIuBlJiNg36LPWFsIms8SFzJ/rF/FIf92jv6U
fb5M6S8X8Eon5WVXlJo+nxihjwRjGhBF3az2w3gztAaPEk6b+8q33/UqEMt4riFs
uWyQrj4J0J+XWhxCm+36fIZY5Kw6ZZJvNFTV5FZNmGlI0YjbXac4wHQAd8xo2w3I
pN1/dkPRm4Kdjvu9PdYQKiJe7f1oju3TZ6bsdFZg2kd8pP25B7RkMaQcn7sXf9Fv
w10go42xxZetdrOt/WrGHEKpL11+6SqZolLSyyaFkAwmIz7AgMib54zAAkNpRov1
+MR9ynD+zp2LoOCtb41tPiab+smKZkdSBeQzV1bSI7Zb42bZx/AyvdGxmcCV6U5A
g13NXeX3gfldoVSYinYe01+WVkiuXHnFQkP5FDvgldUnALWaWZygnKklht2l+Fpz
S5+eIMwJlBwiAo5wlkDPH2G5ci0b595/ODaogbNGcu0sjzmiPqkGLaanbPUuBhe9
8VwMSCs9P90FaqcfNvDqrfrcLnVXGC6sIT8z/aaMNUEzPrxHDOV5lUk6ajGD8aRG
PAhJFj0K2ovsa6gVQW5Vo/0KU0xWTaOr8OlRu0W/hcGZ/kgraIGGE9++3C4QocZ8
OoHp3Cb8Clbq5l7zlTxXbq53SfUuIhVcTj47O5OE1NCgymyu8EgzImnY0x63xAdl
du/Es8bsI96Asws9svgqb7nphrHOvS3u6pFA4Q6c1zyWAa2CSmDuMBGJI6ZDgrHM
ww4A7Md05/QgQOU0w0wfp7G+P9YQ3amB5qFAiwBJbL29yRPe2Cr25Y2OpCzZrkLl
FmKt5y/eFx8j5MJOb4xJvasWWwJFY5wxCFW7dJCVF0JkRYRvBFRlOD5vl4VFMHFM
TnfpZHHtCBFnXkxOBpEamkp+1a90dv6BMfD0S4Hp7rVl0v1iQuWiM5vm7N7IGXgT
zx52k/jo6YRO+NZWAkQqz9rTHx7B/6Z9I3IVKJDtg3c8i3Odof5W+KOzGPkySxJc
KW6u62oZ5Wk9Pz65jH3IoLS2FeV+7n2aQIkTIrvGSiup3ZTF+Yvq3g8SUvKr6FgZ
1KPSUDKIlu5E0lGEsU258IawKQzOgggeQa8F0IVvn4kD357EQF9BvjavO5yADMW1
aaEYUkANjVBmae0i7Dftyl16gR4e3rdiXGCKPYTywH5T91pCsKfG62AtXffGOL0P
n6lj3rRDV+9e/PFeIMhouYDNLD8ptk61y2D2R3ElLN4S49Fkgc9LKCWbHlN+jPY7
GbNDMUJLZoMZIgHPWJ2lWaGVKSsehyfEC/RxArl7r9vPBDcZeku9ctDNOEZwUMGC
pasqDQFknRH00AGYjzyp+05YXzpFkBzLR+gD+QZe0RiMJY0RnCRT9fHKqLog0/ep
AwrSt/ZswIXAgKwuDfAsAehmJykUHO7AZPLk/xSt16T8X8InopJEaxwzat66L8yo
VScvDsS+KxxbCYvT6Ht9pm3FLuqkp9mJa67pZnvWr4pnXknmIHbasQMKgaiJ0qwV
R8urFeP3m1GVJUrAcy9xgoavTq2P3KcrUrIAIwK4s8PxUbJiaYqwOVtBVa2A8sHW
59biQeaICxkx81AevxOqa7LP16xb1WQK8LQOW7VWVv/Z5aADSyKb28OEn2BgWz9a
aiOqlZNrd99WLP/tRhOio/eQpwnuCWnfUDJRq3ZcSWV9eE8yH8FsuWHIkPO1iezx
HI5/cH+CU/0/2SriNUblA7WCiBMni/mlaQqi4Yf2w5C6ZXaKewDI0GZg43yEcKIw
ST69AXOcAytuVURfkMGPF/PZZXdS/7VDT+l8MSiBJC0XJqEgDgzJr+vPKNChgGEs
ukPvw9gA57TB66a42RBU1Uqfg1gXyHOurXYJJXEskas8oeMlPKaWoOn/3LJCXoQ8
HQJm/StA1V001nOEGJ+DwmmXN8Mtd0dSUbf/LEt7AfPBTAcBjXvdbfkiWslykjC/
uqPHtLrpVDFREMFa44GSThhmR4D7WqYCG1PgT3clcnsYnG3NCDA1ywAfOa6PVXex
jKXvVWcuGrzAGPJuMpmSqjf6Z73JUwbMhxeooXEyRs42O+p/FqKRIGxfrjsyPZH/
jVFJHlvqfkzH+Sj3I6aWy0CUPo3pblZYkxGy79GHRvgX3gohPxKg+yMJjpawr94u
dca0ht45OoT5I0CyKIXYBrF+X+v+z+9HzGL3n6c7LAQaQFZZG/ydXlMGqnwFplXk
SDwMnfI9lOgD7y/RBZZ/VtAh1FfZQmqAEBTCsdq6czKnsfAvp4MTwUdy0gEMmlnF
B3XhksXUU+fdnwQ4sEtpmhU7pFgwiXU/Yrrh2lO6I7AM/L2ZdQwXzuhS2Ymj5Yn9
YYwH9qUzElB1n/4F2cAlGVzfTxw92U8E7ko7K1hEAssO5FTNPfXVezIs4n/4mZ3U
6V6ntz1IU21jte7X6wdYmHKFh/ZLrN5gX5mEdwXXjQXZzSRDC6gc90zTCwlNFy/K
5mW/VI8AkMyLkXUdNOCIbVkh2ytlXaGhRGXYk2sDsbTxHF8ZGQxlItlNBuD4uFG+
RL68LtnX0TzW3JOTICsGEb1ly743A7s1SVfXtHzNCobMdOnbn54cDaDYXghjbpFm
pTq0JQNxW2+7cM9eOSJIXENxFhv8G4uRRetG8G1j+dMnORIor4jeJ1RmsXHZPq47
vuKMGf/2L9pkNqWiVf1vkWMWF/3OZCWZbPSW8vQLye3Pq0A8mAdS0Y3ILCetE4d2
rc1r7bejZkDZyNC5iHFFv4KsMV5HrWII4EiWS58P1V00THj8+uRUqHSIoGd5yTVW
nkhOVGbkFejFiUL8v+zWX0dw1HoozdX0eFc8S43XBwfULdrKf9OsF5Fj+BtRLHIc
FzKv6Sq0gciob42NGRUB/hbIk/tz1Oey+EqkQnmivV5EQDO1+2bs8vTp0MGZkPj8
2EWwkbIY9iGvmFUiMyuxUT75MI6PGhCkS3tOUqYc5799hnVHAT9YVhxYDdMNOZSZ
JdfJ8qo3F3xLdrJxmTmfkW80wR+/oreWbFyfVp/6TC1wwECorqDZUczi/RNfEVT8
g3QOJZOSL9Nxu0inso7vmlIFyw9oiNw6+b/wsuNMrowsQWcou9fpmUG//5sM5m02
XtdfPYyw4Ts2LK3EdfpAPVK8EKfQDn9G9uMQiqyQil2UF/3uV2ZUq4Dfu5pKBWL1
YR7Niy2wKl1F4eAucm0fDHIft6VGlY1mBNekE3zEdTTDcFA1VQbyrikl6dok52tr
MZhta+/0OxVDRvASmUPlGo0nUYlCbTZaiQcMNp0ipi82XMc1ER2Ahlr6fzcbPAxR
0fsjFn5MejEovDYRDVenhNPVIbgpt+LU3r0/heTYUtG/grjc2gB0KGYuzQGqCoYN
8NgM8aP/ldpqMJVIAX8ESVJ9krlNVrNcNP1/yUhuQS7zC4iEWDX4Fp9zq/nICxPQ
gaAV9QDLa9HeJEpoH5yQL+6Or7BVWb7bYDPlqCPDdtLvxxwlocxAYOCxSCz+qqvJ
lt7VH4a6d1We66AmYF+gM2yZQnI7fnrtoLQUnz2r0xdiAaBo5bIffpJ4kvrBGRkA
Zs8dEBowA7qZ3SwzLSe3piS6+QDfQ5m+7+uzyjv7c5aJAKLPZt0YTOIUxJDysq38
wHmyK9lptcmbFEP0uutwvXGeef3KAFyEe27O/H75wwdNWcAHXuOh4+2BTwfYzoKE
3XH3jCvjQq2lJvlTmDGFzkEinV7MYc0NQysCA/gqNbZERh29gpgWuGw2+oUmFaYC
yrqG+HiT9kvJ6UCVlKR6GND9MNzGxnJSIPyIyKhNYXhqsAb4qPAJ3O1CLMeKhf8g
BArTksmYv8CZmK41BHRc8zd+mjDwur0A0BJ4K/p0aWoqFb8wWlnjckVWa0Z458iA
2JNLiGtZ7mox+fJVLnGGF0SPaC8xEUKE7uB28WkJBGpKFpxizuvrnqPFqXvY6u/J
qgoDBhXtmPDZlPn77QHRVZZAQoRbpOtaYeiwZr8U+m4uUHQbuUPeuF6edMjQZ3PT
T0ihVJZND8PvKJeOkK33/dQRjHKAhK0caq+5NA4CCFvpWOei42nUs26DDAQLJRCY
m/SSam9cwwVfnwwOHJQlXVM1OItm2WiSK7RAbaSLatK+PimuW1YqZsQvC7oJg0x/
GvyExjLp7dF1iDhitXCqNjKMN4cm/WXHR+kbY34toVsu/Abk91/dFotVHKiufLr1
NVsYzJ1EQKdZuZ2SujYAqRl2bXTsPFWJ+/gKUCC5e4TRvJTuPjF3xM5vq9wbNkP/
GayGOst3TlTF3y7EdiLsjjv0KxjNzTtxkK0F4Bwizs4IHtS9I0c5UJmxdkjhIpVu
bCAfF8moW/F0ZSuUkAYYONRMEUz4D9VfG5UrTkJ80kkvszmEEvFZW8Ty++8cz7hV
YPbTrRMdTsm55IbcGQF3y+CCX46AwfMplcutJLTlYlljIqFpskhL7kQ4OHVAgQeJ
aDkgM6Ttp2lxkArb7HIEl/K4grYCmsiIMO83Bwe3R7u0AjfDM7anpJ82XJDP1Qiq
p+5WpilEZuU4JHk0VQ/Xu+vCxXWkOwPGqDsSmZ8tPRo7bTIFcNzGcboBvFSm/6q4
0QHQ66aHbui2IdRYaOEqbO5oVY2EwQ+sb8KcRKyVTk6DSuw2SJ8sdJ9eXU8Lt6vS
VM2pEhf6hq/7dQLTkAI8HSDzJVxVRjlGwX7DqVY6NpTwizQ1u2p1FAlSdvC1o2lm
u6TRBBfm0ahiIAvDpY9fmVY/VmZOq/CJ5O4/KOYFMbqnVMjrlX4APXDj3VasgErc
qRwCYfOj+f7HXIv9X7thnPfi7aESlAWe2dtX3QCOVan7QcA7Zur/CwwsgIYh83mw
8yrPS92FtEYntl0lE7OEQ/ZNnbMeIeTTabSKbwP23aJKBqPQLVYv7J5EaPiNgSbe
ldoTecCv5gpFBqcliRg4SiloQJvg00u9jmWJjrvq2vDsqCQEIT30pAFi9wdOtJmo
OOCHEQgSckbMao0nY4Z4Q8iGen1VUYnNdN7xJBEc1OySaCBwzZiPvAMDzR57Dgw8
Uy3PPK0BJ/z3/wUhyFAotxDxIa8n0v01MDccQ0YjdQdUJe3KtB0P4QHlOWwuaiCT
nmVDWRpiXVVYvNplSH6/NLTJ6wgsFCvbsdXLNqJEiUbWYHvvgbsGuwc3+doqI61k
ZocUFRXvQhKov56qs98WapE5lUi7WnRhnDxa09qIIeCb+lrlLUewQ9N1eXzEljRp
jWHCO+Vc5KvkWyhnBdDuQf/qhtSPRzbkzhKLG3e6E2aiDsJUCHixtPH9QaSdTadC
eIEjDZeRaGL2btdcYk2D2bcr1IlNmcEsiWYbId1MC3JIxMVeMpg8m3lqdGdrv9OB
e1iO3nGw1S4d1yVE8Z5BZomeT/8XjDD0+qPaoVEUGvElzHbus28BobW+gogCC9IO
Jx+gZOyDEprwhntxVvjR3fnVqKZos8dWf9BaDh4hvn279Wq3Mto3zkwIkcRhWXxa
xK6X2gRvgfgfJqQOedDXZdauWWKE4Bw6w9UYnyD4c2U1tbE3y4uDK1sMIBG1iQ4J
7/vKftaCx2WXQBaDew1c8TWGGouBYFy03iNozXPic/oRDfozdxjQWey2YwRGBi9s
QEX3a1rZWZ7rwf9Itprzl4ALo9XSOyRg5kF10qhISK2kuMpmfqdt9phZ2rZtUMKo
FnulJMcguLmQfTOD9JwN6xKAtAUnH87MCkcds1ol7+sHuUs8GH+rVjY4HOKGS0Ji
PP7aczlT2f+ZOGH1B/iYLXAY0GR0pUZZCvbdO+kwpz/g0Bz7J4UC+mEkGpHeYLlG
9RzRnGSA6jO9XLsiPKxrzrNKfEtgLhu4d4mSOGdlhgiIi9fsHf7exwQPzg/Z+X4A
7bsvD7OXTbBX3Rga2e7Qaa0/hte2Ybu9NaMN9Gaa67skTYLsSQJSiTK9IOc/R/0o
PFoOZXD/wcP4MTrsHDuQutjzn1nmEwHvOUg9kQhpz5I5rZyKNnxUDYgg6b0k7oDq
EGlQZPS0HBut/REDdbcMXnxZLwutJN7urGyIRyxnySAqrXWKCQVIzcdM6x4kUIG1
AlQnp9fJ9GLo6UdVve3uwTueuzTvjLx579bNpoj+CChvmv2J3vdn2v4qG6xzoQzc
cmKFEpfFmNPqTphaHXcbX2xjCHzfUm6OyiAfue9mEDp5qW233S8rAF876FLpHkaJ
H6kAUjlcRWvYDPWyDyvnY9S9zqcMXD1M9OBaT1vnGaEfwgJ4FFXMULn+wK1ouu5i
A105/Mo0YSs9onX4lPUPA/iIJbRPqzsEJjPDnyr/Zh25YdT2j0xK57JyVpuyhD5u
IVboMlCLJVL6XT3jqW3vY+0WvF3rcK/5RRHMWupQ2aQkdvW4BSW/pZ8MLhmzJX2g
I83aGzr8w64Yje0lePmmXaofLJMUxW7HKK01W7S+fbT4w3OF6bP7atH1QWac+WFX
ssxcxSxNMS4vvSEK39IVYu4SIwboWLVWlPQX23dxcWnRwVrLxq+tcvLKkX7StSyC
Pcp6/QXaND1MNTXtnecL2Wg/iyWDsDIJVQBMKCoXfmEU5C+GdWRXitaJuX4z2v8X
XvVO5nTQmb+F/nVuBw4KxGnZZLw5eVLiiWlMkfDxbiwytYflXbp86keAwcnOB7cB
5oHzfAjuSPsbWXVLU8eQNQCQ0Mfhx0rElyukSEYpUFt40Jwi/hS2IvPHlVYDEtzS
7bDO4O1PfW+IWB/Jtl/YHGNQuSgMaIlMw3atUNjXT1AJVkCfmPNbYLaFswVAeW/q
h9+XI4R0mcXwW+khWjuTg3k0BCjvjf6CpBw7d9yQ6EkCMgohfgwsyXJDTWg/HkAc
cLpXZTE3lIXu+owzgJ+RzvVk04DEOxTJlhncdiqst9NHgbgbN6YNcxJ1efLfvOYA
2I6nGqA2RixJNzsXUT6znJ5Kqqai5Q5u7kIVNLgpPbqYvSJLiKvK1LEYgJ0BBHVW
t/Y5qc/G8YSmsO703QEQpghOWlVM08YJ8xF21UNq0SYaqJNYq+9UXM4+38s+Af+9
0BaHpYkJZic/WlYAROcSkejudkmfEJUEYclf8dHwEkc5dQVTNDgtE9TpPNFbhW5n
NCZUL3DeRKbpwjLSrW2rC4+/xfYKVU196h0QikXPX8pN1tfzuvR/tl6E71P81Wlw
RJZuAyuHyT02Ym7Fivzelpm6KDtt3DDIqRsXPyMql5kD+rSWy9JzhwLExLzoJFA5
vslOt9cYS/y8CCpshWb2ioGHEubcQOvIVxHCw9IZvnunQqttUN2Vq4nahfIjYPEk
wRZFhcFmmXJv6azOnQjiYkGixbbzTxQpk0bUtPHKG1viHkQFSZbVLjBYS0L/z7MA
Y+RJ7s4AOuECZCQ8Uc3hEfxf5gLpE59rUQFVt6ex8lrLaUTAQPNaNh5oCenzIixQ
3GAajjC0phg1L8xsCyAzOSkMDCRp9lRFW54++xGLXqPYMRc/LAzPuGmIedWuBnkV
SCt7bYFUorTYiVb4/Z8k5u00W2sHFaxB1IEOunRcxksbhkqcScqcfLplNUjdaUG4
ZsCLy9HHnrMmHpP6sEYENAjY6MzGgkP/BkuAWM5ILEhhHw0Cadp7Z+lmYIbxoY7V
gwqSeYT/yh6turtL3NJiIoRkN0o7PZJbEZZXIoiHGmJlZ1ZseBIScKqWXUpWrOQ3
TCl1vNubVr8FWTUN0O6g0ObnWbFzAgtoUl4xzDsybq9QuYD6zWvlKHPESK6vdbGQ
tub6/ITTk2F7tDFrWH1r/BrrnsHCXZRjWCuWoRW+pu0xFuyUw2INOEccSfUkcNZt
07igKe/qUbJlqjSbUxgBXlOEhTAnsvSBBJmL4+/aUT/smuwsfRVQz8HVyiJ1ukRW
N3i6RkHL/Lxq5PpIrlz9YEsVj0xtC4YJIbxlsUu8+4ZNBbb0XX5xzGCc8lVD0elx
NWjzUU8lngsrqx0rqba6geDxyscLcysXqCtmYqbuKNOVlT68PRJ9t21yb0gs9Eks
P+vW6mzqrY0qXASN4DnPaEnQRjRynkgwlPtUqWLqnKuvm/w+80vijE9QbVyWFSqS
3lSc2Yf4KCFj6eEXC+OWem30l7Qss+kwA9dZ8CDyy89hYOzZmzbFhzA/J4X5k05N
qtgO3RyOAJBFNlIW3C+2UbLk/alQODILwZ5h/QQK1Rdv0TqjydRYhmOj51fW1/9/
IkfhamgMvFjWuJ7PkHtiNuJ10iYPRHGvPI6M8yfNJcYSBap8lxEFbYLkepmoYxoW
uFGy3PXLlwn2lJr69R8OIFLMjDfjzxvxFfJ1pJByi81epXFbW8y/X0PFMdCvbnju
Lz00mPQ7X3ljJmMSN5KdGSlcpbPot9x60RwWmsk1q4SX1yzWBS37ZR7NV3Osagta
/4KGqVq4qjP+gAhHsG3lLaREvl6AwcYQqiJdj8FUbovnFvafMLBrCg1fv98wcv80
8cfy5DjYc1amJ8FW3FOAeNxn6p8AzT7HuqEPk4XBsRWNAzGMGBtjVTBvXfigQ/3F
4q5K96voUF6anUBJ78s+AxEC4VMb8x80LPFxYvV5JxRRzvgZFPrCv4xOuE3Tif3J
jNRYYAzZAkiW5VTstr6lX/cwDMOUptqFYW9tyIFUJpD5bER3kxsFRkInVwcrjYZd
JwRtxFe4j/MwhcobwtSFcZ+uSnDIbZxGkLL6rMmgXrA9tv0lMB0I+D2xJd13UVus
FGnsnStQvIQUjOVQLulGY/wEV8T5T1YZTaifeP0rdZ1C15lDYEYL3i0UVQg+ui6l
k4XMLaCHA/CBS1KM5ZfHfim59U9cG2ilwsbh2c4eMZkyjX3/uvjk1EpYmTJjDemW
vNHU7lcdS2d1fqU2MW7KLJ2rhRhgMzeeSjqD0UY2/TtowLuFETiSF8s2azaU9uMZ
sDJP1VZOwfkde1KIvUFgpMfGrr7YyjDir0gh2NyB2LWSNXITl8U9MBFnr6txU+68
4CBTWkuyAsmdmWdiu1YlUoa1kgjnq7OEeFuqfrfEyUfVTuNpPBefBeUVkALYXNk8
TVNdcazHKgImCjluy0H3LXxpQJG9/JTxdkmDkSAQ5+uZuZGhfaEoWlznDA7pjiZ/
ZllmfjyTKPl1WGS5Ba8BOO1rEv8sti4ElDY1TUUYnwOBMLDpdi0m+eY+VYDAhB00
tYRyL0R682BE1L10ORq4+tQfXJSyGlnqsdjb1qZVhK0aBoSLOoaGb6ItucuzeK6K
JlM+1FeLDpprFVG1da5i8iI+icricIErgPHxmscyEhSh9DcA1+UAA1VlRT6kQ8oT
CwOWZ6CCwwJmuCqmEXwHcPLIgM626iYw2k3WLh02tKcizYvGl/k92lEALb+S/9si
QpX5fpVaalTWaB19CpgBCPDJV2NbhKdu7vaxCPtVjZgu4QzCLcvajZJ0OC/zuomy
cJeqsnw06tRl7tuhJBAqXDO5cL++9lhOoFriZyJSDktNSAVGWz0X/XKFpE28373m
QpKOIczRloKJ/pOiR/KX/eUMzrFVlKcVTqqrzXhNJysdSUlgCfLYQnHMvVajOhkK
tmNNf/50MUvZRtSIBBoKXnCnnE+VngsiRROPxg/doeTlY7qRNbQ3S/wJ+ur6MLcX
7BPWYrpasfBHQR+00kECWuolMGoFVqSfEZbZZRJB6KLSAVEzTbR8OHe9MQ18+bHA
IBR0159miMY61+5NiMvdZ617hVNXa/SIKp9uXlRou9hNdO3psqOxAjpDBzD5j7na
euw7/bbc21OMJrb9NwTNq39NuM8CepfXD9Ru/4t7SKQ+xpebyNfSVAZiGNcVwW42
1zjsI591YPCK6BqPwgEogO2qpuPSYd1QntRSNWVfo8d7nK2QY9fBouCoaDLP5CNq
SQ7a+CFsJsaC+9+pethNsWg9/JNhyt9cpJaYlRAZtRS5xLYrrW9Na7maNfxBRQe4
Se9ZNhSaCYsY7WT1gl2EYEODPmNAJrVSfDENQVx4Cyp7OH9ABzIuVqnjXED0ld5/
pU2I0Mfm5DX7Yw6DyFj2iNub7WGEGGCNezPpM02n6MjPlIbpj4uMnKGJMNoMvLLt
wfArZ7XYXyoBxM4Xj9Og+O9hlj9smKY9PHxnAM7cwbsq05uvexzmR95cUPid8z5K
S8xrTGx1G8Pag8EnCTNTwTBunIP31iu/6WzW2xv6+HbUuiZrJDCRBvuVQWLGd9/K
refVl4zp1duDJ/2s4PvzhRm7DCUvD5TJxbqogzHXUYinvFcTIhWDdkIQjdv4HarQ
Gg4t3xyb+PTiDmNXpGTb9nfPfcoS4iBkU8HJe26EZpaDUA+kcRGv2OjT5wU9PF3E
hNGf96ZVhW9VyvjXLbs7YwDV68Zimka/OLdNBmvgnpofAVd2W80fhxMXhfcQ9Igg
u4Bap1kEypSciIn9xXYvSFeiJ3O3YLaIU3BXwvRmhd+PAu3N9B1slKuhTvxq6AA5
v4qrn9pXm9Zx3O+JqIVPMyos7PMjw/mdl6sqGwaRdOHIp5PAXLPN3qpnjBbx2dx+
wGKPrKAz34POS7rAV8VuTVbSf48agxKj/zILq/1/8yoQHkTvafvJkKNi3smzU41a
U1/AtAMg10cVbGGcvVyxbLfthUK4Xt7VnYo52imljjOCR2/urTUh49qrgROYOAZ1
SWKEE/gH8MS4kGya6MgC9v9pcyGQoVV4u/PVwl1SN6chnc59dfY6sQ6DvxYfhELC
gjjG3e2XQUg77j19QPeI56AohlZEdwpKu8ycJ3eBzOr64WTnyDKl8hURNf1W9MeC
bBRg1XE3lHgxYoeyP5guBggEFVJqKvYFNXw2VLqXPd7SXIF2LFv8GfbCGWk5T1P9
WpW91NgQvBMTL5qBzP2BlF+ecdzpAXTCkF4Ur7hsCImzu06YDsd/MPxs4hySIp6n
Jt2KiQHX/fQY722mgkoMORHAoT07BhQKrnycGD33RmBKZf1hhE5eJhy4Cc7SNaU9
hX59/G5yftQz2XvpipOLMKR278TxzKuc+WWOuIG+AiO+9GOGrC7nKueinzdMNC5D
NxlByOABkCEUsX0piQFjIt8saRQhSTqDQDja93pn81UUjXdwxW0IOteAmWZKXTIW
5yMTrGbUtlA1f/NLArYYIOO9tkOb9b6NWaZxBarjzRG70M38hlSemMpteAaXyTDn
kNR9rr0Knn+dPp+rUdKWWPoajM2e75mLy1XRz5O6Dm8rd/XrpLvlWE8ueBd8dQPU
Eg1K6mrk0AlUbtNCq22gFgORLvLIOWwdrwyU4nTYD/nv+fIc5JzrXSKguMDkbtlu
V6AdioMYvL5jyJeBfGQDhHHNHi49YBMB9rL4g7i4BCiLdyCzifzDxN3Z8Js3TKG3
JGPaUJVtM30o9ZMO3u8eALhejLvqVzCJ6bAj6/Pdcl9JYQdkbjpLUxwqpvNEn45I
0uzJou4avDvbRH50bXOQUFSgO5nNceoEvddAtJoRNMce8XFvjbpYbak/kgZ8hJjv
18D5q3H0B0S76B63gkLX+quwQsnPxpoNU+jXlanXQnnKaptgYxThHBI7F0GJD8Ti
Fc8pXLWKxE2LuSuJSoL4KyUDS7McjEBsFb8kewZpgrsbtn5hFZRJ0l0E3KFEVIgJ
UFtDtp5mjSQ/gfrjnx1x5M1HXxeWRKkZgpZR7iSMOOdqpeieH9+Ssh+OAgXoQEnm
V6Xb3QzleA7vQejhQaTWiDeTqqSLWpzIeEbuu1CUrHz9tvnLeAmMcUkS4wswNyqU
v3FL4DMhcaaTtCtc/Ro8/12+viB/OCRpcqjgS4kpcy4bRFK4ujQqGg+7I5UTNMjs
E1Wllp1pKT5foHhaV634f3g/dFrLXMT6MNPPNGFl0VQj6YleMUmvVlgXvXZBGWvc
LkGtc3SJGeoctGaeggmkMlZ0ukNNCZnJFq4IAz5Hs3mXv5+1KPC8kXs4cugKPZbL
JVPoQBG/Jk1cqSyEacCQcCqAzxOUw7SV0/M7mzJlKSh1hMBG3VnF9eAJCd3SImzx
edmt7rfHVINk10AMnAl23R2fGKSSH+ysUyv9NHwvSuV+lXGwmAq1OP4BB3Qwd5NN
LEn0iZROCLlsdnZQbB/TyS8Dtfgik0vD3QhU79jqDeZUtp66xCqmBHQq/hcfRA73
l6qIQ7btMOdVMP0KnEB67ycdWhJ507hnmWPJqlLPw69RoqrSq9Q554sztrYNWH2d
DKn8FWFh46dw5Vc5P78G3Bek6rTKNK2CldEXAhOZalJdL+5r60Lhu7XPfRXZgv6H
y5Q4zhuPb+h03v2uyskhBQZaOtPJoUdJ2AgBAZ0NzYjeY36I+K0qCsGdf4FGqMeO
p0CMBAQBITHjo71L9+33pesZ1x4A5Q5IQRSWpIoyCkVbHjVWI4ITj1scW8LpADfw
NH6srm6ETbR79Jt514ma5qfjuIxYHfb18Pafxst8/qU4fdq1FiZ7RI1R/GlyJLJx
LxRFHc+KiOqvah20KraSbd4nnxRF3JDX2AU+G4J0qXBbWFrTBvGIows4TcMsBPZ7
evUKO99zwxa1bN364YiJV1zdigCJIzFbPKTTwoMlptxB3aVM5ii1sXYpC3fQDIiN
YVENs8JBLO9/fd+2K9k7vINYs63cg5+BNwUkQn7dzm/lqX9Km5WaMorAiSXu7zmv
phCyE9jmpTAnQGSj4fCGaeXrrzKaPNiwyhM2s1EVzfGE6YKlQEzfiHUg1QcuMbLv
Ow9jEnQMs8Qeev6Oy5BOoU7CQ7kDew2PQET1oN7LOxmL1ItvWC2m8orWMDe6jnmq
oJDHhuW7WvJ76++JMd2wBa3gwOJD0SWjUtd6nhytqD6+9ChRLmGMOqWcEvPhzS4y
s/eq2VT8XJquR7JP/plw90ghmypTgLVb9nwn0AqadAOC2uPXqUD0zmJ50OD2gllW
LC+LZUodQsp5Syxv2OiltFv9b2KuZ6DXDCQLBYgcuSxg1tLP2OTc0R71Gy8c68XB
n7U+iSKkXdSqtTGIayUe0pwsX7OTvPR9JyITvtUNIkpN+/lRlnL84mfyPJpZnM/Q
uGIQz2QuiOLaLJj/RMD15z4Stx7eOxNRZT4gJEBkLvYi10VobCuSpBZVFIAmagGQ
rp0bhq1SXYJKrBk+bfNHqdJPrRha1vIEP8NB89DtdYyux+tqjuHVPUfjTzOexvcD
B90u6yJ5hEMliiVf4TVbzWx+yf9eGdjN+HV4LFzAqs3yyI43SwtgUPFhY+LZ0r89
uVwfH/NCFIREW1x47Ord72fWIkwSwW5NprHcgsNy5oLYsG+ZR5CmfVl5QfBuz5PW
k5SF5x51fY8Khc7eLpZkX5OXV/Uq67/3uWHv4hw0hH1R5p7QWAQdHrWhKxs6wFn5
JJrKR9HRfPF9FDVLUMQbuX05GYm9ZUs9b6almcwupc3fVjzhUEJJZ+wUZFe8RKD4
FAQU9RJk5VbA6GXBS2WNJ4eYpRGYUwPqZ50jKyxaRpJqlcQG6/dYobklhPuylDui
Aou6XmqDk1NFzdvuSmfqnx2XsAEJQVo/1X7g2R/3YssSKhkvMr16cioGRqGIqH+I
0fUrPzT5xqPeExDoTtB8oDEnKTdShtpefIR78A6+xQDTNWy+mBIjLc66EpqmD2Sw
rz3beXJ282gPYNTO3Xt25NnVVxbbs5jCqIdv+CL9FIaUMrVw1a5wPTs6ZdTEzipj
c+fgt5hMyzQso+PB5LTwkBUKmf1DRu/L0oMfYRipWpcNakH+cHEUG5iB5LPQyc4X
TyVy0nC0wgXJyrirfxesfLIQmLYeQDBI5uAwrn9MKbgmr9LvJmwGYIDNr35bsk9C
HTeFCjtWjy652DP1AWG9JaBlZugEME8j+BaF/sri2/YZ1AfKpRWEXixNhbssmF+H
lIEH/WXfnN/Pf0ka+1pzgHi8JaXkFGrtLWWSjb8McnUgmSABzxdUY/BcIyhJ8BBy
vnwD/NqdhIK6qa6GwcHOiTikFRl8zTkayJKqNirJdJzqGjKM6V0Y6RDOrIR5Nx5d
yBkpK2CTB67OeSz7FO205T9zGDieCrr7cI6Bcf+XPby5N6D0IF8Xz2JICiexRu6b
7UFj5NIowR+ngMNESJThgKS8oPl2SpfkHPQ0YSlDIyZZtx/qWNrMoW5B/MiT2hum
9G/vGBH1EJTYApMqzDpglVagKZK2OPDmAtlBQiY9VwERMPS32cMyy9HxlzkiaA6N
oYVOKP9EKP89dn/tspbLJVLnlUmVUPtMoGkfBKSN5biHvsTvxiD8n2bYQCo2Pf4Y
LjpwSxpmcVu9snVWl43cyDMQdL0YURIWGy4Zjb/pfrkZ0/JsnVJjxIrSS7q2aM1C
oGWuV/U41tCu0zaS+7+KV68KqqSsMvwF+9066vZ10x/bl5cXCRnMspZnEUNX83ks
qkLSMv4fiPoPu+fDunIbqYhn8kCVWlP7mNEYQ07QVf7z9KsJ2VuMp+SPmrq50yXi
Z7tyB9eUw8oTRyOjrpVhg7Ev9rgpWVFpx1mJFr2SCLWywc1oemlVnTUS4YwdDjgl
vAVo5txEbK/du0x+Do8Y38auKTkozZeFf3PNUs7Cpe3EzBTWlxFdXYwx5cOQk0eS
QoijROXL/YwxOFFHn7THE2eXserB4U2sJHI5dzoqVd31bC5b/l1sgjzaQWYt4a5h
ayLoQRcgjaifshZYDJYT3e69eHNuuLG0Nqa5YkH3IbOpbBfg42Aay+BiqiOYvDQe
LaFDu9AQ6zENdli2bpCZH9x+/7CwOsKazPNldioZeZ4pTk+YLbjuFtR/VL+cmM5z
cOsNtKaAdH8Xj1dEms/rWz5P+nGDG4Maar1IuVfGE/QAIm68v5MlI2HdjYEEgknO
m8k1pqCaGBdHRWZ0zgyveWBWCGm8jSgEJ4dfue0cGWnKFxMtazIFBx9cfEtYjQwX
3+Gv83kSHbceTn2ml0RgH0RHiiprgB5kF73ffKDgmwvh1KohEfqoQRcOmokzG+KJ
2eyNsru1+xKT4cCfkdAPqKXarTqq/ORq29V9F08Z5lXkDir30a4wX1lYO0cSpvVN
VTddXT1hlJuc6SqofHxdrPl48c8JTb+CNDrxyq3plvAz8gds37pxhh1vnJzk6AeZ
U5vQZ9a/jHFzSKAE5zUTcJjTWo9wdJoDDo7Zf2kKZhzSeIV6c2pe2axVje+H5nVJ
wsFvPq8HVlJszUpl/y2yMzm6hpIqFiLrtIxaGBH/KmoL7G8q2MFT7W0z4tUrduOs
ha46wKVd40HjwkTSQOBf2GD7GVTax7t4JIPuYCx+0Lvw14+f5WumFvmbmNrHZLC0
nY/ky/lPCQlS1+8rTUoOXtZN6ZI4WDtUDz6fgDvwgRIqcfhDVxYfQJ99wLWPZqXj
aC7/28xJvCRIhNBJQ/ohq0avacXa2/i1WXAGGb42fzmSuOGpDGp5TPmcLTXxSV+N
iDTN3RQzMwuzqmzbo+4ozB84kJN91ZRJeWtbkfnT0Jn0BWwfp8FpLe0djdbbnymy
3Avu2BbxkptC+GKH9u0Vvs23QbY/pfFtOcFg7+o5QCBDT87EuIra9n2KOtADqIa3
L1wxI7h3/wU5+uuPqiNWRI99uNqsMoL3VIiQsj4aSKrV5ItUkQWYuUle2NOV1wwc
GQ9cbEJEKgtu+V/ldXL4sBF7J6RTwCCJW+fbFXXWdtS8rHvfYELZk020l17wp1Z0
diILOCSDAFIyw1TgMpnEclyaAmJ/8mY3BGFtnbMfQ7i5cXuZnz5FRjOYUl4C8efS
h747k91A3CsjHkVWjxf0OFG5RBBxH12bYseFCO6jT4wawjIWDoC35zE763pj0KXZ
hytM3Sf059AxEYU0xaEGlCrVIETBI2hqwC94thagtO9kGD9xoEc0fddTK//Xf13l
e+vzTSUOtnSEquiXYB4CHe0U6RXND2xa6BTjs95qOEcC6oaPG1kElScyjhRdOo/A
El+Kl7htqPXqfgFX1EcBMksuzefyHM6dSGgeUIxz8aTwcM+dXsa9y2u6gUu9+uJf
F4vmIa2YSqNnIkT4hiI630p4HXLp30FFEUoEOI6WfRBHB0JgKlYf69aS9Fsc8/i0
mls+S2MDHPN4beFIClgNtDWEY9vb89fe4PODxyIJyov639nXarxE2MOXJAcbRhAy
EjT5jhhNSLzuwAkloA8c6o/jBgy+7gPTbcZbVwR1qqAbN6iYiNUGja32H4tpzDXA
drpZTjKVKyOHJH2NJ77bj82g/osq8UUbw1au/oOvYfeFyvxc+cO7BMAu81SsGO87
uriU415NvwCesUM/yf6GaXBO4Zjrtq35OKwol9MQVvJfRy25isEm+2cIi65Ld3dg
MF0I12PB3rDi6W7XSdykC/8mvQyT+7s2USrR+fZh2HeMLHUFO7EztDtJ87BpPzbh
XewtFlrdYLkvCriPR57S9Jo4fNPZeumt69gUpAMtgBBjlCowTOod8qQTSqrazwYP
Q/7dbDsV3IXOEY/pE/wKQutzJpAjybmkH4gcX1R7PvunmcLbS6UG3tAzWdBKl0MM
ctt7Edc3V18HU3RTgSIzZ35zK/oac9w32qg7eXs9JCquNPZX7SUMmF/m+jVvmcM6
0vzh+xyP7jfNf1t7eNtI2FP7WlQj5dcR/Erf3HhmDDv6japATfesUD489gD/lmHe
4DfUDWulL0DMZ/PF8TdgDr2HSqfHCh1wvVpbNDUDShwWPeih7r71L8qExzTg9ivN
DWk29jI1jIo5wXD02eFQp77uJicmvY9189xgBv60JJiryWo+jToZVwQUCTDNbH2E
F9ozKV/9k18pFOoEsBd8dSxk8ZZ/dozosE6lFe7AB0kfL+BtXHkQYTdaFk+rCk/z
W+ncLVGMZWbgWdc9DmhXsuJt9VXridyIKu06ElanxPsSAqaPV3Y0hgMReakw7at3
0Gbi+eiCp7HU/EiEYjvEKq1Sb1z0yhs3Hza/LV2mNI2EdFj9c5WUDx722ToE/ozW
i/RabYPC01MUSqVDEMKTkVWP9ra4ZPPp4uVi8sJrSZQCLyAWoN7QnbKzeZ93mo8l
f2+om8AfnUdYry+Ao2ZwWouSPpm9U1Z1DOz0a+5oGibeyxix+7avrqQO8LIR2YS0
a75K3Kwf2ojuRB0i6OACRXL9A1V/RPaR17SODPAf4KfaKJYSLd2kiNsWD8hUHhsU
HwF1ArDVDUjlOKu0W5fN/Ag5lzUleAghc6vJJ04siCUkZl2SAdus7KC+XFmjldvA
QGF056lvEA9zWldOUekvdcDaVDhztS5n59e42qrpn15Ey7K0e0ywmGMHpC2J1cTZ
gCXdE7NZTvKaqhgJrfXRk+cyqoAftVm97VXC56p7CnHFsJb2xQPPcHdvVEj9Rn6A
iGxQwr/yrlcxOoSQiIa/hwFqMEkx9IfNMQjWjKvtv2wt0xpOJgmR2d3do7SR2HjU
Vp2fYED+T2YJgtDgSnilKLRH2noH0IBDrjJ5IrNAPhebD11rdYd4bHO2h72SOCNo
iGaXaqMwxKumV7KHazw7ChQq7TrQkx7Gw0yY0+3rlK8weFdytq0lGtLGaokGR/Dw
sFwO891lX/wz9udMCCtAwINdxvzRe5xCSWPI3GUU0WounqbOw7Ssa/aRDnGWpSub
E3tfbWsM5Ds1laMwwZrlxQzG0QWNsfDIPM7SKOZhmUCgL+zu100R35R6E+chAUk8
019B7oMpIRwL/EP2PaMRGerTe7kQrMu+kVhBj0xIxx4LeZedX+wwhhvErD+dRQ85
CGqX6NkpLa42UoMAbWKKkt0TGAbhMTOFfvmbyZMgIz2gpZmZ4zdwyElAU/xRv8Cp
vCmqm7WUZI75RluTorA1aFEMDvfZTlfg9xVXcfaanFyNlQbZW9HEcrg0SsqjfcZj
fWUVeKo7inSzinvX1jP/4DKBvsQF2hiuAyvBYXdy4OFAFnCy2gwUkbJxxc2p1wxq
VLMIXN4/2VrGqMKKSZH9sAp7yndIfDOfDF4WIgSZxVNM/V6zXkngjrIg1W7PKcyC
AOoS54+3x2aNXvjJAh7c5fKuk/zKCKfS7aSkrdI7e3+HoWgIDDNcgkfyeeWiQuyq
YKtuFU/6jW/7+XoXAFjA7HnK5kz8TsJbDPxSBrg3qjinnVqjhOkmZavH8JIf/Qom
3+e7nFLYsAXs6NZc+g6eY/DriT37HwTylJcE5346ftfWlePhCJptOEYgZvaI1RWK
9px+KGcUhByLnO8H6whHzrUaonevaVR6WAYDfHsTMOn72TfqoNDkrI8BdgUQUOv0
DsGk//bfPgrwauRRa/XcnEevFQpiZ5Eq4/5KMXjP2L0QhjkX+4+UcWGn6NYeQM2J
/AVTYjOyX98ebsZCjpweYdFSPeZrtJNLQoICB34XjRR+IB0hmjmW21eOSKib6728
tFpm4Mz/mQSzkoEixCFg07Tp2+ivG5IonPim6mnTQtWmNvFJ2q3ecO1RBrBmGkX1
IjKKE/u8bNw41cAuUT6Vc4TWnr4g85wXZgIldaQI0glvSCn/WXRe/3LPwr7sOVRt
L3EMC8EREwivBOanYoZTz9kiPXmKlYwDn8cLLWp40b0SVDtbRcZbsEsMRYlBY1wI
56p7Gq3/xv0TkU0R2THP5JVyXzY7N8iH1CQU2fiWoQd7SAXLhicY0NpbiVf/tyh9
5255jwE90eqSvv1GZCVT7MT4x7wD4OS7z/zQ2oKIY+HGFNdOHL5YkqFPfm351Gx3
I/JNAHXK3xwTLzmMFu3eXZJsJISLExwESlQkA7Y8o7pYqCIz9Y+jBfrno4iw5/py
o6Ky4AvGE48VV1MIVotL//ivzKXdH8YXj7T+hayfyYoFTx2fjkKj31gtZWUwH0We
t0FRiyLsC4TNP3H/7W9wQkEmmiasNKr4kuQV5v7xid8u6Jb6Gn6qG2b+KUPS8KlV
9V3Ls+2AA8j5tlTHJPssf/iNVfcrw4McfBIbuwMn8+adEecp8AkXDo7PiFQ/GEZX
MhjgzvZYBhiGRyiyACymu8ZL1aSkOGVytHEDBrcy2kZ/kGyqe7JdzKvkmNIDdV6L
myYfC1KPh+R9QnAFphK5/mmLmcnG86XDdSGqzgDDaV5552J77sYRuq5gjOQ05iLY
LGjOk0PstVs222jzzvZotJpOJ3SiX4TJQxEI7VzPZ/HHMHvh1cC5kcsRv8YTEJzm
DgVvWzJEVsurhkm+1w4LbDV4sH3PP6Z7t1SslxgMke9EVb72SWA4tbPmiHrZTxBd
F9Mr55Aoy2Z44sIbNMogL84I/SBHtaYcsxLxdC+LSMLtRz+eGOwUtVkt/V+v59Mr
v2rteaMKQh5DQMwEoGGlzs73GuprqLKt9elUT8hQOY1SzdHjviiNKlmigD3KwF9B
JdCWfH+1VNGAQPjIbaD44MfirpAFWdT/fDrpe82GbS+zb4YunpL7ybYR236B8RA5
GP2j0BaLe76+ejNOpWJfChqwKL/noKtviEN01qAjomj0hbIxEnH6TpxUWxGZUy6W
bWzNC/Q2Qbx+//2G4eZRIrmIM/bWqWHEAvebzb+cgqotaJsl+1hoTq1dkH2GvYm7
qNZ/pOJhrKmkoIkTHC58/xSQHiggU9ceNjMHoyvJ3Mple6/0w0U0m6+UYgO0xXPg
womchXPKhTV2cZJ6ZJ7rR2yV9BTgHUZoY4M5VrFwamf+G6aHwhKgXm2ckd3EcsOa
9V5bqnNbGVOqf5qCcEsFxEdlwOwPN+4a73vxuw83PkJ8lQ1fN5rG7zcSrcp09fLx
Up0Ry8j+dr07tJYEFRSE0dTUdtJMm5t+zGrlWrl6OvcJzegkdPRN3tBP9SWel/Ac
DHyVyuR59l78+8eGQnv5lNb2pDsP0Yo9d1uHnqXzOa8LzwxJ0kFpRC2XjUjgGH2J
N6tcZwW8a04It2Sk4iBnvJlSn8wMSbXptG4i8dFimnXfHhV0EZI1igi/06Oc+nQo
Ie+fal/xh55rRke/3vZMsClaCI8XNg+JUyhamWQYPBvCZGTBIqOhYEKK3nzTDcXu
ttnhatjXIw0RWNSPFfTb56GLI66ulrP8PMIb4KjCLuH9ejmEP+jM1bskGCPIHCh5
Mz5/2L9egDFKFPuuMx9WbGDGuPSygcgU/s5nKTv/UQXcT7juhh8iZkPJp0+CJBbm
hNRLOBTyIC/wv0/j17FIRe+pSXrH1YlvOUMiX1x0yEP2Kv186scNwzITuJBduOAY
mxwSozUMkodimEIClWZNb5zUxHWASvcwLIzgy2we/oFMRz0/0p9azD2hOWt9Kchu
DuvVYhqLaiQhurX01VurvBULRoicKYGgoP97/ims173YoCVdgZQ8MOI8XVqfYZ2j
ecHEdOvyUSBblUV1UZRVe66A3bmsTPLGD7m3tzqIhqDRY5r5f+5UyHkIJm0LGjU9
B8BRn+z/GZPmc0cKks3FMhd7cMuao9woNHu+WTiGBcLbM8XUjSkH++lwFoTj1c2e
xM7fsTfyL0/f7SpUnozA0BH+VTjH4EtWpXm/V9a6EePy/ObPLJXVaHRd8Xyg8JHX
9B5l9x7/vLDNFptqU5c/Qt6BAq54Fs170OcdZ6SBeLRila5zOIBsUsLIPRJ5DUIX
wJ2n+6el44R+2DmS+LSw9NAwYy2CuGWGR4uO5J6H3xilpuXmxQhAsr4/dMrZhbQR
89aHayA3C09ZeeapZEtvIsrC24hh4FZkVt9SkbejKD2+RR4D+7vreyIwpK4rImhr
jkocAQBKG2EyGvfzINuu7qN3GF1PW6R+GQymBPEy+NyyIa/qbe8U3xmHYJ5sixRQ
NF16/9Ff0JsY3k3Pp2Y9QdjiQOtlWU968dCtNBeLvVd+EPF6hCtLC3N/z4OkKZJR
u/DBNQhOVRl0Qj0z/IKIBZGGFJfo9wk8UNHXBFAXzSTB/ubFmMWfgyuCxpKMZx4R
cn0J/2LOsqn2V8DcQIC5SgQRJu+SeFKZyFaOygcjRhI3jT9LQvD6I8lTwOsTjiBS
Rq0HF1H/TWeXqmdFUMVVYY2HkKWPBjFd2qJImLZGU5rEosn3cNhB6kcWye++9g6B
hsiZ2oM4Q4CWVqXxP8oMWYEkzNpkPC5Qy3xY11DR8gng6jc5omS+W2zJFpAL2CrT
eti+/Hsl/Ft7lu5jfNLiDhFh3Ft3A7PCkrTdumGs6xp8Wl7ujzEcp5A58BezSFw4
G2YqHSbv4Ck6mil8Q5cTDkoXXY+5/fN5zn9TxRTLD+aJeLBgvOL/1oh0sM0A5XOA
VqMWKxahbtqLYE8XoQGZ9kkm2A5vWo7SPdBqAdNSg5TMfDuYjWoaqt1y4zGXQ9aR
sspC17tFG0C1kR7i05FMYos5dcVz2gAe577jgQFCBXoRD0EcCXzdkiDcTmBJLS0y
gFl6qrMNxMaC4le6KGpDVvmWZU6/CMUydEq1eygL2I6MQ6C3SZuXWb5diAIjxy7t
zgVz0hILovbuJ4LzVSb000+rFIaP88TYdD7E8pLNe7U5gG1SJ4tEqmTMh5Zd8J5R
+pwDE9zZ1IrJNcWNH/OFOEoZ8d+I6l23mbDUblSkNxLCAkLbTZtvKGR3wbOiz/y3
iGpLpXzk6r+MlRg6QW139NVwD2wnaIl9cNGvMSx8WsKKCy7/DgboG+a3AbUSGaJj
ij2bpJP17RM3nZVsbD3me4LETIX8oIH48lxj2XY6H6vxLL9eMqFF3B+EDlXK8MxK
ed4K6a/xIgzT52KB9tVDmS4iZ2sKZRHXpo8iEy7104eP+T0BJ3gCosfQaLWadBse
P4dq4c6wH63pW7GKarSChvwCuqmc8YbcGZmIwcCg/DYBNXwwcjxuAXWU0zdstxdT
J9xSai8GryQzGajK5+lZYQepC1fWoH+5/fdrR/ECalLdAuxM9TdT5SdzB0xieZr0
c3gXvDHnIMpAkERnh+cY/921uaVIvXxGgKPZw1zFzTF9oTIYoaYH9A7mcGnoWQHq
anoXWlVhn7At/F7+cA1yhhsX2qcdMpGWfWQA4/NeYf3HaOrofouYXbzr1O9TNZO5
XoXKQXwbdfx1nKEfnokvUwLNYeJvAY2bIsbOr7hIghRaBdhk/7il37LZOb+W2n0U
vF+uQ3/3bwOcnt8CVe6MmhLmG0O9aQGj5w2IL/mcGMU51pPCkxVR7FQkpHBkmvvr
eeh6iqP6WVx1XPWXTtn/QxxPxEsti91RZaN4Ath9x/FnjCXxx4syui49+EqRtl+1
ZvoTV7ZVRxGwh6zrAf8W3lTAOs8YJscKHaM4Mlkj9mRrx8oAD/idlRZnNAIo9rhP
1nloBRVFIQO90D91tRtbc7wA0ErGAX/UcdZFNljwiUaH6A/UySU/huRCR+ptKvrw
Y3/opxFjnir8+jUQQQus7JOhH9tciJmDTGstXwdE0wd7BGFFgtkEnjqAzahMcZJy
f0pa2a0dPzD2QIik7e8dsr8tAJ9D7sDwC4Dhg74dhriT3inw1E58F+17BWEttWxC
XDegfbeQSQs9s1W6tdQpnnOYOj9V+KtgtNJUu8BL4IQBrgZfL6TfXgbeIvJN/2y6
S+QLR2B/8riIYWRUWwNlj5hZP72WJIzfF82fDD3pVVRNTW1MMpkQvfXf3X4XYs0i
uMdn5olqS2d0BCieTC4gy/RC3bN70iDlhXE7Ook+nslEuz+vsu3kfGOyS6dlhbiz
cRavtJCMn6qcd3CDi+IEbfCTW5slRR0+waAhq9Wnf5sSlJeVfAZFnW2aqaDXxYgT
xo64vGprNmHAIAhOt+q7MCaZSk679ZZAYlxcBCpxVTBGKDfQ4UJav7TQABdPHtzy
cRwgcqR3pRihabhrVpBOZcsNzAlfppJ1DXjlfWwIaPqBh8QDTmF6KrKFIz9NUVk7
wh+OB1IfnxAGdSwYrkl4107i8tiTff8fCtjnu6osL6H1t2Ew1ugc2AKj03IWDNFT
K0WTXqa/HU9XIVZXBAF4H2Lz13LGcqTq3X/r2quLSMPdVq+Xei1zMPj2Uull0iG+
L7WgmBRbGT7ZCTX4PxSgQ8/zHlrl2gFYBC1kwm5n9lQVMwdNKiwqLy6sK5UBeD5p
NNFazarFTf0jf1RAOufmGt94UYIK95SqGdbD5mcxlWCL4iEaAaCNA8v5dM7XBZTE
ty6rqFYwiun0DH4EgfnibgLfUPOLY3SDJdGL13oRJL6D8h+YDVY2ls0/6IWGOGH3
Tbdn7rOricTxm4UMNfyEvOr/HgxM7//pCLOGNZOTbhvcMVeVMCAUmAxiWoCx0F74
SdgsvRFmAmkVhDVkzpz8bqlY1/nct4HFKLkvmALzHPcI7x8IDrvK/KES3yOxDKEX
BCUZb9TWCz6Yp4BBfe7RqIFUxMQ3C2vdtAhL8M32U0bCSy9DsWJgRJbafa/s0c+A
NY/kNei3Kh02Sv/TA3wXgbRjJBL30/fks5uOgWjY43gPcGfPdFsS9IHxZkG7X4A7
GZI3NxBTb+LWigHY267ByyhMZF8k89IKq05/weP9PHnIW/putP6UfjMXcd2UXdPX
0PF9Wm1XUgg4cWLTCPhiwjGzzBtxRPex54d1jBbrR78RW5QXcRcE3WBGkX/3dJLa
OlZzt/iHcypm/NNbt7scenmE68n15cIUp7/HHd/12c7a08HIhMvnU9dHuEYPoTLo
DM8EA+tWuRZpefaV60YFcKpoQLEkSkCFmJp4HQW4C+FllabGGC/OtBvAUBOBjuyp
o3wp02qzuYWXUEGNu/bwdKhl01vHfg6IFPwgtMn13E3UTx2GdSDC28bufk81AXtW
ltU5Ebqs3v8IoOQooPJhsZygwSl26xNUTjINyu8ZCIa03hZz7yuP789EPV90Cm3x
ElKxhesLdtwh62lxTZdz0ZsK5OxOIDdo0C8QxxOn3oun1KhWKBoPzlMAH9K6bI6F
Fc6RfSPbLdp+J8aME/NIM/jyicqQnVqFYUlrtyZqC2qu3SNFi44NiE5K0nhWHP3e
a/O3+zA/6s92t4byOqXcFsFtkd3Le02DsDvsA3XbmB+Y+Ijz0UWHgcGJW8BB9j3W
1JqHi0oyZsqzhEpMwOlph474zeK+iFQVondRRIDoZyl7+hV/nQ0qsQ+tKoZQNjzd
2tR91lw6khW1O2uJTU9o5dp9CSYuxRDqXM09KvOVuZ/Gi5qxLXo7kInoJzCmfCPQ
s9TIMAUgViZtF7XvoJSHvv5XtOSE0hkjBGHYOcV2DgrrkjlaZzRsJN64CTzh46nr
duc6dVFnHronq7XNHE+7ik5l7Bd8mYjN3v7IrhTU9FBXVoyPUBE6oYCz823qLuCA
3IoF7WR2N+/bffPFY6wEP0NLKNPnShH5NSURyrmFS8jBaMWf2FdHewVQbEQv8rqr
3OVS1PDCFihyNDWMVODqqYUL9qe1cVT7RHIjOPWN9axgkDOhPxt/1o6V7dahmrMY
5auR9mHg2+SLHr83CFw4NTjYWD2xQK3bhdSsVVaeB/m3M3L4CUd8lWdi5MUDwY2L
qGtUoq33x5cw6NMMhQpDoJDRUAWZ0Hi/BnZO26VRvz7JZXyqW+hwd1AS9hymsr5o
Xck7zvs5vJK1IxZ3fDzlOsQF7dG+Vt9azj54a6AExhs+VWKQr98psmSX2mFSX5hK
0W0ALP3araQ6zdYcMfEZTnU5YnryOx0EyqUqTrFDI4f3oCmikGq/ggP0TMe3dOjM
iMFJHvm0WcouwPAv27PrAfGBu727fez80owg5+IFsyFa83OIW6RtXJ8f1O3YSc6P
t8pdFlzSHBHcqCep58CvPUgO6Yhnu4srnIXkhl0pQLETH4hKxNj5VABakQ6yE2eI
ZV4JykT7cbXXT5afETRKFLM9LnI5I0P1v2FLpQqheIL91lV3JMAmXjl2+FNzIXNu
pfsHUI6IngYNrdMPQMPLSM3/XwlCQVnYMerR3KpRlbaOv2dY/ZYddZst2tQ86rb8
rJsJefnJqTkfu+WrFVnoUvk50TZebYc5ve3oOczM+lL66YAfkPLtH4h5ig8klR7a
laqwOTRQ5aPoDmb3ILYHKFY2L6YmUBEBCmZvCfh/eATOQk8wJ5ErXZLRk96uZ5cB
P958tUE19ppWnnKbctlJsowggQpbCteuaFMyUfkU12LfbgNah9X168ZGGAuVczsd
/3E57xgeKdUNplVqicDPz9yKJosMH9VniY8Ci28lXAee0ZwW0Q360+oDuw+rs11+
7hX9eUfjQKndVXSlFsk51ZSbmUIzhp8sig1LRywFudy01b20knDBGVMy8fy9Ux61
BVXHNCbbFCzfHUvWibUpnZ+Zjjsp83k4C11JOtnUf9G1aOAWOUOfLAfmvy2Wfr9W
DzRD2sheTBOkKG6aTaVIBzWOLYyS4vFrYXFptWfxTGCIU4T32abA8HailzgVsjKy
SUxulpHEyJnmUEd/jdgDJm7+Swxxny1eT7uOoegY6AxfUy/CP6biFZ8SyzZIbIPa
pxGLGAi5fbcusbpmSFnUZj9ZrFmCH0rpf6MQpFmE5p9GrbseQoruXaF5gvnTCyJb
4cFeq9QSwI+UOkmQgCWEpQGC9HBg7I0DJRE0iRl8D+k0pAkq+Y2N7bg0L4HIwodD
N7dMhFG6uCq5F7ki93RIsxcVD47+mnWadTeDpLvW3VLtkGgaVM37Q8TQRZKumstk
VaSsJSHjCkHU2qSP/TVYfqhaHPVag0qrkCrHl7m6vZjD0IdltLMkwMlidW7oALN0
Nd8/0wxE1TvW4KxIkT1V3GxhgdNZYH/TGYm/FH5wm/ZugqjXdxOpDY/+R+y98i4I
igK2HK1qvBM/AiJPyLaZyq+KBtJPuaKWMLZ5+LcCdzLCWczQsFhXA3Hvl9kelYRP
I6uYiV/l5eWW2TNx9tJh/1txllIShjMY5zyO2Cq/dYDueib+Am1fBIESZ71BQ4MM
TybrnxAbv2bt0exno8kspZhiUmWCvP95wDNC7XJSvKNQ7jgPvIhCKGGOj92n15eO
AqR1kTCGuP+GINkT2s8ewmTZnxrRe+qydzqaJGYLI10zpD0mB5W7lEaRoUGQzzl+
sougHk38W76zmsUEir9cPd5pl4cme3i8+PMFoeT3JVvIW3ot4hhhmSnth5SJqXok
nunhJ9XXoSB3raEbxUFzxL9LFrPOqX3SGpziT9jO0AYJC6hwkh2Lw0XcIskNcNEH
hfqXXoex12+4bpmjZ8kx+vAfBLIiIDNtqnglp7UQ7Bu2veM873sHYfHoWthb7mlw
92BNc2IdTdDSrumLIaKUAXqjGdkLQp/V2xRfIVrv/7+IJAf1kBqxrDpkzJPvRRRI
niWNG+/QB/oAh9RPph/meX6PAxHM3ORPcx6BJwVXItAdNpWXv/xTVldIdbjhbrCn
ILBRQ2eWpQNHl1xbg9QWLElcbX0fgcVtuvuwr3tFvl65SS2ZYSxKul8OlnMclrE2
+87rKcHE0PmsYPW8bftWoFqPTKZdR1aQ2RbmTIULCNkJ/PGHSEdOXqxi89a8vPGe
L9llOeMmz/WX37JPz8Ixjx8FUw/IEhe4sNwUV+gIokAEs1zdP/z5pxegxwWVEUkA
54yYExqM3EdW90Nt86/mfO+MCp5d08hAsIP6JcuKJ9juytesLexCG/zw7cqNgw/l
GwZlDn2TXSM66267cOGxgaFlUyy4jq9scNolVfUkwaDRIns1P7uw0a6/aoDWrbcE
v3L9zMKSDNjIRihqq09gafMTt9jo+TuHQxEOYjrjhPUAHPOIOTaP7lImZiaBFkeq
QJG5xnUgUstJhLoOi4+L7HtshkOCaekMLx0DefPQV/MStDLu77gqjcQeNQVjHihG
KCm/LUyLap/m/7TzQTOfRiYwEJOJmi7MEhNJ+MFsF+C2UE8CFIrQgb4+wX6VJY1t
S5dPlnbrA8HiMli3AninQFCnfXb3zPxCVSB+bmM4COvP5o7JlpFVl6Gc3uqRFPtY
NTWiapUTpsh5NIJvLzxKSg4FbJGor9iHZ41f8SDNyj1WGQiuhzPzOmE0uoTSb50W
I8yNJt3BxFqV+fqJN3VAkR8ZoIeQZQ0P/pDumVc6xZjLLBsjoht8PgDPXt6kgOX6
A3Ou5rHFIRG4xiMYHnMaexc3xH5JseVYPRgYSv8v+K7buAqKUyGyqooDzlWbibBF
Mraec+TrG2UCGCWu8BKj/ABtBoNlL3JxMGnib5YzL/jEi1hQW2ahKEgv1tTWljjX
OjADBho0qCI4X9BLCHFLmRDyAXn5s7ugGuBMwBC2hpWpVJpPupAHwZtwUe/dMezV
VXkfTfMUCybYqLzVTz/NNXP7N8ie57lQhSd4bjfn2lPoHbd4jCAsWYTy7RpcScI+
h4htCb1YMFy9niFYBJwegjH9EGi8y7Oi9aMEskOSJyDXaFxCZmaaCEfUZGqoRQfx
R55S8RL9W6EOtfcB3JGcU7u1emcnGiCLVLSeqnvvhU2xKEcppI/ct8Xd1bo0Lm/k
X2B+SFmoPrgH7yo2AHsH8X96XaB0nOrDzCGPAQj6xkqqXVFZTJmun3OE0gAlraiT
ShOusrVa/22+6bV7D9qruULM9v9oXO6uDjNpLHgR6RD+BwOdxiyVTObfnkd4cnIh
TmDqHzzZKlVm1VYPljk0WkIHIo8pA61aMDH6J6cw3P1OHDhPcONiPE0fUMHzR+G1
nJtUDha2/oQFYDz4Zr8660wPvAAu/Hw/z6ZtgVE12NNQrSHFu1twrrGTiAy54G/i
KlJkSp+W1r082cX68ojuF1rd9KIs60n+tSVloR4MuU85D7rQaV7Ea8IDaQ5lFCzm
x2rwxx2ATNmatQ0zvrDvP9reHsb8LS98jt8bN/BX5epVW/sb3w1tbTQZ9byruUqB
fsLvBT/b8l7DU+ygmkd2jcexDr8nfQshrC8ZeHudlMusXSMoh2qp3aJoff8ZbneI
ZyWkVqGt0KJqvi6aZ6rIaV5qy7pnLg+idQefUNsVJoSIzNXyiCboZUBJ/gECmlBX
ftSIOzg7rQcD4j21aR9k4aGr2I1GR9MyYMtgXcKdCNf4FcqJsx3Und3oQpLyPwDL
L4fZa95HigGxpLFZoJf6QBgCYzAuEOBopVx1bnKszrd/rFL71sOcPS4ZmJaYfmfL
LfXVV+p8VAz3FZzVynxBiYscHMbLjZmE2N6pKIKV8zyKaNj4jqdKdlp8sGKVwn1e
MyhZbdWueh8cPY3JzvxFvAw+CjLuOJv8BM+Tr0OGfxtR9rhl+6XbBcHFM2LvpE90
n1ZL5WO9iWK2Ijp6wUAztFPnauWtTFMiXTlrIYXENTsm5IIeYBJCJl2UAoyLJKCE
TiDT2JG9rmD9s1PNMj7eMtoIKLTBpoais0rId+3m912EJI2hnHsb+xmdNrq4Mz+E
o/POgEFA0MmTxgUmk2u4Rt/7lJbiJ/+F1fHKwevFvuMmRgyjwShcWYOjhP8/hhnm
PR75UrlhasfIdS8JD4ROPEJuiWcmIVYUIeLwrrqRTSxPAVwx9JMgp+Cy6p10qef+
zM+SKkTxJSzibpq+fMP3zy7XWYnKed43LN6ZU0dSJ2wp1a/I9buLx0nxA9omCEGZ
nJijOocIMOOvlYU24hFS5PjouWhZm7brCNBvuzpMCp/bnfi79r5q0/AJkIANhTRv
B7y2wSHifpNCuPoIVR0J4fgle7NLobmMar6zokdegKVnaIqOqGXvMLkb7et+j5eQ
FzW11dGCxF3HPgVlf0pVCoh3pVHYxr1Yd4esUBoQlnV2Pir3Yl+jbYD0dRDr5d+7
Pbjabk9tGVfWZR5QCqDweL7EvI80DHEXwtvZSWWo0UkyRiL1Y+U3pYIR60NJfLy3
flnpQDduSpmDzfyAkfjKsM0p3/ZfQ567G3EsE9VTPRFi5pm+oBPAWXX0aOLm0qJa
rKATHJl0COYlf7Nd6+CNXRK24veNSZ2eZ9Mm89cb9aPasDIVRMSXyIb3th4AqM54
S3x9cCYtOKnllU0FGxpbpVraZj/XdpLl7y4cMuLDuP+dMmFomvbpBbShpmMgOmxg
GYKL44zKPU3l4tQ7wt0TEqvn5KHAYrPAhBnRQtuFWinWWPiLUXd4HQu2soJp4cE8
DeOi7Ga+u6o2FMnEX7uXyeb7dqqML+SNE9Hudgn+ZD54LF96BIjKj6swe53DES5v
NAMBptXaPhnveAqxBup80ICsYOw9KSHPgVYAtdPJtkRLj4rf0VgpPhoOyJP3I1IP
dMRBBn87MRx8nvCTA7dxPBJ9XmFEwhBie3lSRQeYtc7MAcBfd2OZD93Z3E5lQCt9
Vd5TjNW8eweo5vfX2optWoU8topEZzVA175uTPCFYBZDTAliv9GMD+4ie77fVoIX
zR+7nco5Bcu4GOlw5/Jc81FgmUCdy1gFsruEL56tjmZjkLrDi7Gzfa1SXu94KBDm
OorzUpwN860VZuBR7R58aZtYA0UdklZRsqXpsMKBWFH34xI4ZHpaobnxzC6Sw6J3
n21F1ytVbMv7VRtE1dMwFPTKCqhfzBmp4KCUkbkNw69N03uVqzfldmJreyIWnz0k
xg9J5397DWYLShFAgWPgEkmqwo0C51lU6rh6QYFEBM0uSxLnfzryddQGOxpcXmXy
AI/YVrJPpYpfl254hm9YqO4Zd5n6qWudRHcJxoTXmuiD9mpsS7XaCOY6mC69SumF
1iKj/3jKPXM0SPUXUw0I5WlzUlp/nrWdo/QIckgqrPeyajul2bQJiQrexKCqiMu9
YNI7qsOwlIkvARkpJX31BGSZq3tTyKJXmmm+z/YCI3+3Q+df9MYFVKnLdasUug0v
AglrRmYhH2s5XVwWeYajrclXfTwLtbRcABpA0qVHEz1xtOUoUADwpyoKW86Y3ii2
hCGK+Kn550KrHOt0KVL99sosPLlVpTwqrSFifs9NIkkME5+a/K/BxHCZ1icgK4RQ
2nwzR7+AQkMSaHMYAG/QmiHWFZ9LVhElryhIV0sRG7TjMRlJ4WZDFjg+zBrJ74Wx
wpR8hBj3lw1+RBh99ZSHzvgKvvV8VG5cEGEWgLPL06rzNAkygmzU+WG+KaLGhDVI
JFTbIbMyu0Ptkw5sjr9M8TSDvmN0c1eogG2B0MlBHVsPP4rzichAf7dQZOPGgB8c
oSU/GVsbA00/UpgnOMxpwkdAi9wveBbgO37lLgrWHWSMlaBqcctpCpP0YldLgg/c
X7pB5HZuFBO4MEaJlUqVTh9Ieq74PbnZDS5z1LKn4Rp6bc/GBfMeiwvytYBVRIF5
zSFsx0ZpDJ0oMLi649EBXY/d0ASufW+pZiuq2xZTnjZjwz9OaB8BGn4opbdGQQY6
p/L6R82s8F7otbonkvdyG6WUDb7iCRAyCeiT9zmgrtzFbUMOw35CU8x5m149N2e7
YAZFP6UTcnidXJ4RxJDTCO0VXi47H4AwxUN8xictdwB3nkQzMxaU7MVb6nbgLXgB
NZ4odMt1xskYY0ka0OVzrE0W6IZAgwliZDrN5gvpGTYtJBPehl/MfHAA25YkE8RD
RtPXilMk9yuCk4PsgCQSNHGUtXpKVWq+pnMxY8VUXFrljKKWyB7xsLcri6fFU6yO
eBZF73/bTw01GwSNcn4YWQeIByIWK2nNH++CL9MaMGow3C3c+4IiUl+LvuIYV58k
otFs7/qtMdBu4Hg26CoHTYQnjg4wCFc9Wv2EJx+mkPU00+CdULI/q2z6DAWqzlKp
fmv5YbLmLdNCIaPgYWA/B5J33+tV/q6ISH5k5QWlD8vVFEhnBCafb3f9uph4WiTs
t5XLj0rcKtrYqmcfX7A0T87cAMXJYbsJH1eNJjeuzV5VtZI79rGAMWyjOU0KUhCE
M8flachzMDjIc0sBFtP0x/J2V1DA9P1PydtlvFSTEDlQ9o3ueRJtgfVisWYvcH2z
0BxnDwLDlH109nb9NBXhcxOyG30YjsxyxszXoclJlVHSnbXG7AeRtE2jIxo/BUB5
vSSeT9eyl6Yo0YtV4ChZtxff9gru7NaZpckbBQegkxTJ73YqwrnIKRWMixUgsvnO
h5C3oR2/1VM3zPv5zczJKI6GUN3m5WyRnTAmdhch2cIkx6hp8r6MOW4nnkDb9bfk
RUFri39J37l6AgY2/K3QNfuBlo0kKRPFsPOPj8kB9EGpUyR5DDQWD2+97CVbu0sm
l5LNWsu4VOPbSxwdfTEUi0+4whMTC7KJzdNmQ5ViVNS5hI3JlcubwddU35BN5JJT
H89NIkI45X7xJBOU9iwVkdTYiMLMrDam+Cy/6Aogj37tj27wbEQTK45pdu1CrlpR
Y6hYlvWtbNvDyhdkxCbnjY7bE8QQJm0EdHaiaWAQnKdKDSRSjc6glFxC+nmDprEp
D8W7EC26KBXnlZmzB2sfI2vYt6Gpcu6Ar+eEQpQ0g+qmG0c++w8mQsnsF7vAxRcV
GLLudaAiz65lzTvYeN1jTKlLvNHt9C4g82s8A5uX6/u/bqfcsxLcsyeinfuy4CLK
J5Beg2q3Zs0hg+jXpIWhS/tEhqo3wuaZlobaLFjS0nFaoygrySTtkrdENklqUaxE
3nY4EP7L+fRxf6fB4DGWNgNpyZaqUWBRxyEE6gC13FpBHKU+DjM7Po/oGLCNsksP
nIj2vw/WA+25qR9qLfkYfj2wJxvhJwFK1stbtLGYxX7MuKJsl43vIZVgRVqsqmls
vjMGVZEyWIXgwe7s7TPGkkTIOZueDgRuWCKN78jPJG3tRc65ss83/Jf+pogqoJ9C
LQdaH25OMVi4pKI2+YjyHgjVigfrofozcaIwpm9NiYdzjufeWDnG8uOt4OK5HI43
lUEZnec3t/TLuRMrjvd/9gDDSXzbmlcSoTOE+sRBDdHOHRi4N22pdZJ295reBSCs
Esimzz2oNwAW35jcnYdr6TRqHtQLr4Yw/Zf+lxctJclIcmcLemZbI7AWJ07ce7/Y
CBk+Oe+fHv+/pGkQlG3jHhRIt6G8FbInnFVW4i3JUODlVg5SrE5wyes1AZoneZLf
A6eUVbQXq88YKsvE72iOalm5SppKak6j54kstMYskCs8UZJNLezsBA+uuny5uBta
lNZtB1qFiOJ9DCmWV8gogytMHBpzZGSs6k7vjt2pdByv/vxVx4/JYCKw0A6daHtV
ZMa1I2NZQM6zbRlzFWvg2CvibfArzQLVJZli9fgpGFyKXbM1ZD/ud/lzHlzP6IQ6
et8T9MmUtGFhlNXT+salSuwUfv4sDLrVBqa+6SXvYU7kQb46zfaQBbJPHrCo+/IE
H7BcT4cOjZAv83XNgKUS0z5tEjXUtoNcBBoiKZ0lT3RoLXFvCOrTq0Pz/1JQ4x95
XjM0pHC/U2z4vCAi9T6WBKVV177yNLdRX+Be/d3WiWglQyL35MremU6k8iL2pkJ6
V8MHIbrvtJdv8uFUU2z6ZBK6opUaAjjhudlezqfKVLrogntdOHBYlUBwLAyV9m68
ICKkn+v1maLvo9OnlbHRCJEFhmeLr0MyxNXsxCgqFRzs8l4yJ/uvAZ8z6vjmbEls
ajyFztavJ8ENdkJzIvlkw3nX18/9AC2I94zzaLSkBKC2Au/6ZaBMcbXAf6zhrU3W
4uVHh8gmA5g3PCLoDOKtYHJtVc1hRlnyOaUQSVGh05w8rdfuhyQc1VXeXcKi81AA
xm36VP/xh34HR+oGLBXTQlrsV6dzU3/fmT4rBXGqdKNQ05xU5fkfNTwkG/g75cs8
Ws2Y0bnUkLsokAOZ9GnMwuQx/OBNqq093dgnsqu6dqEZQ+rgVFvCRT6lafY12oVa
RpUZYSgCw08+VrLys2rB0LfR0XPfXdP94qFxoF4NOR0yoKjs/0ss7O3KD34mzyc4
gN+fjbgxqIPx1Ja92nbamAWQ2DJeJXNqnPBz2kW6OZWzMy7yn8c+kfiVgLKbMeOc
947fJoEXnf0xUASEOHLwq9TKuLjUq6jYCQ1uznrX1Jfadvpb+MZC3csgpVQ8mwOy
lkXtakmPIQXaNEg0ayTDp8WNJ8sLXYFQ7dF0laC6NYFhAmwyp9l/PjhU4kBY7Mch
qSX+FGItZDoICGixHr+dAFLC388sCZp7RMs39kXfOrP4TksD8CR45w9G3dvN+RMU
Vidrwm2//XIw6YiGceRY+3JXYq7i8SK9Q/ZYNtAVbTlUKje3qpmYOpuMfgDFsxox
RutXo5wS3Q6fpRfHLnTs2CGoYTfVLYQVjtb5q9S4dDDsR1PPdDQFHoim0XvicyuM
M4gx35a9LXYTardNoNYxR5KLbAefVlRgneXEygrrfWK3jKnt4f9VniezA37NXzjc
nouVRyrUcy1mkgYN05iSzE9aZaZterJ+GzEpD+JlkX2cv6UhEfgm4e40B1mxihYx
keVtf3akTilqYERUopEz119U2dr0y4722RCqsIfe+EDewGWEAwQlrETspC/Dxy/j
MNi3Hk0C7MuMGFfp67DSE0zZ5uZQ1qSnZccyyet1RW/L7snJsrAxps8H8SQEDq0F
PPhieWm+oAsVR331C/hSHz6Z6Wp+fvPMA5BGVcshGoXWvky30wx6NlQokGhET7W3
Qy+ytH0WAHqTZVAPfW4MG28zgFqheTGaoPh9hmSAacoM3NcgOetycxwz86lSSOsu
1OqRKabQ21PjMonPNbShKuKY+jFy9rsNwMDFphEOADD/PFFdJ7bR6mMmPAA6mxgS
xAH5vX1ZdmHHu80Zsk6MZoyFX48hj2un7NjUAWLVdrojX8i9ihDvmqbzpvplB7AH
uAZHcXzWhnLVatUv2FlUXlIe3l3pSenMB3X5enOCoBaB40cyPRUo6WzPBSrI+N6F
2K894BlOkSkqk1oPoBZZ7GFQORCtj/MUn85OeIJf62rWmvgwePgO5vRh+GSKqv44
AuJAHo49j7QSLGgBgmbauofhGHD17sdozt6B7sKOpG0PrE2pIy+FmqZt9CEO/Y36
XHwSBM8wqOqOO7GYbmPB5syFfB+fEdqTcd4GFKPm7UUZVT3JMOAtTn+ujv/8RG12
n+kt2PMKqTHh24rAIueB/9oeo88huTTw426UiQeZJfTD5/miDFdakGkm+erXuM9o
f4vme1hPM5mxwpS/S8dtY3qx7JHkQI31PojhASv2O/HgXu3O9t58SSN+5+OS0fuZ
3vQHFm+vgLfcMxMajFx/HO84ulR60XTArRjJ4LULCaNAgaivSyF7JYTEr5DPjdhG
pWerreg5PPsXWt/pOj5YrtSsp7U7oCit+mvOjsz/qJhOutSss8/Kd+Nnf/9o/dfa
oimVv0bM6VDMcKHhaGiop/5Z8GfMOvd9IKttXVMcognzpdAO/DpjKzyGdbfVmr7a
28lKdScMSzpA7OQOwIDS1N4QXUo8cm5BPaOz+rJCgYzES1X1d/BVZgezyn/8NtdO
XnGJg+8LcqPgSUXcM5T9xAW1AxcT3ntpg/JVAXCuZcKeJzcYnEPINEPp1NNT4Dvx
5Ay9I7EGu13RRif+LUlA0vv/X+F+BU/vbNAlx6myOHbsDmx5naYq81H8P74+ehBT
tc4OYzIfO+zihWXO+ANCxfsGvaJz9V8IT5tf8CmkRkZ746U8Obs+LXBml/K48v8s
Q7B4v0h74v+NvF+cmX0HVe0GKGcVkmRUAVztliGz2e4AaUfZlYpfzm+eyX4ImWsx
dmXN5O9FEX1hNczXI4mobmS+Fy4CfPwhX2eKiw0bJOLFQBkQK1Z3QWzTrPrfCZgx
ahFQuYOM7VZzSOMPyb1XvOkcZJO9nHqKWvypcnPOco1WveWmHHbi6bn263dtLmuR
XAEIWFa0w015jKQB2bco2q12mWPXDGUXWcovVLePKxKR9hmY+B1L0GI8ucfZ1Mr3
M42xGIqRQGdWkTdqwujv7ki0i+Ky4WdST7IJX41qW7ySN5m7OW8WGWDvEQenkwPu
OAk0VSqzhzZ69Jc21M8L6DWarzfv+wilhzhaQrYpADWZe3C5QzxPl0Xfv5U/0i8J
OckmoChAq7vbff19zWS2N/IiD5qh76lyo1I59xvxJy2zQmUCGswz5FBHRCX6//8W
G229q5RvILN1JHiB4V9279VXzjFBMbZOr4yCDS8EjfxpZxDBRoI0SLKG6dpEEdgu
/CNOeP7/tOIPM6/cKA7rTgz1RmyF50NwIe3U6OkIApnPrLrEjiLSQuLgQFshPA2H
Y4tho5toaccxrkBLFJH/fNxWAAUcaZ1eI79jiARSYORjJPHqN+WsQ+6jAn7gFdmR
TVZBvAw2Md+LCybkmKHmKqUVrFohMnydSodkmXSX8i8q8IF+NoerNbnXhY5aSHzU
s4iRFr0YinYzd15TYtyjZTu61d7GusBbgweuKU5hU5PSt3wsNjECdEeIYGG8Uso7
ylhcyok1dcBNzE+lzLVTi+9Pobl6lt9u3tB+qaxaR32ANCv3SRWgmxUHWnHMuXPJ
HPvlSJ7L5AaY+QVeWaoFCTrk3OOJQ1EtM3yqfyoQ/remY9XpV7FiCzvUjkICd/2u
xur/TAN/6ccNblRL1Jy0jxvdPDKIecuF5IOVsYuWy5ccm59O/kIKXwWfbJa6Muvj
8d9X7DjR/S6T1WfCYMfcUF5Jycw6v1UdLMKOQfdtE96IRS0yfWkjXRfQo+Y/UbbM
HjMohw9P9ufIpLYFCzDcOyD8r3B0ngC6EkczTzuBbWZZTPy2ZQHtDoiO/K0Ha9Uy
MTeHsmtko638MM1499qWT9A6aU8ItbOSozj7LyDM2G6uj2s+kdl1lMHMkzKsFKx+
SiIrepIdxTIS57xbwTfMgF3wq+7lhH7dMusi0353w7SkvoGLxAQokHVad3xQIRln
4Yi1q7SRdp8xig0lyjQG/ewCDQRWlHRPVgdSoTnPSd04Dqv7WvHp/iYNIvo8oz/l
qAKMcjbd0137mJMuLTJf7fqUiDhlbbeFzZc6kVgKZeIgJNeq6eBHdFzElcR3EA9v
PbI42UUOxdakWstquyWVpBhS/QVYtxTII2f962uw2qMclfaWJKDL4Sd4pfZoXg6S
Gjo9WpIjv8Y1Fw/tvgHlAp28mZKEXhi4+bjxossEKA3314Oo982JlMEp4hg303Gq
rMAaU99w4vnw/ovtvp16I1dpAIlyXf7Iy3mwmvNXg4tBSFoTIAWf3/Le45FLCppy
I/8fyM6jMHejb4oYR9632bmx5u2ev9pxcmuCfywiZIkRmTE8a1z9ULL6YOFD9oTj
t9nkqnynzF9Nr04808vzs8wCYT3F/d4v678z2H+b/OE/tnZ4uNTW3Lmnh64fMp41
zR0ZTkKUMsqb61l8mxF2aSTBq+RsVGxKe0BnfqVIauD2wNwfo1Q16TYkJ8tfsDfM
HAJ9rEzwIqB+SJslCyqfrzMnHc52Q6DAIGPJ8p8UETIhpDq3oMerF3+qLRCK9Cpl
Y3Tht0pVqcmuRdJmPR8MqdPrBRA1M1YhEhuNyjQvLmiiJK6Fj9XcgDJ7WOy+G0+E
erYRdB1c6hnhYHA896wHBx0skG27ZOSiyq7QFcdAXggfEF7CS3s3bDNR37AT82OZ
yuB0LjAvnrcRbLUosscBET9kYleHz2SkgAAoL6sPfug4UdOcVQVmUtOKVVM8UDOj
s8nk7R/iyo85pGu19riWcaLYBTqlmP1bjOkNxp/kdoS3H2oRhG/BJihHyagm4Glz
9Y75yO36zzJQvJHuU2TcFd8TW0mq+rMp8WmG1+tcDg0qy9GAQSfn/o8Km89laCpv
eN7cvdHK6QRqI03GvYwhrSLfPUej8Qpkb2jG6SMBTuA0FRwRxEv0KYiPtfYvZOZE
FmDCa3UDArUABsolAzxAERVKieG+zuPc7CGFpotoYmOVm6dGAqvYoNOw9RK6HTcO
8bizDDtHHcejRP58UvrHYwGNYS/9RhkOEx2cK+HhRJB8GJyKFaeSalNUdVCc1wzz
DRxmuAyHoxnJa1kFxdlgP3tFBfcBkly7y9/sD8g04In0EO5Fwv2g+YrTgVCIIubl
bwOEMxnQT6q+2K7SuDokMo3xxL0qdmpoGklrZwbvzR3pSkQVe/RFrSjCjL/uW8OD
OLN/jrvc8xV8xOW0NrS99rUoZiNv3YvmT1yTCSgr63MRABgFG5z1QFP6Ky269sVf
Oddd3cFvfFNq7KeStNX4mHEpsx5kpy1LpRYKuGNzVyhwcYUxZ1JWDiJp+1EcTG0v
cIB0hO270eAZJRY2gnFe4SApppEvymUvM8x2E8T3o4UkDIOdPoq9DdLKvQyaJUTT
/5wbowQpTOErRjjCbASoz/2sbIrNihm76J5aabKAqStpH5KfPMbbaeWETCQVGQ7h
/lZIbsd9G7pcrxkwOXE/8WXQ/UaHVXmsYVySm4DnJGiRuVjB+F+aQv3X2PqwsrDz
rRzocaH4zz15DGXDTEcqNYrDZQ9iqqrQpuIXAZs1GjGDblMd2j2i8X4n8Vo5ly9I
wA0UJaKYHcyZsDl/uADpxNcWj9xqyEur+ae77bt6U/WxzdobD0L7z8M5pjQe2RcB
9aj5AUT6cwsBdCEzruS6vVhbpC9J95pVvNTM+7RqwZSRJN+5Rov3bvpH46+ZoXag
H4ru5vgsHOj7BH4rv+rM3ZYia+uqq9cPUmXAUxMA5s5gP3Hmfn1aYhqDNvA5piF0
m4TS2greCIHUuwzkP98a0/Ty8Uln8sqWdPj+8ecdo9UIuyR76xwudN/q3DRnFiF3
EdFO0FIRPI/pktmKElGp43gPb/5ejuIqxUZ9JhLQv6eHB18IbbTXKM4R+GbxWpKw
VOk1Q2r0u0rj/aHna1m803vET1WJjPXhJWV2wkAhHXWE56wblJnlRzJzByW5zfTd
pwNhZmkbQwvyrE51f58jv43J03zrIAwDPb53LGz6G0VOXS0bDfm5uJG5X1zujArp
ygd3HrV8NrkYYwEKNSvoA9BVJGOeFMob/Y2YG3CYL68YO2bTQlfHc0ajz7exyumG
c6d3G1SQqe9UOk3K1I866N+enYCJiNSXKkWYCNczxo6obqqGnMyghW5nOwrY/yeJ
HPaAnRIdf3k7b3DiXE20ECiRmvZb0HWuCtjls/EpJKNwtKzxn8CCh/eTAXzSMr7Z
JuI+PaS90JzrIewBHYaj0LvU9WZNDJlZY8S3eRVYRiVMGgRpwtvmk7kfj8108qdn
j3ghs8c9BohToFa2/bee+1MWFvNNavTnF+7aZO/0tOiyyw27UrwD7y1opAdH5ta6
2mHjpUIKqMQUbXNadOpH2yx+oFhTeecggHoL7ckzQBDDsJ14kvnudEhvc2gVCOUQ
VU9GJamicOJWV+VeMScDuPq9MN5A5AwrpSgpGmYeVj7sJd/ql15LfvHhNMXaF7aA
5CA30eR7kQ0iahhe3JU6WDb7HssAF42PsfsGif/cM8tdqsQjDS/77eSWMs/Hgtxr
Zeo3OW1Ira62bDAJsY9E0k5RcXrJWr8bm7TSgkI1aNFglH5cxuUvM+w5Z9uMLFfp
eyW6qdmUFPQYoJ4Wt/FLRCV+E4HruDZFdEbyF04cS6ksy9q8BWGVrlnXW3TZBhV+
JBswQB61nqf/srPmcgOCpHQvY0QSSGwosgNewDo0pcYf4HWG1H9V1lxmeD0KSPX4
ogBvEs4INkzajooeOdZTb6bLDNY29JpPgSWj8M44fwh/i/tgJIPmN0LLs7icKTay
3giHjCjZG5TVQVsD3fZQqPHW77OCYkFkqvMkBS9EWfMIT82MWfgsXga3NSrexI7E
VtzcjhVSFSrOkO2lO8YntWx+CUB7FDQZaXY3i6pwROWkiFKlRb+ocSzb9TGN22qe
oWeLX5Zc0gUnyt0qjdbHk2gOeT0LDwWTt/+nDkSs3mkxPvIP6M01Wf79ZugLTbxb
bf5HKj4JuVPcG9lgl+wGuWbW0q33ByZujUPv+ruV2kKsBK4xtjqRVJ5nyiVSxmF+
T6UGWVGpntXELJeMHxVom30lnK0Ko2VfoL/cU6SKOEqt5PleyDFhzVcuGHADnsfU
lUYUTiQDP3gmQ7FF+TsV1GOlRtlrBtOqECatoQHsZuSReU01w9YZ3c60iJJCqMiD
RSZTLq9p2wslQeGLP3SGlJumCKGWn2ytCvcpQShEH12or5Xt+BWRKsTquUMCswHc
qTeHfxBnNNCsNiuMtOwLhlFJAaSRbSiOxP8pidw6lc8SGvf1cRbak/xEc2bEfHY1
a8/Z9Xe/wQsgJviWZRG+B5cfPt9OMA2/GCh5kTqdkPM+KcRjbfLhxTMQ9H+BxWVc
MR5XWQJCVUaTDIjR8WzPKpUCJC57FTuJFiZW4W2h9dAEI2R40J7Ob0EnmxH+QbV1
DSY+jXRC/ro6+ws54jZoekXy+7Ncf1dKxLJmMqMaElfadDVBk4o4SUk2dfmuwWyj
kaSNsvDyPZafoyagmB9PQaOb38Z/6HuAfjsXCaMAE3fSUY4IeCXktMk6sdAWRNVD
WKX7mKskHVQFcicYa0UX25sA9vv/7g8WoZdB0XFMAF+fgF3RfnufS9pFhPpI5k44
AJSu8ZGs33QuUiwUTkuE3qil1DHqk9+28HmVmCFpRurr13LxaNSUi8uY8+hqVIIp
bZMcVSivET3h6TFALqMt9mJXFmDeqoKZMbwMzGxQIQ6UNWpI7fCdDfE4Rre/hA/E
hPNHhIhijDQe2gJzIduKaLiY7Ek+p/Os7jyHx3xVHeDERzcyjn+HiZY53/H3EB2U
QWCLWPUHk4eiBqQL5PTpMEGszMv9sPKnST1+iaTiDx+uLiG9zQreKNweQnbiPqPF
ekQQPbi0Rgk5Z2HCtIbpBE8mb/9lU/fB1Hw1iAojJvATNSd0ckky48927GdZwZf9
vSdl63XH8Bxl12EHgsCRQQGqrK0hZ540jXoumphlJ5njBLAgEuNpdpqdabbWjQkc
NivznBnKwIpzkn/+131aTPYrApAfhDcrpHSknPawMMkTpYl/oaTIAXWpN3CSVY0P
3Uu35GJnKSV40hla9IHHe78go71U/ZQliSMzbZgTeueR4fuTOPyEawauCD9a9kvo
sALVjPfT21MTBcbecdb9s4au5RLhtzh58+24TGmJEYwCVhcC/gWPKYNUw4d23NI3
dHmC/HCN8r/bNJFA3xZcPMTYLkNaOjR06Z7Pu3ZY6JeI1Imj7lBBne+VhDMFC8c9
P0t9BsIgze9QY9jCVYPvX0HlbWyWQYQKE5NVKQDOTXFgiU0liLSlItkhkzmpK2Rm
90cnay1M0RmqDHCu7xMvffPG+AoVDxJfOZrDSq3HJ2iciAZHBKedlcZ/9wRXAsoB
0gDTH0CIxKrVEmBFBZHbXI15QWPwqMxJVozSzI1YB6zMJ3OVDJDUK2ido3LMMred
Hv7HLEzh5QUT0SjrKNvFoXYb422Kb05ytKerAzX+PM8+5bIAdNexUTsao++PsT/y
8ejkMdKr64fY2GWb44uh7KvFlHCjHYNhxAUx7009fhtEDDAnBA8oLA/qdfFZGLuV
sRc78bn6R1wEkcZfFugkJ5ZI5aTtQROcmGkyTYvDNJvCz2sSo0C80f4z9mxIthF9
59H36WvwSioy404YgMjtUaSH01K3bQwfUXYuuj/rci8LnkCVNug8qErR/g4HGazS
ryEAfKcQ1DlJG7n++Y59K5e6enLigOA/0UQGu3mHSOQ/DVRKIBjM6MujDfRWmz0d
Vs+a8qDR5rglojO/58uqOOoI4UUT2Vf2ZUbJDxP1PLPZWPEJ1gWaCh/Ihp6PjLm9
rFx+1IfSx6Rlt66OmBAMU7WxJhTTmvGqdUnxI2gW2jnR9rdTu9Apsv4rHj3WahAJ
0iWO9k037kPLcEtB7RUDfvQAam1Z94riyf1CW64s5fm+3hDK96eMjoAGyg4vNOuo
4MgQbSm6+c/uy8NRp2tBQkGpS9ea9KKVrQxzHBa6R4eFpHlkVtfdHIPVqSXT1ShC
AeBGqWswsvr++XXS/htcm3CUU47DjjRZF6Z8loSZ0GM3WhJOfUMM84ozOG4imGua
vE1BJlBfszqXucKKhjKAvRfaMVHQ/H2iiGjYr2M5CczrBr8mtMUVYtUJO+ajH3TT
zhIPPeNKlkODXu52Pp7fE1kBU9Q7Zm7O7bW9g66B+JrWLrqSfYwE1+fGkm+5ytus
TTr4M5BAu4nqJvdNmW3PhylKe95fnGARdIMZz97FQ00L31kbOHDoHEHSAYEgtbWk
zC+//jK2KDG/u00FPiaPSjXQCbJDG5ndUGO6I/bETaTiG7oDSVl8dM4VDhd8czTn
iJeF8lPd1KPLoUI27fqdCJtSCJSN7f/piB8uq8qn+3P3jjecmz/FGPkAHEh0ZbUk
jAV7exA3qIbkmVXjwcddxhYjkp7zvkkmo8HnwnRYPQfeqHehxCpo0Ziaju13kDlg
Hyuam8msP/AxJmcf0Eo+NNY6mva9pYA19whaRqixPLVmmw1Vg4c0M3O9jNohNEtq
hgBNFEuDaT4tVdjmW9eiPV3CQK6MvZc6tyQ9wnGu+RudqoI+MPGwuKeUS34GQ/Um
C81NvsDBd+8zDNqbx1BAkad5bDe/+O8POiXxdWl5rb2r7Rp6ygxh5m3/6MJV9Qit
cDeFtGNSQeP7si6sSQmxwG9p/Nd4Z22sWwi/GZVXMHdlFAACnUJulo6zHLvKJF0H
l01anhnnPpun7VDCeN4y8JmGUQK47dR6BcHUa23ej6pU15D41vMFIDOv88D8tuII
blMfUcBY8V56D9rJs/kxeqi1XvIMlDscEpSRprMANYy0eAPaZ7QDE2Vvbj0/MEIx
wGF8JaONwgfVyghBO7wAeHMPX99/vN5ceABxhmBHwwevt8vufwGzLey+cfwdphue
YU2gD34EJBPJRVMvt/1kbHHSXo5zP0vWglAABB9QMoUN3eHABgs9kYZj45iDqkO3
MeJA5l3HVzRbiRzd0dyKUHYRQ8NBRNs7CjL4A7qmcVrizG7LRdXWv5LD79SLs2zd
I+5LaBlND5hRAdy5+knvy3dDN1ekV3f+KgSArUdSKTyZi1zpYOK0qjZO9lwGnq+1
nYOdqWHxGAwXpP50ak23p4Z0if47CegLSha4k5JspSI8gKg9D7eTkageLLiUAGUk
q6wyAYp3SJguaDL5iE0ZBoEpiWg8xgLN+ld/6eN/7CrrW/+i1HKyJ0ieBtB7YGJw
ICDth4aU94RPQ0pQYYHLmA5hRnLM+/yGyJYvLM2hg8oZErLZ16A4Qwj8mMMacJVO
aUGQG747NW8F57vyZAdf3dPPmjOXYUj6sGEgmm9+Eh6iLDhql0WYua51efIQsFu3
QGHoYGTwvG9Dg1tf64ImhE71YlfvzDhdqLlwkgnb+g/TcG6XWHvbjTc/FhDhwu8y
/TGhg5TciXbBD+ax9zjw8wjDcNg5OOq0GqBYrPkjtmpOSRIK/7pCv8BD7/mOG+qH
6tekPMUvIzglSw9pj3XE9iydCD0h+tBjmuyt86uqdjzAIHqr4itIq9GE7Vx1o2E4
+tcUMYX/e2qu/L4ZA3bsqVZkvUmLC4gbvM3z8o/2MYiOV5DJ7eA8ssCobHdGwKrd
+doI8KEdwWI3aG1ZlPn18obiSecoYDZQh6GnMI+p4Ni2iHaECE0yMic1/NrDyTSz
gC4zFkNVTBLudUDnaZik8Ro5KQlFlDQRuqMyDPxyJiB+ueIxFxMv+JSqB7ViiFlv
Uii1kmc8r+C1auGL68AkqSYbj/0nuaCMC/1W7D7cY9RDXWuiB3zKIWPiwemsmbLA
Ztqj0rdkt7jOVwdltRPi4sQ42S9+04crJS7moVPJ3MAwBJr9s89yX/bD+cPqxxAG
RBSQwxadQJX/VSTUx9++vS+f6uvtoZ7aImFDYoD4difg7qwcZoRlKdbNpHtOWiPN
aBo2WvAXyqHlxjCEVqyF5Bpe3A3yGQY2uwO9aV/ri8KczBs+AXJ/K4O+BaEJggss
pTnoH/4GUnMfTvBh5u6ULfghoSayoHu0iicBkg0F3eEMQJVAXXTGNXyaH+v0aUdg
W2AK6EP7UmYpDCmROwtJ8bcVU/hVRVja68GbVvdiJJ6FeeOJU0yWPpcn7Zp5gcPe
MI22HHvpiJoF1khRaRxa+EZl54b1vxp8UiOpO3cxN+aAJfLZAK2yi3lvICadDtRL
dDEXqcUwv3m25P4/Uxc+KXNm/hGKYwK5MlUr3JJkkj0wl23TItGp+xm96wx390Cv
iXkwpQtea8J97HAIvNtXgO92DrFtKM7p+5O8uYxBPozpcdHvvw6xM2iJxA0u0alx
XzrGbIS94ntjYXh7qaNlnj4QUKZ0H5CTrfOSav3wgNnV6wGePz1zxvFYbwzq2Lkd
ejyt3GJyPKYgjJipu2G3ogqVVujxO1uXFMzZO1wFApaXRrCUUPlZdJnRL9HRoGqu
OH3ip5cU4mjzOPlFzJwn46iWOhxAPqDvS6nFi46s7L+0JIPSSSWz+slBhNzyXcCN
2uNApS9oJaQ9qjPW9rcpdw97+G16fwUMbymCeD0l5Ghyq0vUcbX+iM+Vy8sKU3sx
MRGcEEbnqiVrk8dObLYUBmQtm5QYJ5T51aHlMtxC2KAew3ULIcxDNeyheZPKrAWc
1jxTT+dWsHwIqELZN7xNgesKqE6s6C74lzqJ0NBpyiYaP6F7pfLh3BglRYNxbZEF
EVYcvQRtIgj6fUHlFgpB3yyF0uBq9XEaLhhq7cXCemLO0mIDNc4h8h1bj4rptYl9
Kz+TsSd6zhaFw+dXOj3HKmmcsh6Y7rLyeo6KuKA0ZAFpXOwrYhfmkuEB/cMm2Mzv
Y2GSDIzgYZR7vARh5461wqVqNtEPexgyhNPYokZ8AkJfwP8GNFbNov1IYGkiL5xt
45z8ZLW1eEGIalM9t+ZaQEVIcYsitr3gms2Tz+pYFjr+fjpZwH8I+sGOV2AzwQOC
L7tp21yQmhmP5zGETLyPSKWylm83lP1mRDi6iAgnAwfD8CBx6t41I+8V8BQ1LMe1
kB0gsDe5dZECI5AGR6mSkfKFHouwzwvxPlHptZjaI3oO2A0CrT5Ibjzj63jqpxDU
bTVUILT44UcPpRg9lAjTvA4ZzYXwzqKM7VU1YXhhFbE8R5E4w0Oj+IbJ0s88Acpa
fwKVVZOqwySPwbTZDV8pg8IPcGd5XUzJpmi91ai49ksfmkZKkMn/Ckq/m4toqByR
oKQGVoYu+AZM98QTAJ192hDPsrcdtoJR0kukpsACd/IW9pWXGW36KukySuOwEgIb
Ui/KhCAffPq1to11IPfrVW7x8N26FDyyAcK5mHQ6BM+XKpLcf9WkGE4vPi5ZvKcx
+NRtHlues3XNa36z/UdVJzEYlyeqbINKJddjWsWR7CbzabGu050TmwJ3kCcQL5vZ
ioqhEq4zvXuCVQl1d5So45rAPX0rrduq91yHQcY9T0Rmb+rR59uX6Aag9PnX1xSU
XE1Y5B8qnBw8qB06a3o2RZVFStT6ucgk9cWxmcWcDq7VNKi4AV28BIZ0KLBuSUOx
wlnB2NmQUnn7c6Ir6mmwKalO2NYJ7FEBNqG8GBWQVYi6TtjoAIpgyqrctJAW+iiT
lyQwMPoQY33eRtNIlaGcCyqLPQS+kmsbgRga3IKqXFnEldrJWNOKn/gFRJwOwY9A
QmZTbIU9ZWPGXhY0s750tiQgSn4wvCwNXN8bOZZHroLm/yW1Tu5DTwcUgvgVWcsd
4F/fqMOTMm/ZNGJQr0sWXeFroTbvJyxjAyaGSTX0FS44dZTRC5t4821X5koyPjrE
IT3Gx1VYrWQalMwWpVzVju6aFc2s2HhBsp+z82PAMPaKiOHbUkQbXQ9fO1wsgcmU
Rnhf9OUEWSfVWX3+SuGGg/N2AgdlDbFub3Idj6ax0SjiKSDFM1XFqTxp8aQw+/fM
wAX4F6oailfQo16AABdhgLPjhRpZNZ99ZbBoNtIw4gbLV3scyDUVj+ch9Ao625yO
n6Sy5SROWgShiD207VX0lUa2DYXoeHbYG3eafiX3c5GlgSK2Ds7jkanVyPawwGkN
iIFp2Wd5xIFzqVrRmXUJqHl2Qo67MfNaRrm/k/K5tsCW4HNOlCfhN+uAaXiNCDMR
OJ1DqRgMIy2ZP6Z536yUxfCyfGsHKZZSt4Q18nNWoYD2hjikwMOnENzCoIoHP0rr
jp2D1geMYTMzr1wV/oEQ7AaAGzdXXBZMMP6xLY3Ypxv0p7umFZiSX4xT9Gb9Io4S
VlPM0pNGEdkIC9qmAMotfhsev+41nqR//cKkuGLiiMQCgUmZkvQ8NPYg30nCvtnu
4sR52euB0LW1BmyLgMkb9aMTDIzwdxZaU94mbL3hyGpbxjhY4LMTT/hiZBIWp60k
Q4u8Bmy5X+3foZ4dQo1QDLrETxF8H+O+w+we+1rXK//tSTsQrUe0WTfMf49TLSv9
y6EiW3Lj2lwkAR3MR7bHV/P3Y0bagz6D6pNtBvXx7rSRwgKu4b7/+iGAKXbIVpus
qBKwdCHFkoaOlM1cEK8y1e/LYdTPYhfaDaZZNtCJZ/dhl7P4Wb9Xg27QXwF57HJE
Iw22jyDrKsY1xkDLmHQLNmCRW4Xz055eeQWmM6Z32n8rcqIDo00voOybCnaOjQai
qm6Pf8NnBlGB8aQrNL6JoMU/YZ+rhMIt17dLT9ekbGmO3RMHVRX/epu+ppnIupay
vFxO5eGDB7lXfKYxzzHr86fYRYXVkWPI0fSfFib1rUq66Gk0PnHTyl0+QhzTxUnl
eI+FtmlRUg8LvVZSerEYKA==
`pragma protect end_protected
