// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pLGFC6Q/BH0d7TWWQZeCsxGwFfURRsJ2fwQKk5dlQyYZzB51slRZs0ELvzwtQSdO
+ZFu3M4WNxhpRbamJXX+oBQDhkma7MbRmZKWRqsh/afd3rr18PziZW2EmmUjTUYE
3N4R2qTTSpZX5n8mJqnS2obl/90e3ZuRy8/YscCYFSo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20768)
mLRaFlwS24qeaXOM+lOGi8RRENQrKTqw3KpWI8BH1Yt84ZE716mJcpkaUjuG0lPO
NFAVmARAYVMyFUDwTpoAO/wMpFddTKwaSz75CArZjBsR9IHtKtczTVJgcqHBZS22
a8y6b1VjjgWCp2YfBDF7VSRHoRn9NUcZJTuV1ts9rJgpOae06b2gzZ4m36LUd8Ir
7Otc424xKGerYnuOfqjsCFxj650xeM3NdNeUzd+czbfb6JEYZQH0juswN3PnctBX
T4iW2TPnXwUjtpYrOeZKxVn4M74DBtMcHuuKV1/062XN/gIvQ5iRDw9LUSeEsHvD
vroRFIX9GjuVWV/kvopOBTLLZZpCjzf8KfPxWc/KXw62Cw0hqs5+jDRbZ0yjhhhQ
9ONoW0RMtOUzMnsiPDCB02vIWsCJVlC0jn+Sj/NMa7ttZ7LmcJnF9HZgL4r7ZVIb
a3xvS4u4Nl9RhXf5mGZHjwqy2H6RYoRF2yy/d0MrPasxmHE03DFG62T+Yw6ASndc
ZcV3L5zGCXDSDQ5X2gv4ezfzx0+fuWuS8n3CDKhtn8A35V9GGzUQlZZp2wnMUAsX
wo7COuFb0GumwQHqZxJa2vuCoCi/OKggKWQn5gMO+dG6SFA/mhN8RzvVaMlVFDCt
JpqXAlN3i8n0cFDbVTT8+iiOm6Ta8Qbzp07KXJy0ONP4pMJGAdx7H0iWoqirF9UK
xRSklBJOdpQZLBfh8uVTq8BqhN5Duy6Ks9mv3SO6mdxix9G4LKb4van8vwOzHHHe
Qe3Sbkc+4kHPG+Z/2CieZwmaCECVLi0cCihrDq0JF0rxrc3YxyMKj0dnhedFW2J5
NKUmibNKK9uwvQfjGhEfb4IqwrkCa8FVikZlrgBIsJ2yQx2jeXC/liqt2Nn+U8xR
zybBn9DYoZoZzLQ4IqCEDWNHDM2+88+6tWrVP0RWWk7oQxd4+oMAapHH5XymkFUz
0o8t6suCEcqXr4+5WVSRkTcCWpl7rtbP+OSS/+RxOPhPY2FRmHS6BAcAJMa0sUKo
AEkCrk31ab4s0g9asb3+B3HYQi/4Y4SlwiAKOrMLywj0kBHhelyzOL1TlLCwk8V6
fyyHuBhtO0KJAKOXWiFBViVBInjHChS6/UERrVeg3k9LQE4K5BqAgIuwlon7M9rK
58jxWs4TUl92gsLFwVW0i4bdlUVnsMWU5fOIlJiVN2Fkv3eNC3caMpgV4BPa/rZE
KzStZ7udEEJ/5P0aoR+ls5JEowOQPz08zQ60cTPIVyIsRhOru0OfQoLJGWb8B6eP
qI3TVVT3HwbTaANx01Swij92TypOm6jvRdfxEu7Kfx6SeB89ZfaCRqO1Nhh0L9WE
OCj5AkSroxFqKdh7xk63y8+SFkp8Z2u0gXz0FL1qaVVS/lfvWRMZDXF6ulXoDFtK
uMZWODHbYCcla0GLseQNn1F1TevLe41a9rBmIugnB6uB35Pf+4jE1FHk0GtEVqH8
WqIbEsE7VXs7J7+jZb6KuBQWXFuTyWetXO17TWoG+6hQxymQb+hsnT+Wuo1S1xVZ
YzEyqiKq97UmF/bAKoedl7bQrEZbZIXrJyzQf8bGRVn1k7yikUxony/ePNKnh/79
jLZyxdE60ajBNf/7iBDjJTzsQ7bXni5mSG7BapSueoVSewKe1C8koVU0HPRcOZ/m
o3Efgp6FAaoSrz8zrYStkoWgZYGv9qOtjZCqyX0ve0yKSnaTo835rgsqyQVIdftg
nxHDjbwePcHv3Th/jv6PpPs9y7DZAXQc7/xMuZJgyuRryF1NyeDzpFyK1yuhUbT3
7IkAlZFz9rXWxE/jWf1SjMsTxAdUbjX+PhGZWIwvoNg3P+Bk+aDGyr9k7dvPO12E
Y1osQtxgLYlgnlLce0zEliyTaQJXdg/n6NsNev6cEkpqdgK+kSb1+SrxmjXzvidy
Gqwr2Ta//yAN7+JJ3hwNXN+7fWM5wAqhkihTkirCCaoMOpDemKvrgLWQy0w6SKNX
E6qeHQvqKZfnAsF4et0zDQxznj96I5vZIOV03jsglfjBa/0/dLk/51QUnMONnfC9
VIVEhn35MempfO/k0u230WPLwDOmNW2zzX8uJkCrqYfNoY7noLYUroCpYU9gRu7i
cMOLyAFd+exZEhS1zZptyhGvTDD9wZmVly0yH41Pz2GuSTB514/CcLLHfaIO1azm
bP8ftViWGNAuDiYtI8pW5nGy8oiMF9vCPnWo7ffEVC+GggvecD/hpPFpdnPmCMTF
qOSvFQiimJPAbHwpFTv6XTPrm3EJzrfcSH5Pb3aVEQaUbMUvdI7hwol0zp/0gCHf
XJFhXeU8UkL0rNYmxNO9hgqWQuZK4RCMbA1iXq+8un6dUFAL421V1Cb6wrLdDlrF
+1Fvw0c1d4wCsFChqJ3xN9EhEkDGFxZyw9thE6uNFjReBiWTk8UDRLmj0JG+6YJG
jjFWEg5wj54eDcqIje5VaX2spDtscTddiY98B4EBcVvBwYTjJ0Qr37Ak7iEfReId
EO+hl1pNCf7QsBhArSXR9uouGW3JmWuO0oQsSy2kQ60KXJ7R+/Ik2xpg0Dsfvakx
F7+BeEQDsAVBk8lqXVpsQnM5iHu6DOETpPVRGwFh+NIcTFBoVazaqnAjx49pFN0v
hU+sA3pUFzKnZ8YKvWu6KvkdhWsw9tEPlWZ3fQEj4mUZZAJeCZcoIjW9pJgdBIyO
d2OyzEn8EJCHyrG2jP2iG8IbIzlZdRTbNOcsgfkXkKPQNArAcxwURa0843YI9hJU
gNcv4kTPr3/Fpl+oUZyFdkJWCn+rL94NoSzmzj6h0U3tc9Kgqk8oeb4hqHAzZ51Z
vnZur6hnk2olg6bYq/Z07iQoXWSoSbL/nUPk7J6fcfyNxWKJFw71Iy6Uje4dgjwj
cw4p1nqg/5tRwIcI9j6Fe3qTJaDXQmAfj32Y5z4pUmz//DUO6zJAkMF3QsaHBUnp
hwaozRUj6U3dCe8bJZyjYWLBYMKIQd7lqykNoL1dVZQUwJpQsdK/8Sp3SRsdo4fz
K6S7jk4VCGH8FJSTH5f2Va3uR84ic9Vu4/4e6yvZOFpxLoRq/m0plFBLLP2MbhSd
YKZuFkUCOEbxNl55BrXvPvvY8HQ4chHVxfypj1yr/FkUe6tusFBp8Tuxz8IJqxe7
3rZDr5L8PISos6WyVwJZlKr1nbhPqt45HvVoeiHPqYx7ULu3gQbdtcu9FyyWdGtp
hydakcweXu4aM45962P+mb5FzcVO/1EJjsrMB/ll7HoAhi7oVBPES8ofMaavHq17
PmAnAadKC0K4u9NlaXnvWcNaV4oqp+6VTZzXDILHUQY2SO7GMEuNh/mToYV8A10G
/cMEHgUeOovTjYcg/w1eMi8GApIAadGws+MueXWzJl3KBnBxHbZ+2UGo3h8DCnff
gNTMNdo1ZJO7YjylUQNsd76oGWdys0Pv2+++o4xFOVZWSjHiYbmMPp77zNWN8x7s
SpcMQLGRSlAbLNlMWZ72onjzwpxOqlz2Wjf++EjVybLpivyLCz+o/hnKSoehJGCg
VaSv3/b+r9RkUOUDzJ/hx6YWaF56d5kUEOi6y8e7LiNIy67emruoT3CsASMcdL/4
IB00KFAYMGVdE7VaWeeQAMW/RKx89sPpFo4z+6Ya63FMiE2u1VVv8iA8CmB+byP/
1t+s8LR/InlsSUqZgwgIZurUut+Bf6ZgxKCJlSWvOHyrkqqv2QzSkptQkg+rC0si
kkiNf2U3/zsbLVM9fGR80fFz01AZAFeYTIYRlv1V5rm0l+pDgl3TA8J7yNzzEy9m
k49TLCIupIAYOYWEA0nzzmTQEyaYzOKWu645UZzVTuMS8AcoHPFvxLJ1SmBQ+LWL
zzvxyWl4BpMrkqtJQ+QbLVYuR5Fz82L0f9o3IfWiOpOO0MwPZkQIWq69uhFbt+30
a4WqqogUVGqvo73yzt+yVlOYDdpHjhQHCmoxh4jFOypbDFw9nKIHk8KzUgH1vC7y
+iSeEBOWdZDGiQA36IzbVTz3/yxO5qGd1eyiVqhFNKxsEeXBltst4eOq2BX71SC1
KcheWfAaMQQZ7Ekl5ZUKu8Hhti0EXswMssiz3cMILpgqQ7K/NqmnsmMr93Ek8c8j
6UGUQs+VEUcL+2P+nCmeLKWPi8dcUZpzWwsRi2hTIF5Zaumn7TcQSCTWCqQjXbMz
FNEYGSILi/dOIIdBKw8vvIOIdrQhbXEvcnk8uRnDqewFLnQAXFI+CzXr3VBDF5G1
7oqJ/H9I++973KyHK87te8JGzV+p+AMTnT16q7vi55nyX0ojY20r617EZGJySQgY
Dqx01po2y2dTUmG/N+u0QA8fOCGdE2P+NRdvq0IzpI1leauML66PlJYI9p0PAKz7
dGLUdeor+3u1+JVltecUX9zvJ3JltD0W45FT8RplSnubdiJzoUAP+giJnui4Ujxn
41ltYT5vOE6sFw8BnXUJOuZBTVtpXnBhBMXN9vm2wObNkWO1VNBmP0imqTqraJp0
3KXVDhf49Ep4nx3kebPThaFTeG1bUg/8zA/y2Hf3QxZR0BgKW++JYx1D4aUbeQ4C
sruzhQ1NSEyx85hKQSAZFOv5LQ1aX4OJ6qMlhRP8VWKwmuzlXWYXHso98rMPvKzd
a6IQHV0kl6wn1ezcZy8c8xZs6M4Zy7xZ1p1Ud9St5ygjYSgNGk/yDyBQxWkowZhy
QuqGhArHlApUDTXcClnS2gKe8HocNDYfmHUBvT7UkQ7vseDGF4i/9uaSyQKIzIOU
oJTHd4c3J9Z99NabIEsMkAa+GkhvRHpNCr5YrdGs0waaW0YChBtY/r7RFoXPJZIC
HviMbzIxnjcDclYZiwWSyeOcTALD2jFicr47KMVSO+AkgyynOwovFHuo8ys365mu
kzqvuLcpFJIaBtdCRwMxQbCK7m6HBMfulD+2h1MpNB/sRRMRRBnhFU0E++kio4L2
LUQrLXUql39CwABFoZbiX8yn8lIomze2iQth8oJ1sa9yfKDnaE9+A2P0GBYmQosh
EStcvBFOU4G0gmcMrsmkD6ueMBkcEnTbHJBAwtdKyx6PzSpqMR5un8yhKe+jwHsQ
wdDxvwAbzY7P3QdsQxMGQpfwRIWPIfFwsgI/LMbH/71PI3mmr9kWb/L70yflGQH/
P0eODbMG1JfJ18lY6V1U+2NwWWI6o3OkSbg+mqfFEP0Ayqb/+Ymn1TOlLn+zpis0
QMUnZ5HVNPfT62zyOc1QthYf7PFPj3HG1vkl+PnYwhrI5uTThTpb9QZBJdPLpuuu
/BjJgmTRdyWVTZNZfvGHwbubXHWud8ddQqYJxvQJ2/HU+vDdk9I8K6Y+4hWPbnC9
Qe+QIvsddcpRviCzeImW6SODZEd7IWkSBq1mdlKU7o4xCy+smjS5ZKy+RO+kniYf
ZBnD6b09XM6EarndiMlZBqX0LnDDXTfQxkit7EQWh3Gw1KXTqOM36wBHJz60nEsb
i0Y+5c1tPq7vMbP1obH+W7DJcsxvl0bbGdavUWvswU18U+CZc4LCvdV03GNhAmFE
WVF/5GjD0O5WevTgLTb1XoVEuTRVr87pbwe/7vLuAT4m0RBMuQ5Kgwa0d3FU87Rn
jT6IvBxREb8uKt8bd2c4BsO+TAtr6TqMaKOMdAztTxSvS1q2OSpul6HeJ8wllPTx
RqA9dB9K2e7W0QFius0S+dapDZgTM1zvDGFq+fp5gxyvXclmqxQ6Y1LLuDFSpY7Q
sACx3jmRLu9SXmkF83CkdfzwpwC/FW0sKEKRUI0amGYXX5mPlW58fxYju01XbYcA
kyKyb2Qv+AyLgaR0xZvrh8c66szQPcVHFLyCY6aeYE1GC1wvTS6VwD6Q+Mjnz6Hs
dvAWr/TnYlptHsLtQ2COIjmw3IyQ6BFfODTpKMkyn3rqWF0nkB+sTi7n00D5nOGc
zRQH6TMxNaXizM5TAMwQPRlc1trwhqOCU13qNoNAVaAtcy1L5epddf2AdT0d6JmS
LoSXvh/N6aDUQLIDEzFaysZtmxp9EbRB2UkvpWmde05BffFEussZF8IX5o5IRuqr
uSgyPfhrt+3zy1lUU0WCod3yt7DhhvEgaJ6x2VcjECLf7qh2kSNyXgZXBEB8Qk19
LtcvP1RlAir7A3D7ldICcRjXP4jUXq0VUWYWkQymPFFD9J9N0Keoj6WbXnMnkTdj
cxcXyWOU2uJ0xHls9hXxU7qCRig9I34YRhD4SEZ8YRkl+q1SPkQWwEumAwnDm1Mk
mPO4R3H96+vlZN/OOx6cz0gDsHGhqTVH7YIWMsBYn9kOrSKn30XeLaUm4tMAqTT+
GdCGqlSkGlaNhvbW/XtRB5UuhUPPKrFM7ETzEfleCy49Qnv+RnH6tqk8mLva4npi
nz6pZzxn+9l4Wob3RElrzSaBiaBiuNE7TCIgo0LLvkaqGmWNaajJxqP50A62Pg8l
Ng/5GqAzUl+X4UBKAD0ssB4kndR2buvK9OVrqS4I0RhBmEE+YlMp+u36LSPpeHVR
Y2nQrxm4iH0JUXrShlSvrEm/HlyIr0KlHGa0HeE/NzzmiIZiitnCTxvS5ltdFQq4
TAnIPT5vtb+12BFpc9RKdE5YAA6RNeiIt7dK9bEc1I3Md3fsk2BGIRhrSsyz/zZi
GfuI5Qb/Sv8X8VKvt7whcnTAODrmMtHnmIR5gWa1WFlfbwG3Bvdvu/sP1kGQawhS
Py4eEjh7Ln69gX8zZONAt/NTB6VHXdiSTGQ/pIFEbxDnMjkg2fnHSKVWf1LsJL3J
bVTJaNfBWuohAhCYjHY59mhSUOW2zMqVKwDmh9FzLO8ovxOASo0umDSoLmjzisiE
0YPZ3x7lEYTMHcrlaZg66D4tIdZXgxlvQ5/uoyxjZzd+Htt79iJWLBSMs114PYuv
il+c57HWRzvX4/FBH/DuvPglMB31DWoHWIQZvwEINHGceLe8/C9M1+DoGOac4+Y0
qwCRLLhgSPoPnKZKMTo2Uro2jyrKEjC6mZZuHInfnKPLtxyqTY4kk/T6qcq6Jiyx
SDgqWBPEDFS8f1P1fN+UsmGgamelZ7cIHkWewb34EY+f08ftC87vdFcZWsFsPcPc
MIUixV+8nRAh11TpGLTri6PA/fhWyO0a2nX6w6na/oOzsdDzLoYHc4xB1lKjdtVa
7s9C+doDdMof1+lAMia1tdu7OqidzBzVXJcZlFFd6tD6nHJsqcnDUd8yfvDDqfZQ
SDZuitbZMrOfmO3Rk0XAvQ3qLeTZWmMeAZCwcMqSy7l+BwISUMjcizjf8jQNr+je
MSQ4i5SjnmM1g+4vbr54+LsnMis7hBJpMmaNiCWt7fw+ovQ4BvWYr34YkZiaEcRJ
CnQtsh3nHhPaEDj0uwdH8tbkhc2XNNs2GW8Nip706P7biYYRi+YsIyMzgbkOu9Cv
cT15E3qQwy1Vx3O6J7e/o55uTvoyereDoST/GdqwU4wvNB7qf3MwSTQ0y8JUKnGP
pFdRWpOMg3CLoiHH7Aaon7vUk4EDOWYaDa/eo58Z2CxUv98FHMo+48nnwQPf5eWW
JzLwI/Z4oUa8FjGA7ZwYm5lk3HDjUIVqRsE5sZIRrvg/lm9YXXcYS3p7eoN/hwBX
Mzy49OoQh19/09/zVteTSYFrNUTiZZbBDAgtBbJ++CwhAi5dVzZbY0LIYcLYYplD
cGcs8cnkDXcmcLiF9bxyYWnScgxPyifuxOVWXtwC2NjPE7VhO+8xzOHeh7zk+l5A
cx5OaG1tmP48UNj+OlwHUGiMLOVMRRCQePWIhECm270D27q0VzX9v0dMLBrGoIak
Dl9R/LANEck5Xdig61CH8fYxJ2PPGg0s2vumIPElc8QvJ6a2oBbP4EMiYKygfXXh
OdxA1n6rvYG1W6eqegBgeXP7w6CQp5pvuiPnxKgn/8gXZjxJ+F6mOpIEUPM5hs5x
Nqn+0WN754K/t6nk3uFseJ0YHlppmObKURGAY21e09BY3D/TpnTbG4vBbRRylIpG
b5D+CDHL/LwAqjQR/d87vI5stTZV6ITDjGraIrlH6tH6Ow41sQcfhVMpuS5CpFwy
P100aoNHXchNVAH5G152E2xQQ3M9CTYh1hlEVKrG3YIw8JzvSPMsP+RnAaYvTrX1
dq2vbqv8/ALH605M0jdhE2/PsMyme5Xeqsu2ahP+lbWtmADnaiMkDaJxZZfoltA6
wz4StKoShsxzYDKWe3fm6EWw6bTOdXmjGlPzUBFVizl7rHrFSAilTxE0tmwSLxlq
Wu9DtUWiWJmkaLOEyurFYikdxJDooGIqx9kkJUwBbuWZB86OJb7tSmiW9+Mv+44X
PAuVIn/Gv0ipXlY/vAqDEIVOUfDS/Vno0QEXo5gHT9gbUqT8RwvWU9uoceVCpJWt
oKcE8rcUYkC6E0iM5N7dgH32G8u7i3Oefd0ieJhJe/wUXnMTjLLFTAeWzFR9ob52
MnM9wpQ3puVaokGSkx4/1mDKf8PNjmM24JSx9eOmHI+vB7YsNHyLVovkjMFwhF1X
ugztl0mte3tHVX9hAvqCWkY+8nw0qEx7bNCX+6etYNUHL3VO+YY8Y6b8lVCMWiYr
vOzZiPIVtQ0OjaYSLkNlzL9iYvoXt8R4HXLqPa8uHNgwLtNFxt8oS31O+TqxlRuP
KH6dKTSnpeD9Ayq0O3n/1Me4w7LIdzROG95QSPSlejgKdju0x2uVptXo6VOyzk+l
DaMd9LFhmOdBFzSexT7jOA6EYd6hxDZ+X/wu1pIWDC1SuJAk0YQZNy3gYz4ieP88
ReCiBkjjFoL922Pkh6Mod2xYlUs+QcetFTHEEtrqsO08KGif/r00ntKdjTaRLdUH
glaB06m9RLxcU2i2/77dl9+UEFG+5cgdl8xhLJ/rJ7k8+hGGe6mS4Xptq4l4YYOm
JMv8W2fu4TqbcJvAcdYLt7BUHK6JMDpBxC/YsK/bN+bnpGmd0jIVqTdvZFO2N/5e
aprI5ZLH+KVEZ43pO2Obr83vh/fOe6ptTYLV76NpPLJ9mmouCX+PHXL9vGedPxul
sRv+NntjxFqGndOkUWgCyOnynls7xwRR4HG/XJQ90ZMGYgQow88OGB9NGo4UxohS
UUKGaYXuBw5EotgFZSOfNJHZarGe4tLf4JuuLAesmX8/potCVefSAxhoAqXNH20O
i5jM367+hzRv6A8Ja+mQjwH82YEpKNtdclKsdWeUHu150L2hUG8YJie6CF+rRcaH
yeTM/Lmii+M8gOi5+CWIQ/CdQoxEQtbcaFuW4DkjbFZ8QxSs3sU5iwe7k0BoosfT
O85AQVJODPKPNN8S+uiLfW9MRAKBV/MNgTZWI9ef+wGfyLE7hWBl+iGy50HlTHav
CieBtr8yn/XwJ7WXZNrH9z51QLPrhjoonBj3IWhADac2DDvqw9ihmSeF9ta9eq/8
akbeQLQXw9FPLuDuFoRJHaMYExm4uLwbnq4n5bKaCFUsbxGXpas8YzAN0NpjAJ8U
8cjm98ZrQlH+Abwpm1NonzIKlP+jSg9vP+Ndv3xMY/T4V3OkiNpxg7/1CO/B+6OH
eItzXNO7T5odXzXnO+TzjHeqYExAVAVb44WMVzzX1CHPBQXaxAkcoiOflOEt79j4
P0DlW/pdPaPvaDi2Htbtsg9L0YmYUQ5lo294PtPwvSTL6IWClUZXn+0RfCq5Yz/7
S+MadTKupd9E8VPjMJnsLemIwif0+PYYmLW2MhBgT4fNR0GfVYwQGn3nT5HY9ymz
ehjlTt3tQJ5SKBaojq64ZTe903eFCOMTgZ4MmDjkjUteVxX3slJjyh7W9n95MOKD
M5hLneRFAkfQIh0VYyD0Nz9gcv0r2bAfNTyJ4gvk/eBM7eNPbjPLfbqGP3/bZXR0
NPEgWcCO3wRwZYPZTjlGYfBNZDzXE60xMHGG05MNSSTIxGG0FNXCedpIT72fK9u5
iaSi314R3N/CXAGgdM7/KFzLsjbJLaNO1HHiP51+kcAV6QCkA+n4Xct7ovX6nIzJ
iIhFoiv//eUxCpsmc58muLLfgRSp/cqkkD9KBKi5NvZXzYBRBku1b1EQh2RjwcdH
Q7c1rUDSigNPQmhXE4xT7/PeNS024x4oSKIbSAfvH9xifbjoWbZiF8Zqxev90fjm
eaSLDgrv+UWPaREuKGmLKK1o25WjhmPUwqX7bKUoBLCxN3kOObIeopRZc6Tnk/V1
7ww/4DEUSXpVplvexb119Aw7Ivp16uZH9EA9nlKhtoaejEQGpxkljsnj9bi5liCe
i5tdrPaIsgyiyF7XEOwLsnLqECXWJwi6Hk97BO8qjhXDEZYmjhgarMmp7d3jzuKr
ui90+PmNWjVxp8raKQo+C29T1AjVDTmLcFJeJtyBJW6TNbpWeYAvNJJcvSa0DUqi
2sycFpsUw8cuGGn8Cb+XkGGRHqrC6HUyIkweoGsw2c2AwdfbMtyRVMpokg594W+U
mLIN5HGjp2yGFbVEZh8+2CNejob1rnPeAJeGy6v4kPIQBNms734LAPgXOLxJhI2c
WNcyiy19P03R+grA5w7myTmR0tCI4mG898RyULmpaB5ANZ7YudnEvaKslb7IjObM
TGV8yYX5EbqFkSj81FsYaRYlB6qlFPo8+A2rsw5h3kFk5gwqlSkqvjfLw3mUiA5v
m8seihG1yoJwmcrv1Aa15wRs15K0t4rdILbKsJFMUoPJIiRGNCY0+zfIOYSfBjsL
XVpPbGzaeudiT1DFm6WY8tOBxA3YzZ5bGS0MSrT6ioBE7wN7u5iVpnXRXDotPUTp
wzdxj1LApsnli5FFDt5BOSoTnfmQRMe5eIjZqgoPRz5C6Yf6Eu628++AoTt87XzL
cmV/TyTjDqpN+mpP7kjStuMaocxK6IZzL8cvvlTG6XY1KZUmuqomeNqb4nrDDeom
ecuKXIZCYNTW4vVZLLZKq41NgxR8MsuMlsE9OofqV181lzJ0RqVgMM7BOurUZR8m
4t6CsYOKCLONTV6zEWCnuPT3lQ72DSYuQiFYRjJOfaDMz52Z8TTgn20q4ENe2SEN
UJ1cyjwaRGQ6XtqBxaNsFX1RxA4LBcuT+RtaMsgSkbF48RUDsTjIVcb0xcoGAc+5
EiT0PVR7MigGmvQty4mHwVKPciVPv581ukUdKqZzXmgA8dUiFrvfqMjPZG5JKfSP
+uwpCCV5e77nCMcy3foPgbMTKZL+yljtpXnhYIt5WkxjdGfyANpQDK3J81F7dan4
1Qa2K99ry6C/yfb3PNirNc9UxCEGHsw6VzW9Kcy70lxyW/14nGerujbA5tfedSWV
zsDGY8E23itdcHTvfgBSWoQQYfU26Yf5FWF3FuiPsBw/EJAG64FNq2s2odMEMfta
QfW01GA+ecdc+ic8S6/kngyUaiejvz6ZhSmuo+rGu2usHrq1Jo/AZVeuac2EJjJw
92rHy6b1LOOS7gm3+wCCCQn2PFHSgmshUzJ7oqx8nrT0QWbkDSVJ72L6kTvr7/Xp
BwH5nS5VLVyIycuZURtk/6IjG/oSn9dpxw2l9qDdrouXH3ZmD4v3AENZgqoPu2aL
JXz/yIInLy2n7oiGoNpHABuwUjElAGx0PnvYDYQYMustnSGGP+QXlokwXsTLZiei
Ou5S4JDmlwuejFLSrj2b9LUDjvGTtyEXKP15muESqhiyz61tgFa4808oDTHxJlAb
SrRoJUEV/sAuBFgCpuwFf+XGY0nsyIlTTuJhofE72kUqPIxTXcX0twncKPnplDcc
TAOY1BVXFbtyHZYYJWuUBpaXsN/C4Gxy6yAOX+1nyp/Zz1gXOQ4+VZ7kCoCa0jHC
u2qNiZYqcSbuIrLohU0cd29x2841/XkYUqsp6x2QEl8zdqjtEFjqc4toGcFGWRnb
iJGHirMnQArhr0OGVV0ge3ydWfopU6saPs2J0pFxF5bY/kvwydTT7IbBaZPscZK4
ZQ6cQx+3z/xVFH65IZOG+6DcSq0/f/aw6IeGyLrjGWjQKPZaA9FeJZrEy4NNamTW
t55TbPOPii52knweNItNp0o9V9hxFtQllpZGribHU2ezLuB3QdLh/h5K24y+Glvo
IQBDb1/J0RcfVhVxoqOkZxiShQnihKC6bvoytf7l11csxaMXzPVnjBrt2TJktAz3
lfsp6cZCv2t0STURHorXs64YjTxVWieOLWgz6+zEevjrVwz5//3byEiwX1pBQDyO
khYjiH7zk5hV6wkajxl2ouXt4NeP2T4MrOb/tjZDbc7kBqcJoMEzfFy+id9Q5kWE
7e/3OIUpa02Ol9HLJfPdfNjRD3B/KFh7FGcGdaT3Id1UGmlSK+LwIIVHe2kbd+jS
g6RaG9Nl2H49A2ipRKDqCR4F5NYXuRUhxVKHdbbpl4LqtuCGPf+eeEYSCoOL5GNK
QKr3McMxZWbbNFcI6mVP62k5C9E36irmFzyMiAVz4n4ix7RWu6wxlYzKHDgKwUct
bwButIzSCIsHP853ydTYfEY/bKLAukCy60wH7b1V5wq8YKkXp9gIa1lGt+iWSNIT
DzqEhWFnInS64a6fOUCCnHI2+BHghUk4ZlKfZaSU9PVvliS2Bh1NUwFa8fuZUMtQ
wjY0kuc/HSwLxaWTGWKooqRd/L183fgowaX/FHfQdEXP9wm1vaa/7V+vsrqC0z0W
dmMmTVC+9mUcvJKItZriqCovuXn01c2FfpkZRgdgdKEZVPTkKW6cg9W6QUL/hbH+
z2HAgL0uPVrkWSAMszA2ltd3u3Us5EQ8DSX3DR4nr7D8jDdfTg2p/YgFfjuFNVcY
xUSK1fiQwEj9dHj/tJWucKk7VkqpeGihsGN1V4ULSGU39Au3pPA6/Z5oQZ8XJ4Wv
BHScS7eQy6dr6dlhnugq4sQA1aKTOnjZc/THHAEsB2GVaoFgdbiotnnYEtoqeDmY
4ri0wFRzU4gNMDeFDXn1Rjj9zvbjqZOhN2NeuBgUJxTUGdCC1HSilYUOf+hSsC2B
IecoBp3vv2XWlrNER5c8jjh86XFCWRCx6C8zaD8gFNI9LYJzMsm0VLbGC+gSvH3k
T41yuHM8RwQtvJFsOkTSaVqjzn9UQtUhB+n3r9x9xobAddzWdLFuob9sUiw86UdR
ifs1QcqoI7S7uNSExiB38Hb8yDf7Mlz5ScILVDTNTwfta8VLfKmxlblnRDz6uAle
QpKLv1R5hxxkESFaJZTiBjO0wAKNlp7GL0lE7QmK0Yw2gu92aqki+HqORdd6TSdD
Dndb3OZIkeLI953Ov9s17WPwKy4zhD+Ynl0DcTRvYXhTLFz6rOvmIZJPCJHAlstX
A2mNnJ4O9GdNg2Oy9XzOC4GRt4BPmOBJ9EohZf7ADR4Y4DlrBuJzw2nr7h2pDxhj
M8zD2EpG3XaQfryBj2Z84K4FIRZERqILhCGqUU3TuV/zSK4Yry5pep3Ig8lnwH39
aX1AmvMpCh58UoorYMAY956VWv4m9/LfObFu5AseL708kxnnxGfnuZn0zDvRbMRU
U5Q/N3I5TjWFCxL83Wz2VXUM3mfXMFoTvJ72mjELPg9UI09tsxEXmLzXD008qUZ3
5EctpySlkcZ6FopHo2tiez3QQ5nR1GNRH6fpY3GSszdJQSWEN8w+M4ktCQAMMKjZ
yFhGr56XvPJNrepNRmZauvOZYtPmejf/tzSTL/NXDkPx9pFPupaRq1Wi2ZyGfN67
N3feOkTWhOFrkYD9efI+yyPbImb/TtIFbM2YG0f3+XlqcbrjULV6DXbdEax2ydo7
JXypQfUA8F82sYiCJLg8XWS1GAqoTKgFzFNV+QpuH2rmbX5GwQO+MhR3JWJ5ug+y
oW/jz9U0Pu26n4tM2dpq7XXtdxX64HSnpGV1ulYTCxsA5dXGcSxTcEWYYlnAwGiN
PfuUEefsByBFTu+nMuJuBouJBXq6b0YVzCadLC0AAZreTYeTa0H7Rbxkk58/67DU
gTSl/o4AC+1QOPV15tBy4ZqboXFjvWs9+wcRvjiidzMl8h+4XL5zMsdpVplfN6tV
ofH6I/pS1ejRxjtp4AKiLIpupGLwG1hooZQdsjSpTfq0RNxORCOOs9TRwumcl3jH
kauloNsR5i3GSxbOTc/LHHp2/UrcUQe8EUwqMBP5JCsDSmb4F4qzJ0EcG0NhMptj
qQdfLM1bPjV67gwTYxL6exQ1VBXxK53SmNEFt1PgIo8oukuaD0XohvQFpik3OEv9
xCr3Wt7FhNq2Kppi+pShNEXpLJ9ZMiEjirMKZQu08gEJwKsenEfzRWv8vz6aYb2C
eAUh+Qyz0rd1FtRuf7FF2IfUxpsxUymK5c1z//bvfAsfPtfFJtbuLO22zyiPEJh2
wBj37nKmh41qfU+Pq8m1ZSwKlpmDYJ0KtQuymgQ33Jh9fL4XVOG+YFaQGlPatq84
MothHaxVpRbNJ5vbWdgotAjhXQxk7PAQ0njagM+zEwKYwddXsfXLxmAFGhUFJyDK
meyGLy+FhMwepmt2DP9rwy0Z9UplO4IgMdFUeuHFu+Qg0zRK2HV48dItT60pZD6Y
NbmTz8BLIrFqotoLJz+cCCXEHYriI73Qc8bxapeBJQfGPd8iwe4CbRtiGQQenWGf
Wo8C+Kw16hE0+t5aFymuIEyuEDZFH+1t15eu16vUvBlsngsJfd3jU/AUgzD6iliM
O6unq0ot8DF8rU5HYBVKHs47dU9D6ZaTlMSnj8F+mXscssgiABZy1xFsEaJ5zIq6
btnLdHFLwXThchG129z3mFUQ7/WcWfnJ76dmDlLsteotWP2qgjSnE9HHird8Sesi
3Uf4mTEj4UumDzK3LrxDi+JqjWSDfmN6u2tUsmXDbjESQR/XMOqkNT+ghv+yyQPy
0n12xYzIq5TSb+148mL1cIx4PLOy1LRQzReaCODpwFmlKGKQDodd/jXmSfrsDYb3
oK4DEmVw0ScRmF1uP4qXhXcv6GU1MlFwt/b6AsYPSuQUxhoxPY4rNRzMYYUnJARQ
ROiSd1uXc0MWbTkX3ivbreu3hRn6KtS7YEeK6zTnPNmC6x6na4OuGNgifyYNNuP4
UJPTQfzlDrsMWbaDtwcLujhmwnykoFdrpQ16vL1lrpbcRGKVeM99LK4edvrTsRPH
4ZnAzzDfbWpz7Y1CuZCCyXcaXAZSOMzWYqYub9f7d7J3ubcbzsuymud86a+ZKyBZ
wwOwkYuxLOKExJ7xLMkDZIoDHo6mbq5H4AtWriW5mKYZrV0NSmp1UN4N7l1H6ElH
vRG6tAwbHloewgfZPkPaLizVChn/02gnI9rFAz8Cw1SzN3CnftW1XYcicpQCeQx6
+bhp7cM6yZpNq2jdOdk798A3E0GqNRKd+zyqzAACcaTLsbP5EVGt87UuVQ8jcmoy
GkuX1e9yjZrl4WLmWDLzYydUBGFSRWXrJ9G+QEKUHnOnBAZaepWTwBzAUOmYepJl
AMIJDKFnfw9W/frxLZvgnpr41SvW92ydSB4sulRkHFuQAj53++pero5osP8iSF3t
wZ8EjLMeZzSYN96CALQ8O4yJtkygfa5qvXyvtWKAo0WnNaucZqt0DU+WHw7mSKnw
XaZccQq4c/eoCrOG2GU3Mrc8bkPTuxpKYIxJC8qioYjD+M8b9dvNT7HQ0qeCgu8O
lD7M9ZnLaJkyJmqtQdQKlJc1f1lp4nm8w67HBx60TaHoFHxc6jX16jfwCbCbjZ0V
xgGPUBNg7EUP6aIQxRYg2hk5FWgZcmOUmuIm3x2B4d6tsXrauXvkR4b/oNrb4/Uj
2pLTJxXRK0KovtUmLJPKMRlP1+PEdT2HoNVJVcOPb5zAa77WboY1CIBaOosfG4JP
UeksnZuSkdt2EkaUgKlqc2M/G0TP0AN/6yFzQPjPnEsib5emP9+gNImhUOHiNe54
cgU1BVNK/JuGbCG3hl9k9SUEaiAhaKWi88UCoKgZw3i+jC0694YWJpV/hb18QYg4
5c49sY0qvt27kzx71cqIjo3jO3Djwe5+JDW2mUVkZ0aAvHGvzOwM2I+SOGnVsNMq
AdBIo6e93oUdB/I9HwxbybU/GPrF+UvXqYkMcekKe7tCjLroJrkhm5EnZ8IkMZyf
0a2eYL7fRuYVOHy3a/NkZG6on6Fvp0gDIgecsBlOkRWfXNkuvwppskxd1PJiG45p
XMaeBX1QcmZsIIjaR2c6HJkF3YZM9fs7Fxxn+SqiR0N9kAMv+WaTXSAefXtBgblj
uaGaK7//nDoXnxJwdmW2JAenN6TasYm2KQR4C6AC2oiH6y5e6IfZpdVR/Xcj3E5i
RVAqLyMJqudfI8heXvfG4niEuxlTk6VZXDnACYh58u0pDHO9byD1ayjjdLyPFkiw
35aSlk1qkqXE4yyfraEWGoRhfcImLv1sO75BgvF8j4holtdvO9tRdf4HU5tkfpHz
wppTkPZEkFg0x1x3k1LKuBZHz+uMn/GE3iFiDwkmaHdgalbIeiY3eDP7UTMTiIHo
xfPTvJtHVVahjhDZRmZkZiovyowk3W8lBhdKU78D0E/lHGeQXw5BfoFKvLrt3TXw
qUlZf9hTjW0rnTsLY2Q5TBLYCu9GyAKXjUlmUEXHS4zZfXV0JyosDoyyw8Qc8UIG
WqjSAHWIb5RcDEJuebsILAXkT+g8GDqS4/9F8anp8shE7WDD/ky1+GTPzBxvDiju
ke4ms1ST+AJvZpmZ6OpM1PSL13fjN1gL6cKQRpiOxEIH/jkJNPBq5rhpyDjontuH
MahFN7437+qYoxIXPwM6iqOFhcZQxImUiPN6kQ6hC7aM1yMjeSnvHBs6YxS6HpXb
A6K3bYLIIJjhMEXqwlMuoXjyV51wXz8i+PaLd6/H2PtNdT2wKouwwIH0IUvZ4uyI
+CBss9uXQXiygx1eJPjIQgvBQsixABehWnDrmCs8zwdrJZQylk/GTbQneQp4dFw3
kfGoISXKAJKebuhlAzyz5M4pFzCQar5MuJU7iUA/yWV4HYz3fzolebW80emHlACa
21Up5N1yyV0AqOuVsWRCCyvQmNMtSYA+rCST+rgtZ7tETXZQ5Hz8WEscf7GvkbAV
VkmQKiDKDul8+g+Y1pMld264lKQHD0F9NdZ0q9f4BDht/kwfGXSwMtFIUUMPwiIp
1hsASAtdYhZ6L+O+bskZsn4hH62dWnHPV7KuFBTTUUyT511vOYz9ejhPd+7AVtJw
vEaFOInBF2Wn6aXJUOd+L88lF23wuRkNlzvSdeJ4Rzup/0v8NzquOtNbsou37zDY
kD872qEHiAtQGJKjTisWQ4GJ+8SqY8CqG2ElYzQMX5Z+2Dr4y1lzpB/+hVBa2uL5
rwvjVy3QtRF1fy9xZIhzraueTaS1uEdnunlFA8uVxoze9Iqf9iM1VmSk/gQvX0nh
9hZZ6NoiKKWlHKIkEzPbNEC24gYY8w5wj14LGcAFJ6woL70vJFYJDomjiWsSptC1
mUQel1UVO3ld1qICD2dTGWVesMiyC1Gux8vDyYvxbYhiJUCqBnUtvGmtIalN1m23
LAub8PBvaCcz0VsQn1iFbehIwjUZCVttUGbJW78g7ptvnpY7c7idUSQIAXSiGyIB
vKNC0a0IVfPCV7T8KBRZiB8hGDWL9FUx5RHUjOyubfBLM+TYTDusZRf1FVFeNyev
k1Su9hAwF5E8vbuv9pvnWWD26woOPzOukrfhyQdsVEUNsTLfJ294hxrnklvAfHSb
NCsptZBGTnWRQ8FReYOSF83EPvMGy1eSlZ5kq4Bai6NpU1MNvE1/YHEnnjiYhO9h
NPgMQLoNouVCeNqyEVYanXvJ8Bo6JM5iZK4or1z+T/cXsMmJcr3MsrXqq66KPpvT
Cw9kFrQ+mzeZvw/jy4Ws9CyROD5eq8KtqFEvD05rhhzQU2jNuEgrJS+XPlaL7Rrt
XI3yXaCtY2L0y1HOyHApYHxmL9DeUoWYWWQ0K47P2JtcdcMbEGnjGA1rU6LwiMjV
vktPoQDwHg+NQn6zou7mvMx3W7GbofUGd+7eliWvnC3CKyaKI2EM84jXcHCpF6HH
FysyfweggHlopPLhRTmI0squn4zMV2XTYInwkegL5/7G59DJ7zRuoXE9Lrmd7nP2
jycc6a4jTsGsrH9VVM6tQMXvO+Eh2PV0pE0N/0I+tWL33NTlvUEQtRCM4ANFSn6N
xTkGTsb95Qu1W5tT9cChU6uSo+5umTRBlKqPxdfm93D4HkqBogqEVyEqKadg1DQA
qcvdvCdp8eKFvTsqrdHfaWmQ1Eh669dqoydbL3KbM2IyafWlAi3F2Fy7Ypy5VjY6
LZx8Tlp5JQi/W/Jh9mvByZDS4wNqZRlrD5K9eCdQE+LleyBS1et4yFWKHMukUlmX
KRrH4iDNGFcVHH7LV1qufpxpinmQX2frEWHaK9BxWt5N+w946KQnCCz+l3JKzLKR
nNX7uMYhDKYEJ+iN0LMYRBM3knUE010/48L4Oug5K6bt2BEuLb9qMttjGOhMegPi
MPmYDM6bTI/7DQwvUswaurElVAONZSt0hMzVnEukW4WhgkVDiNBOmqXLJRyQXIth
4KydH5xtYFYTtpJiDb1BQixoOdkDZMhDSHJ8XGEWGzIpjhPuIcvThGP/5sQnNYHH
jvoA2QU2Vq9iY4OgqJMg8gyp0gJbVjX+0vP4SO3+3RQdw0zMloJm7vD90blvAE90
Da+uM56sOL1bRZ5VM9o0yjFIdCrJbO6niejOWqWJtikNz2NrKToLZkAwUmt1SZ0H
Kv2ZslKe4mOpvZvbEqJLYcHNmaxgifGANLKBGta9CoHC+61UK5DbrkVT9rzdsVrU
zEn2Ucc4x07cWIXpkxvpz4rxZUTQes5y06OvVdjMVXZBnqXwdZs6lpXYIQTlCxey
1g4Yge7/7o95Va5upf4Qs5BeuiiUyRCom87xfkggLAbsjlQoPnPzFTKk29nE/d7X
fZDVhkGwB8hNYoGssobL1ACoAcaFwahwkkdRu8neWwLT3M86GgsKemgpY7KVRp08
hS6MIWCqhT9309b0kSIU8C3hA9VfibHLwkSiTlfHTwlT/yQwF4bubcMaO2CABZsk
yMGpnyLFUFUgEijLhhW48OREZdjs3/bc8m0fb5z1ymgRkqqwmuoxodoBDWJ7WWYK
V5ZNhWlJGSXC6E6gl+QfjBsCPriwiDrqKiYS5VuwnJ2m+2NF6YqkkRlKIsSjCx7p
38/BlGr7xPG5ueD0ietByy1bOVZtTDZzGW8tB1RDmFdh+QzU2FaCeNIAYbiBDWEv
LJVyq1ZRSkh1WXDh5AV6T70xJup5O3w0qiY+ma4OZRDt3E3j8NBm0mxRD/J6Jyc7
VLmJr1eQBcbJYxYbWAgf/oYNf7vXflMAvLzZNnGkmCbYcfKnhkDAJPA18B1Ukgsj
67j3dVt+xWpu3MpO6t3O1eFtdMNtie46Vk7IwfH7FkIzc7SVgaTg3syOxtspie3N
payLWPsnpWZ2S/tu5mZ764Y7BzgmmL5yPL4+NLOHdEZqHYo/meaIMoiaDIWa4cnQ
VP0Skhp2yipl/arSm1KjulDlKqzUuOv56wN5fv5lfl10876jtbxEDGKHf/v/C7BV
CUXdr9ei7q6E8gGnzvuSxhZQ3oV4YUwhzPonKsYv1AcAwsgsJJwn7XczU5mZkFxu
T+1TgYZMBmF8GBAVgC8C/rvJ3jsWaqug4xau5/2VrdjdZKI0O+5yISwcRa933Ip0
TYyHcvZpNYB8pYjTJZwywlCJBjvyBwycG5VLh4ED5mt8dAuHtATJFTNADKJY3gz7
yssOp/evcMstqhAB1zKqz7VBvAf89eMA5L8t1xCLewN8DdGfCg1JblEAnb0H8NHG
MGFa40olCbjod0tZCVLA/VUlZDS1iXQ5bnkT5jiWUNCmdDK/3xUTqsV7r+uBv3Sa
1wgy8GaWn+neiM2u5/JzDLJ5o+lRvjcMMfnUzdc40ygVV+UCQMNVQPZA4h6beKA6
+ktgqUlW4Hc9tRNM35oRO27X8etnU6F/cQ1TrMICeDsLLGgFXNEYGl4y3gBPAuwT
jZErCXAr30DV6NimgDfGpVwh6AYCH1+Ax/LT9C2FggP6IofAGKQJVZlZzPb3ZLXo
h8MFx69hB3Ye2SIdK57gz3OBqA0qLef8Ss5eyFFoLM4amhG/BHhyZ0ppKbG2oAsC
CnSqvAisRaTEfqnupZuWmgATV1w6oLz9YR8HV5py0s4ali6EJm/3kNME2RPg/0FI
asRVo+8zPZImoNHqSKdPUx+Fglsod6EA5oNj9FJE5+maZ5D/JjHqPf8Dbcqj4Chh
PO1/UmsFWwB5HHB79l6LvCIpaCVP047vbO3Mo9qhS4GSpFW2npDYngn5ORRtlBY+
kECIlOIHuDLj6zkyl2xMg+Xur4Jrn5FWmDMtwr+yxxXfEMWXvwynqh8d1sQdywpB
mC6wTyw41Z5IF3o2pXz7CKIrkZVFuX44AM+Sr4ZKRterNnENPe5ycbJib5XQMOXd
XYxEy54GVyXy2mC9a0etoynSL4Z8/nu6m4lxLNeisiLMxiK1rsHmN5fNZ/2H2HbA
9i200wRt+OCJBGJRTI3zIIXuHu2xc29k45fs2JqH7i9jRey3nN2Y6WJ4RfkY50d7
8x+BHQgqUJ0bFw3Fh5qTa9qiOSz+iXnrWDLo0msSUrcsEPnZD+h5zQxcC3wgPZys
uL722hy5SvbRoU35Q9Mr1a/jMv6kYiyBOBiWYCsMgkUBX3Bqgmykw6ZFunhkoMPR
Qs5lqBY/bQVNBGy2Nbh6/g3nBqqjZxFIx2fpY+Xy2Crgv9L6i8CPUYzAwPxwc3ll
7JM4FU5948QJYlR+bzA/yAV4roT+mnd+GCFldvSuHvQzxpC8eWldAejg52JMYw+R
cSLwtpzAtfFB1MhEFqw1ZRavKgaI+6INGXQWYfOpEHYEbNx73eNsUE99ZbqGDMz7
zlr1xGJuL6GhjV3kQd/xPZBn9iyXDVyUNZn8HC4PocB4MIbNU/22Th7viJ8cHsoZ
iDTEM12zn35KdqrCp5TI9YYdyr1EILnOy3YX9V9gxlSCSLn4m/Kh17S1Zd0I6a9X
sai0ieqAnQmlupQFfGKgC/u07JFFE3IC1FNpHmRPALFwSmXzJjbr+v4iz9QveCcP
v0tJ0G51eJFVXx/vvqouzE+B6vrczT0t52GT0YS0k5BrCktc7iukLZ9rTY6U78Qf
Fsas4o0gn48E8Pm9/6/EnrwvrAJ1sMuDo3SDOm+qxR5aTgPd2TUUKOKW7jPtk9S8
5gCOlSeIpxMB39TgPZTiJ3hK0KeScnVZ40OVU0aKtCawPbqREJiKBQ5VfUNHxrUo
vgzoLtgokuCi27t0DSGTanAaLoCtTPPuwoPjCY5MQgsEXk1JO/epYI88Jh3KpTK9
DpwezZIlDZ26tOlHiJmDr9VHzVI69ejWl6Gpa1t+er6pq6qGZR7ZO7Vg2nZh/YhR
3PSZgl3rusBCtgf3A3MZ60KClkjEglKFVkUZ/YCm5aUF6+j0/BvS652LjCPylpDJ
6kmx64bHnikATkN/5PxLpUD3kLdfBIT80irsXuPcogeIJ1IrFFXD8iQKVpkEvUgg
5AiVSsBcExBLhmSGjQFQQMINDZa0sYTfF5kRJKzzPjD7lG+mvw4797rzkcQtsyCo
mBlJ5Bg6fh75El1Zlea90WqzGbHV40fjXEypUij2RtdMF7eWIf+eNgxelqhChBuu
+Qswj9M7HfsSJQxddwELHDngN2Q56rBeqwb4DCsoIWeIV9qYlGUnlv4MC+nCErcq
4OhtiBDA5H7vhX3cmIMxBOcI9SyIjc9nQRY5NPTBfzcHi6VLEgfYn37N4pLOQQ25
gxkT2EL9YhLLnlscI1WA9WGOpOX5h08qVd/Q+KsPbnD2h38TXuO9Na+eX8bpEiUh
ZVjLQNxRCrozAMWlRmLjRGLi262ifuKg3FRwbgD6NoyWA7WYyA1ptG8KdyJc0Tif
FiqW0osbB7Y/ywl7rhXP67pMNyx9QBES/3nn9B6MyELNE00gpFFKqOXiYP/EPFZX
9hOSIylDCijyvI1D8Y9K52Q3TZUvPrzbBKpiQH19FPwX8sf63FQiUhcFvFUdeobC
ammVN5m4UM6b+mQyYSCrS+h8qzwT6ZU3vNjIF3gxYm+7Xw6eqUIRWLxsLjS9dJdT
5KvfRn7f5Q19waoA0IG0RtiG2NJMm2mTyIxuwEHxyq14VNaZt29eKUYOw27t3Q29
tXtPg5rApHhlQ8GjcK5FBE104Cp0TLPNCoS/Fg+t6jZuWBb70L+LYJaFVxUhX3cH
iQdKhv/VKXDzuMGsvtm6q8QygF2Dkscgmbfyu4TWvXN7pXyh6UwJlX2gGei88lDd
rrTqNKtSzAln6xL6INLb3lcXwl/OdIOcQTs3TTUgOfHjcQENv14UyEz4oNozFMmY
09TfnMBitKWnwwfGTbhg8N/sDdnhH8e0EPA/klhqliEcnvr+xzjlBWLm9s83dNu0
xlhEBWv+5i1+ZqPpU2buOvxiBL/LfCvAMmejb1leABuFsG8Oa00+AWa1XksP+XPL
X1y6JP+hGxvgX4SZQ7xxalwr1f3vCWX8KsrznNf5zJYgOLzKD9S0fph+lgFB6peI
i3Vg/J4VMFjvK2hwrVaXKAtgAw7q+Nc7TLhpHbf96J2PMitz35fH6uYaNVVNyy67
VYnuqUmuxOz4gx7/ja1X+Dq954dn+WE05rwwSQT3b6Sykj/Q3lSB7ZTjwmDrfueu
C8UQJymWt9e1vA65sM2hzv+rwZIY3D94LTFX+JNtxk1L2MhfrfDX+S9Q5+vWm9YZ
vNDUzMno2aaFkEu87mmQrvjKb7aLNEqYpg6+5RwqbT9hfeX7wgieA8Cedl8fLdbS
D9htqV+y0VzFK16PPJMx91Pn8yG7lAU99ZVi3rX5cv9t1DSNdOyyvIlzizokOitS
oKSC7HH4F/vUJ+KIecn+EPkV+obDjacHaekxapqzzOik5xL+m8t+XcMggDNCaZqV
mmFJxkRTBQElC0fHP2fHcep6XT5CD1ZhTv+ecPiIqAgwM0j20n8rdN7PTbFkDey/
8zrX2wkejSqU88l5jrtrCp7Qmj/V9PdWDNq9o3ijO8aIPA118+gzqWPl5A/cNvYd
GEsq31urPZqt07rAjv7lSJBVmvy+zpd2yTiuWIZqJkE/eFsylz6c4ORZ3b24kEry
XuLgiCHDFI+lxp/Dpixuy26ck7TVSFf/57QA6H4DoLB5EHn1lpNhLuE8lNuhIGeD
DKcn4bH8EvaIY3c31YSmmvgdMPmiUUYYqU1p+CgOlgKJeTWqxAXjuNI+bhv8gAnh
C0ygCX2QDAnNT8PEeiOmemIm3vjVsALN+oaPcoR/UjXTrZsoYNAuo+HgqChtEtkB
5H5ULSvLu3KCZJpHedYKPVDo88Tym6dMMV+P+CMoiHBngeAXmEBpOFb1L5K0TgIT
kk0nSqB2niQAr4PIQcevwsgfUX8sOU+kLmh2xFF24v+9ltzn2CbVJWHDs86FGSO7
hSDtNv++rW+cQazZwNwH+BDNjCAKK7btMXWvRNIAtmGEicpucBZ+MMFHx4GLxa+N
ef/wZfxVVOvOrjiU+OoS/8CcRpZzMWNqPWP7tnYpQ7IOhvbkI2iJz0VpZJBej+Hn
AfSR/5vdq8nWLmwOmzJaVTpIZQmdH5JKdRImlv54gO7auoHIB/VPOMmOZd38LyX1
ekDZdpJBUArzd7TaMTlYN3WfJwSiArg0qoTuuBWIi9Mly2vYWvp/dk2WLGCqrmQ5
ptWuomGA8TIPaB9FkVEEwPnjcdWtHugceyNleB91t1cT1DmauTGImnQ5AeDy2F2O
pkQW4rf0uZO4Fe0fnceKu38dOEMxUUl5IoOTUR7l7j2ix8N0Z7KUBLpyhjOW/rir
b+aezVA6OS7LCbpsY+4wuRZXSctvY/8WHxcPf3ugjf0ZA+WIPxIK3OXCZZYCO5tH
WEkXrzhjYk+Ya+8m/u7TDUF/YAy9tha59JVXIT/rMRtAREjPN5PjxakrLitnp1C1
eRiko6TdJ/cf22FcNZBMAz2jiA9yWo4pmQMVUp/uTf1anmVdfyIF0qNk9uLM1hM0
Cm3zZZfQj3mJYvWIwJe/dB1N3/JBVo/44eM2itC9qfksjX+X8JcttQTjJPPdgkm+
UTFjoLKzSwMzd8pTIF+myok1WOUNsUOiKQheUyn8JDkov+yTXsJxLNIPS6luzFeB
zUqkzNgJfdErGqtpG8yRTtiYcZnvKStjuBVSQK3ymZ29wWeQdcg/07/miwWbXQaV
Pd3NmYtq/k2PhgnGMS8cGavzx1+fH1I5UqaMVYOmuSF84QdQkuarqT6G/O3dif93
xs2UcdbahHQdmO2bl0RWpwT5eMfxLLithbMMEsxoeXhYtEuDEP6/xL+XxYw5PSO7
Sf0I+IdZHbqgL19yWedC3qZbfPaMysMrwHxIeSO6P0jaYw7DnYxaKaFXMoi7gIRM
V1VJCK9pie/k2WCP5Q5B7d7SVrx8soTaDRbMebqdwmoCc5MGeurO1XHBeGjf6wTC
Xqr66rLJiHEBayaEnKL/ig67ugqMl1oJQRKjpduohsYnbZCg0f47WJIGo4bvctOi
DbH/cHT0fcG5kF5oFaE+GDYIcV/iI28JaMyhA06mOsg9Im91Uz6LD6e2zUkH3Yoj
z8x2jFuiZ3s4cY5yzD+Ftu5TbURvWWWzx2Rxy4Q2TM29CVDXh1URsz90TK3p8sZt
aAUIaGWEarpCXlsHUChpUHmiXscYX3+dWMiaByqjl/s9rQGSV7yDtTYNeFyoCxJP
Oq6FALCWfJNzkgUOyF2/KbqTSLpdKkc2BC6dJj4HA2tkRk1croGulh1C5Bn3QGPY
C7Cj53wCnPNN9ochmYbI8g0/T3RpZogIE5rucmhdteuX1UdrjvB7zwbogfwAhniz
tljZ1Vctz31IsqDA0AejZy0fICWYPIq4M3HGvS99HRMYRoHDuqAbrOKrMx+sxG+9
2VtnW2WP01JpGhPafX2/neqawuAmwg84YPfiWzZqZZlZuX1QJ4rnitpMybQ4g4YE
92vEmTl9VNTqDZh1neYvkrAwcGCySsaMRj64kl46EvuXnFEQtELU/GQRsSpvSUIl
4duK8Z7oN2tI3gV3Ei8w9jjpJ5GR3XR2DTyIA3uIbCU6YB7Y4esojPTmaD5EeCgB
8yxujSxKtk2p/JuXpuk7V4FD7E7K4VAGd0uT2WTO9jYJk2cinB27z4Yt7EdZT+5m
bYncZ2L0uJCELtYsAni/Hursi34nMCFUk7Chim3abuLq8Ey3KMydvj60t1jOb3zk
UbjfJWVHD/0ZMs1LR6EGprVHuZbSsG+JvOlLCpsh8pPINImMoqaLZux2KwLYEvpk
TpAcgJZ1BTxnHWt5QGm+sd/rrSOD904+vYvsllZNX4Rae706fM4KaEeE9yFuOEyV
lODF8IP9x77FSEU4T2gGmfYgXIsG+3ALwC01zFd40qUYUH1WKJPW0pjROd2ExKWh
EDAvWSYOjWCZT60AmkebTg7cuhLBIQYbGmOvvZRjjESXdsEuMBKLhTm2AB6TZ2wS
gRVuf6WNs5XOnVCU14qUskRE+wUNtgn8pBC3mWuwGiZ1zsa+5K59cDGvW7IIeora
a+LKg4k8zcAnwkzdAU40XG855l0g1brh37N7S16w/51UvithfFKPdz3S1EmzH7BX
d/I0JaXG/fsUkmVZWtVlS3kgrYunLU/5TOb7XqUV4gp19fosC35a+et1Rd/Ck/80
xnZ82O3XBAEiZKuM3cDBdjgg9Lt7E6FSfMEyeiQEzLXLIpsh/CNG3HL6E4ZIhm3e
N8CwkWcAnKKF0EfQHxNjANKFyoK3E7nTMMLf0f+sEim5deNTGpnkzwYG1jHp6q/h
Ff0lZu9uZqs/yOA8NTmeCxI0vWacubOdLTq4tcZhtrAZTqXYsrbmjnD1Gg8cOICO
mc2qqku0oyRePFpfCSzFGKx6O6lqfaxdDjsPd3ntv2uCKriR7n9TnOxICDNedbXq
8vBjrmLQk3RdCEGJ5zCU7m978rQ3p1Gud/MZo5pzRrvCo0XGkUnJtU+wjhpIPI0d
hLWtXjQQRt3zC7l+CtYuIXqpk4E1cis94mPQfjFNCuz7AzYn85bwRROa6+fRwTHQ
3IHAGffFAZzpqRs9vh+KgiyXewDcHx+mSvjYQmrgmSrIZNUiPLiUBeg1s8aiIp92
tyoWtWhyn7zH5Bvov7t1cypCPgHFCagJU6T+iqaCOXjI85ojgqEvNldrzWqQ3Kay
9tcbBzspZ6Rr+wXl3B9sY6KHVOPjtnxXmaOinIdvhtrV3gi6IfU60AAxBx/+rVKy
KzCkJxPmFYI2UeqhE8vdKwGDCzKeVzo1lRq5W7Aak+SMl0ChLmf2l4FE7jfRodzC
a5UUqXCpDZ+xzgp94i7PUkT0qxd2G9nfEr2N3ZjQFY1aEBbK1yYFyLTy5VrcgaXW
cmRYCrk2okys5nkSNikp1lQVeSqDN2ew8kR9P7uvBwSNZ/kvjk2cFJ9nj+Cnahs7
cSZkHMgZ8rSucbA0A8peS9rdoXM6N9gklfGWGHnC0YwZKskmskHX0cOwn9OnynFH
Nx84uLIClBOMfB5E4Lfsa8niPMmSRJWGqhS3P55Ofnkd1mdSCctAvdUcTG4CITpq
PXH07gVGrZfL9b63k8lHc6MLIheCbZfT5OlHI6wLaI4RYp2AWcp3gHES1X/DaYI7
ae9QXkKiNGRVZxFFoHc9kIEcXze6hGu7/elSapqN4PFgXk7i7Ze/7VjbQfzg7+c/
1Lv/cmnjETLbKYdykIl3oeP8AkynEMMhrdpZ5wCA1kAYVKt/q4h7A84LEV47jtFV
uyl2kQvR/DuCFnIppeZZTIHf5eHFi85ppD5DJmH3/9h2RxxsFYDw+xT5hgnYUt9u
DEeM9u1F3ejjrE0leFDv8un238afoabqJD5mZkRYBoYGv0jiBb1P6+lIPRCSxrqc
eyRHSsYKrRbEV6Rw0D71V/p3yYKw143jeyPotIldpqcYTrrRXtDwwdMtA5czBQy4
3m1AjpgmJGbX8fFCL37inPf9UihKIM+etWosrt8ZIVNsLGNIZ5Gz4F+9NzWFwt68
sd/M1rmJRQLmTy+wyZdlAzWuutyFcetOhdQfpr2Ehgb9vSo93CjdgZT8bjujK2xw
UIGXnhAmwjyN0SE0p7wS3kgSfuwa+AGqSTJ+9WX7J/p1DBpPQGe4oqmpWFSPXwX6
oZHddhv5g9JKN2J2zgmT4WsBBwqkKMvCkj+GaZ8oZj8Ae+aSrcUmIXkuCqBq7g06
t6kee8cRhWQZJ89Jy1i4xg+Oic/xUfoJy70kLyS16nxctxsZHv2XKgD6kv6rolS2
0qL8slgWC3a9OAKpLckzH/+RoA7hECkZOVq/Qd60hB+wiI3ZmXaNYJgUIR+mr8vj
vz4xAl3ZjFKd4/ZdpJ3jQ+20dAzi4yKpe75izLQFms1gzTV6BQrpXMMaQ/0BdwgS
VcISzs7k2iDoC1z7812L2SmV89gwtcqVqkh+gl9gYJQ2ubCICqu7hCmbidThmdwX
VoDtDeFpoN3SqiRQCSoid2R2ebiqj2Yl9+9qeU5Z90b/I1Acw5TEPxpM/r9NpVr2
4VCEintB+YkyTNMhOYfE9OmAMCU2Ib4hm9ZIhCzwAnuFDUHgvHx6MRiKIZVJTTph
AxpP7FWi1yZy9e6UUPIHKVzJwndU6l/zEFkWYTyQZ8RSnxB4AH6uZMfwHLbj2Ud4
EGb97YwHOs0/3jzUmPXENNmlRvRSzU0xr8fg/Ixc6UQnnlbYWR4p2dSPpuL4prke
8eRrjFpheoSQVDeHyqfm7QUbqL4TInJzyIMnrkrhVr4GOFhE8no5qC9ajIB/sqJa
EdBUixCO3JjN+faWC+c1kSKdv6wnpG/9nkqEgmgILJw=
`pragma protect end_protected
