// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aHQFNDR/XCARL7OqZ48bLX9ITgazF3D8cQuRYVDAzeWHvxIvmJUbYljC92k8dQB5
UuVtOnoxL/sVcX0IG+w7zCcUPPF5cn4WTcc3PFrcJQO/al/uSHJmL1eMlt0zWzBi
5de1MCJidYuuHqW7ToP1owj3iJZo3/Q24Y7BDa2wUXM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
jcoittljwPpToMmFaYIsbP5m1VbQwdbQ5ctZUTAibX9c1MF/8lQchrm/N5g+nlN1
xhdAEEu0DDSqQVMMG565vuU+OvNJPv3QpveYlSiwbD5P1cYU609D0IUR7PRUhWdJ
mhbko6W+aT3A4EujcRpwbxknZHXrRs/h3QDjaeR8Mnxgtgzpu1c19CoV+F+idSW6
RIOECE4hrKVBSspRe2qXChiWwv7pGE+3MM3OsdUc+dtq1qVJsQHfdO8f+EbZyccx
i6M2YaYzge8FOqjO1C37Rzhtx9Kapn6kWaE8W1VLNI3RUhJi5t21mkipB8sC3Ms2
ojRvSEWfs6jY6UU+AqX+biw46i7AXOztC4wgdwSKx9DSHpDp5lb/xmRU2R6y7HqF
CCwjQvfPyBEZNvBlVMYwoLfFQEKm5oLuZkaIbRwgs+cExl3sIQ1S68Bo/BXsu4W8
N5IPy5rRrrSieI6DckkjDo8dlJZ8qaRP7ubzhrE1tI0DsxC2UnqodjL3HWhSjQuw
JdZcsK7kOMbVcS2+u+gwJI01PogM5B9fbgS+AzLMUOoSt3HWJDjBoh3pNLk1kiMZ
oqDq8IN9/CT66fL8R4ZN7KEzexxQ9smTkkoOFBqqKsPPgLOJGlZeE9Q0iKsIiyDf
7Ah/51GnyBh1nie1ZWX3Dri5WXN+WpQLAssD9Dxso5lAImVE7jHb+TGn/Sm93qsv
IhGMPNWp5D33mGIZFHxYySbNMJdGUcxHFNVtjL1RTlVOWRiFUsBx0iC0AaFxp01W
NDQd3B9uL1J3byZGIqh1oOqBTIkx+V3WpbA3XcGjpEjiX7FHd/U1Kmz2Otodf1t+
UI3MX3CZLn7fRs24kXH1BmkqgH7wdJhTjxolJnQR7aURTiu88zezLNtYLL7CM39x
snmcnocEZgamyXDhtEb7BKKteuZwta68Ic5xfaN9CWS728+l42CNJkVu0AWdS+nL
G78tDwuPnw8W10pVNel+MT9xXAvAvZqNn5MJEuWEMNiFNMT2YlA+f6tGUprRoPHH
1u4dM+AUhB+MwUc5qgdIRpALncoLTBoGZcwske+y76+fNc9bOFS+NjZ5e2611wtx
ls487/IrwTVH+hTIJvxJrkrF419jFXbKpI0gf/a+bSWN+r4edVQdRgC4iNVHz8/8
xpKcdEKkKjrsCdiylJYa7+bANe7g6BapBV/mHdyJwRtQ8ij1jabVQKETK9kmzLcB
/b8o2k0uVaCsUZPtMwQ3PfIRgrx0iAv+8VNbj++VTaQ0N+MDaw6yuLJEKNsStR+O
6z1rWsUjsXZyev3eMMxSsqrq/z44sj0cv6QEkEDuLBZ52MmXxcEaImon1WoL+nGH
6wuMUjp0xlCVBV8Q4YGFxq4Bz+Nvd39Bt0vcxghiylh6Gfyev+LPCvPadU01tMt0
y9jiJWedETVOubwrZMvuT4T2FrVassiVqcZ6p8LTepC/LChelqYphrAgCkSaLf1P
D+wwkXqgtYDS/fu2pg0ZEwUtQODIOsnwVyfQeTLfh7+19woSTn8FqhlglXIOrp2A
YmxrxAhORMTFfRHz5OW2VMcwMMuWGPVlNCGhaCyM5AXDAyVvGugdvS/n6aj+AiOK
CnzjSUs5CUBCqtIKR5GLZZYyURqWOb5Zs5GqBFNR/7NUuMkrp4XhDDmysDFMMtaO
U5UJYw0t3YmDsGHXYT3mg5jTyeXugznjWilFyfD39QbDhvs99lA0YinEeIzXwkR2
nZ70lvGokozlJc2lZ8DKwJaeTy/Y471V5tys8LW3aLGp0wJPS+KPg9TBNNu0FK67
KDVkBJmEjiE6fl5swPFKnv4rB/68OYP5uEedYioFGWTKyqaCM97S3nHG3eSAr3Cd
EJrnkTow4Xb5kYvsy0mtsafNt+bicJjYMlPx05ThDV5KjZaeQRDR00OfLyXCtl4i
HHruzN1ZhbPjDw67Wvj8yQj+wHxfOTdGejpegp9E87oizpt3f2I25DgIis3xAFLS
CZ4IA6zNOZM2+9LbGhP2tUueaI/7JDNFtUlREr2ZO6A5n96ZP6z5IfkNkcaKk/yQ
nqlEvqzNIuPQGSIQVjXjbpjsYFLXKsaAdoDej8YenoupTZp+Gv0xbMNdxpVMq449
8DqSClwmqj0xHT4KUZy1dB/KIzDnp1GUsvSUtyFu6RadvlD7Tz505F2NyYm57YNR
qJ9WjKEcDliQqXN45iygKCODXR0ey7yjHS3Mtd5AFRu+w9Xz9ZPeEK6/6KI8F4z8
sFNUEGqb6PYbs7q6h5gi8x0uRkWTFA0jbRL/uf1N8BkRJCkXOA2W6fdNS7Dno4eP
643AUFvLXUd0RIAuiwQ51eSACf5++3XzRfjzXHP6H7aXyiZsjwieVBCppGODORbI
TzVNk5C3/Ku3BQzcvXIkjsoDpJHJjNo6xXeLV8YzDQIMyJFJUvC3jXg2sJ0eFwDU
BhT4p/L+xtcTysY2XdULKQxEehQiUjmaa+dkYg9XvnZ+T4k9tO59C5sgzBzJvTLI
s4HGsEO0ESC1hlb5r4xVIjdT3be6F7DInjSQm3HEN74q+z7WWA2XkMkhNOeuuBYJ
tLjvoTko6tFWPZoGVhZ6HU6yooU2m8IY5mZBi7FlATpEUEHs+svjqwfnXlmLHdBg
x+Ttbq0T+CwnBiF9KERVoUS2jlTmdSK2IbLytb/FEdPlfxketppKyXdg9lR/FkgF
1plRPVIm6ibbGcY4PhoxKIEnFt04O5XZSMHJGbIlcTBtiiVtDqTo+mLZ0iG+GXy+
eCbGTO2rHlkjIGr4FHdESRmlNi0bH2phFhG8HtZ36pI8KmXNfWv0PzYlllpvvMVh
5uXIuFHDNzxzue5GPNiEDTySv+sstjCFyi4ebyWG6ZvY4LU0FkSYu+4df6fzwCYt
MtTJ/lNDEdPHRH7af/PkFc4jYDt1DCLA+WRmczgpz2Yrld0C1tcV4QURFp+vX4WG
Uc230l42Sq7DbH80fvIM3XofVS4K9FqRNnjGoPny6qnTohXJvT4Lj97Ku6UDtXbh
0fSAKi85h84lxUEpVnQ5Ixcym5Y0DvpfxC7RnH3BiGXxsIdbgpUytAD5VZvH76yz
z6hieMwPhp3nDgSRtuQ/EqsFYQW5dmIzZZ0y1JF4ZLIbxqoZs2kqpH4sA+hpGDIf
WSAvO5KyuLvPUD8Ag00+omsE+WnXuJD3oMstsM3X/d0wXXt+6LzD+IeyZn4JDRbe
MpdLQPkp4BeP21SfHcdIWmWjQt75tb+I4PG/QRI/JaUNBBfTSz8tciJAh5lJpCpc
bYHAjA6AJaUCccwKNyf66cMndGUCM8FxHsGz1sXeOwcYcKvXtbjl9pGVGM/tVtQ8
cAuRh2EHl0g77BTeVwUo/FAH5RE96KwHWL9KEgyXROrLtsOUKfGExZrrcWhs2D40
+s/wUQwlZ5MVqcps1tCON0SiN1lhA6lEFaxY+d8+J6xvUeuiRaLbJAcAmXOxZ4i8
XizVUDUIzXjXcghcRkOHbpLYBgLb9TTdJgPC3uZ6J3K83sVOmZrJLpiYI5WEtHH9
LtRBxlJwcNOmxFUjawP5/r4dwaIbv7Yaad1ZdxhP8u0wEsCEZQTRd05FlFJHLTCE
7EQrMWuiFCo1YgvR9IjjyAWzJImJ8NZsJaZm4WaYIiw+FmQD2wCjs8gj5/EcCg+x
gxhDT3VEs1CWmByDIO/ikbi1diEyBG0rkXiCD5hKZPeWc2dkV5RJTH79y1rJjVy6
UWXRuBwvx2kGygO6jiRFlH4FCSRKlKxI55JDtOgXexpHUxqivJ5qM0dZqaBRPMlH
YU/qqDX1FhNQFRngOkMVph+0PubufCA294B9gDAxXXUQlPlowLsb18pSOoG8NNsr
JbT7sftSbekbLau1Ii1pkfM1KW/b7TrRfzonQB92nBVpKj0QGNy3LJ7zTaom0+FZ
YJefpsAzUmQ3sj/L9MffJhV00ktQfn2F2Mz90bPaWFB8OZpFsrlYh2GmiSFYR8O0
/zLqLMkVJDbqGaSzahAExwg7DJvwuaP0hgAJMPy8bz/aWaA/4aYtpYB5t9xlFUYd
QlffWfMpieC9sCqzgBRv4ZhNqbwHseg2BeBJSf1lsMrFs4xO/B/lcYikfOMOl4V+
s5aVy3fj1GqtPmYGNvoWsR4tyq8PADKs2waEN/aVdHhWSvWUZr3N/Ahb7cvQM+/a
B4/eZkNBCXpNqbSU5LdCRYDsQR5FK1cNc12r+vGmUvNNxqcJkjRTS3I9aeD3+E8b
cUuV+ci47/KNEBUdpByn87rsOsPNKMqa0LbCiAKiGImeTj8dlv8Efik9mB7xYdjq
B6y/CsUAqkBskET/8rfNXzStHHHkyL3SYNei//BNK9yDm90kmkpDaK1KqVXqePMw
bniuDk9ihAfiuyx+cH2Le24VVVDF4C1dzR4Ax2EVXFkhCIlUG9/ZOM5EqBTVgaxI
2dVhBYeB2Y+Mx/UF6s96DpH9OtxZvuhjmIdqILr0PZX//vBX1KihP1JcKQh7kD08
pFqZPccl1HBb+jm7vTzDZYYv28x5xBGZLCUiXq2cvaAgfDGzrfsYG6uye4nA6tLl
5CbUKFpW7bOQu4i8rU0khS+0oVwNzRaZj59K2Krz4CgfBSp3IQoMxHjZpptVtwRI
ClXXavLfucJsayVE1SsHhvCpwSSyJjD6jzmc2/MQNwKqTIeUT8US1M9rOJnVoeIc
NYE1j44Onr36r2KlmU8jPovvDnktHEZh+/nETHSV1kBCSbEej8DJjBd0nnc02HrB
lYJTtz8yNnFzM+y/EL7Bu8BCY3oRiO1E3aXdpk7MZ0tnEyT+zmKblWMYjRUohOmX
UBvDqLYFaPhKGpJvJOBtSsHAcOp2tKVh0oVKJ8dDwuMC4LMnmdcSsUM+nnsb9dBH
BCi/ziC6Tu7AGSOnv6oTYrYa+1v7wO/qCZAyt6/robshL9frzSNTtrqd4smCc4/E
4TxocUxvxHLVESk3YX0iNLkfbeL2ZzoppVtoy3L3rSb3vZine3Cevlu4VptOA/ti
0D6ToRfQvr5L9ClUANFTeH93aK9nL1vz4cfIm5f+zAvekcd2ph69xmQa3usikPq1
JMTxnxF/nd15LL0dkJoQzEmeC/nNii9Mw+joB6Up7dwDoJ52ODlvq+UN8yk59jCF
qDp1o70XB5MpixR0zf2P267d9xIg9FBNpyJfe+DEhMVp2yY1csQBAgarr+1U722J
p85zuXgScVReCGdulcNpkD8gR8GxUx16rGRiHCeB6IT6quKGowI+KJByqlHcSjol
g4uzEaeRvnXswiL6GEUyGX0oEVsDvGxk9sjLkW/MNmg/UeoAIcFc+nS/4sUGArVz
8a/fy9ReartPfRPpiaMA4vnLgybw3eDAG6TFqe6XJYZpc6UAeL5u0SiTdBIGvh5B
QjX6R+Uiyak8JalIH2Jxu96N9F6U6eZyAcx1n7KUzaY6MGEUTEneV2qPRDMVYO47
iuKyXyNvpZe7QwNjeLhgTyt8wv/0/t+OtbCz484iGJ6jSd0/VGhYdIdAXFXgN2lm
bwKmcWl2ZrNB+KDxnxUHm+TiHgENpIIsNJbs0T8v0FSnoZH6sCTo+Z9NumaofU5z
Bg18suWM4hbzcKQD0oQXIZ/gQ/UE+/V5ic5ArL4tZlXjg9dWVWwZ02kLEIQhN5P2
KGI4gZl5/Cbm6rSe4WEpr98l53QPORsljX7K3qRKoRGdDQ5DK/Zrfs32WDOrfdzj
Sct1uMI9aVO85tnqa8GaHuvTJvaqPlYpIQ32v3rycOHQf6gYXv05eE2BgNibLB6X
YzndQL61x7P0SksMO+8gXc9FBtN9pU+Y3OARLA99W+i1nCH4GtnN61cPJemJud1a
FHFObrqsNPp7DUSqaywOPdeEuxnomjlRH4y/NWxexxmAN7G/oxgAEUjoOzAtCFvd
J7c/hFIqXf8Pzd98wP5u23oTY6n7oPmvI2KvsjS8hrSWZqaqMnAcUourwqqXmYDh
s616m4bP2U3xdUxeKsJ0GnhaQf3M6SFim4EC3oaCxG0CTt+1VaSxbwPun8WZasX4
KiYPR5bp9kekNZRVng+Y1IxZDTDIyzoyDRxq+iWlhcGxN+4xRyg/vf5EJ36SLBXT
c2kKi6vHtI9LVmMWE/NjpugM8upMJSgenJodGCvsj6yxQt4Lx0PZNtSC3xivC46Y
ONXJUB7pwXL8ZQbEIES97LusmhfusU0c0becvx/rdxYlUrefSGNKKwprwx1aA3Oh
UuTdcOxiRVjJC15uTeHGhjVcY0WRTlpnyEjwjiMLo8bUjuz1LtLqC80J1uIJPAJV
+JzGi57kcEhKUHrMwoOrSEPJtx84eSWjTkq3g9A/YxFSFtfTfJz33q/X7+oPxDHp
sa/F+P8i7SSxrTZfXNEGUz7IFPn4FaqPkBYGs+ovyNEmiZgx3PgM9+cAw2+Gxdiq
otmHxWgtPp7Y1wOYk1wfKE5+FeQT0xNvRTHsoxzdB3gLxy3+Yj4ZmArXpmJEzd/Z
UvndueiFQ22+NoypzjYG2ErhSinwoxumpjExkB6ZmqJs8NHSwIX+5kL829ovUtT+
mZ10a4iMyeGLXwnxycp+G/v7G71y+R7O1wWBB+AOutE+TC7QOJ8zDDmOsrI/M1DK
xDf1di38RtRdd7vjTrm9TUS9zFc8JMmTUA14Yzu4HtOZUPKxIeBTZqYrLtH0pidH
lO+UGRlF3UrJeZLZiMlDwyQYCG3S7Qc906UclLXSq/UBa368lDMK+7k9wokKzSeG
jkC2n6yo7Nd9C4+I6Yz2MenGMIgv1DbF0kgyOJ0AQarUTEEaC1q9cflbpTjVlCi7
9I4927wd3P02kYAP9Fw0qvpqk1H9mTv9iIJ7X61WKymkkvtVR31TBur6JrUE92M6
xgphhMVfGxGPZlCASoY5gXqWWiEBTW/3Q0gpfQ7ZygwHecxkOprKeuQ+VAKsRsfY
YNft9lLJqV6ELxHWuC0xotxX/wF5g+ORDw6/q/sjNwG9k7Do5Aj4TmZsawgUpGpE
oKE7KwXXtvAFeUZ4ZR4GuI/vi2UvonSsO+QsSW1QuExEDZDeC2XABBABW31+YMU8
FK3/PmAUHD3NBFjxiAgvAObcMQKrSLYk8ybzej2W65WXnfaCjpOnISybKBEIyZJp
2Pr+dLgy6428bJtYdIJ9MOX3RN7h4Ue3HpFSmKkN+cEUQgbc0jvNwK9UP2Hepp01
hV6OpE/wYCzyhHpD0VOx09p36wYII0JxbcJnAdZ6BL+beZD0+SeaUxPHAfsjEqp7
XLWZOawwoGofKAyxlmpUhQ8hU4477fK3zBNAuGB3U3ldwGDYcw5ogCyVq9DM/svB
eJODvRxvfGLx2gN3n+q6u7yUgIP1RuDQBC2Pn9EYiosBhp6VJlWJTbjlR3OS5/CJ
8h87op/6lVitpZ9aWVGBooY+KBYbKnbOapiu6t5jKkuBRvJX66d94LBjcM4VtdOk
ClbKCrZuGKSlH3wEY++h5OU8apoIpMVb2GPybezbXpMGSWkYrHFy1ZvQifEfVmRc
bcX7QQXRY4sBnuTI1ka8grM1zMvVOjUVV/3hP80GUcgHtAomrIfq60MPtceuv9jg
jYgaec+SBvcnGZQ74aXIzTXECBKuz9basvKvSZXczz9Ae/yWR281QBUfaOzYIt1G
W7k4cuX5eY6kfNmQ7eoRpQ2/bgsGv+5tUBUBJC2Op0zlIfPs6MUOfNqPMZlLaCap
ipTTLSwf6Vv+cq1XfdqUlvRh1NmeUT1ywdRfjfyASkoquM8P2+Z+luFHOeXoOh2U
v7feM12JKSic2V8AJWdy9yNjZMOj6nR61Zx3FK76dx5uL1Yvyu3IiTW4pyT8lkNt
SZ1vBpKzbMfRPPQ0c/qP69aTnKSrwhhTujiUeh6Yc8AysMvQoXgiwjrxJCZF8+64
fIyok1mNu3MktFrvezTxSdqLd/UyjWnqk7GEOfVRPOkrvPbwk7fck4TeGmYsbdyq
4d4Da6bpayh6j4liQLy63M4LgIzt7mERJhgquQwi0t8hk7HNGzPETZLFyY88JjLD
PzL1YE6r0/D+n72oXVyWugHrt+5EsdMAkaM9OYH865zIIocOZTylBhJDerKwvvTh
2y/sxdXwyW8fEO1CpG0YK11FA4udaiug8cUJf6AhJhVTfZcyzjRuNMjckzcVcU8k
QENVWPXXPqJQ41ih53n0uO3lQ9an2mcwhP6alNrxbypCec3YaYOG2RrI7y01T8RT
4B1t3Hbswt5X2QhPvbgL3LTN+gysS5XJSauDYd/n3VVJ3TRC04uGDbpFxdRHfcoe
bd6Ki7s/PN10CiqI/zV/nrU61z64eufFHaGVh4H0cobj5QiQ7+MW0iAT/uKViZhE
V/glvIG982nJLm2iZSAHUoqVR16SoRaO0gNG2GojxFXn4pugwkj5b8/B0badmE3w
dzBBWqbt9/LNKs2+c2CMiDAT0lPPHN4jcqKR/28DS0Sj9IX0ygBMqGHGY8lducem
NpWNxhODKO1WZNbWV6bT8SCyOZj7i3Nlu0XXfoYJQBIGGYAiC4WBeoibcHJUzDrv
yAH2ExgH3zpFr9ekI5mi6jCnrP0B6glQpln7LYdUKS/aXa8F4h6LzcgMGT0xYKLa
CIwou6LSG6dZaC1Rz1ns7l7BO7cSaGAHC/7IvNBW/fX6NedOj3N7sIGWSxIefeES
7E/0PMY6z+mLzKX+ZHU2MvHa9HY+g39pFhAvFtuAsH7nwhWnAyqEOuiI4kHqZLHt
yKLOSwy6uE3Jidho6hwzNPmS0JRNLM8sjzi285KfPQJ0Kff/sCYvyElOsgO/P5Kc
XPCb6Is4oVmvv+tT+EDPlbsfGltZnIczI8+XPErRVjdHOifWDg8kvWb0wAyY+KTl
6OZMb37v8P94nQunN2mBE2HoytLGTg/m0kFMtFS453V5Vj1nRnFVzVynL8Zh/cLF
vBckFrGkZCLCdKNy0JkWqdINuhBySCNfGphK/nYsvihjviUM6FNqKY0uQI+jRgwN
V5MzGr99CF/eeIrqDVxF3IVSoiyZDX2I1huXAmvX+xsfNEPUHkWLR63Rn2Wnf0nX
uyKhCgDYXGTvr31yq97aXGZIuqrfIFOg+s9Um6hdpq8Z23o+wpeqJFXzboVRNDln
VIkWhVfVRCiigsCRQj/Hbg1fl2Kd/W4s587UukWeFlfhsHKj/KPTI9jH7EMpioLt
1FmvbOdMfdwK+N/y59ZeVIqDzq9VjGUP3tHgcJ29BO3dbw5fMTm2yRH6ccnWJKrQ
/AXHsm0gNyMk4pCB0l9IYQe6piQc/YFdG50ylWRwd1XW9GZq/i58XaHssOv6xikd
wjLsM4xoyPZXV8oB/u2ta1IqZcbr4mLBtRcCLCh+x/+tQ5d6XBmyYiHlS3w3w0ec
ErC9REOS1ezHT9d2HUrujRTNigIKEYw9nYJ4ZdChV0kNKqmwdBSHO8N7/7ufO0NX
fnv7I1Mi/4iEuBTgV2LSiYu9yOzmAWUfJH5jRnXEbJTWluEiCLdsOALJfxNoTiZ9
8Z69dKTW7UPBVTg+fVCoPRp2awl0Sx7b8I/nEvd6TSKeK6TRMqVZmzqGbiTYAEI5
D7oqRLjLw1DuEa+L9AE8WCM9bY3aR99prS20w7dLxM+Beo+tZiFV0scurOCtlHl4
58TQdfzRUv9oH+LU5MTE5id6xiruGk/hPCGPxhLhjG3wzFGIOJETnSLDLyetusX7
BeUP1aixZJ2t5AmsiTJQC8/9b1bIhJyX96IxNW4w8MTIPGEm39TWthF/dsDbLPzZ
kzFELsnY98dISokzhmkCLbLO6vOCJnMVq4N5kB78UJg0+briwjrzizR84/MS/lcA
p9IWJT3sQnQ4X3qon+F/O4OQQilkBqYMC7i23BbxMdPy6wgl9jkhBaN1+2fKRj2L
5IpjkdWCQsrSap+4U9b3lyTkkQTTBS3JMILQtc1akFtbYJx9TdtoYf+ea7E6rvme
FqFDLaRFfHDxkvpLnRBo57BSNSl9ij1ZBd6plM6nQSbRsjCLxJd1NxbohkcdSQll
n9u+JgXntGZl4rRWJC6uWdzeLf14FpTMTtJYOkGlPkzTBIeld/LY/sJNsSeT99Km
ahvrOxOuw2tQOKtCVIb4GqEWX9lDJ6K+ueJky45TBj+ZJX21HbjmGs9Dv30KyXy1
Ca+VH6sfMM6dV//nSvsoGhAmqpppC9+wtxqbVg8xa6zILnEo1rhOwtaSLdVCvKgu
PeNLwJB+cPVLg/0vNIB56SYdLEIIFpEaR+MsXOJ2jeLzf+4T4LrgKI52BhZLojqB
Fplh/AbIGAic0Y++vbDjLcM1EecMkygbghRlaVKMBJl5Uwy9xOUfbwd7lVj/a6HN
BJL9CUO/Le302j0GGclTBNJk7TZ/wrDx5g8qt0cu7sr3sZ/2VH98enta/mIvI4+t
KLZTBqJcgly96wabkMiagiFTCdJ2UfUZMxCysHtQmmxGvp4siSKy6RReeyy+EOdQ
wA0MfNmDEPZAkxUWfWXxl31RL+2AqX4EhjeZoFSRSCMJ0EQyHjEDgCDV4BvCn3lK
tpuG9nV0s7DAmYRomItmys6AXHN/DVJUy7a/TNxo2w9DwOIly36uP/BAnt/em7iI
sdSyK+LrzeSmdUxIqTHxIOSe05dR6W2yt6znUR8bnA+yK0U0qP2how/M/lSfvFty
4J1ppEZbCXlRls1OoyZvKXpgYezp64d4E4bRh3/xtq3LBBUx+Eyca+aMz3QwtGNk
JvzOjkxPaqTo7ucaCG7gws2XZwNL9SPJClznUq/RUKsUj3+ZnJ1QG6ftbtdgZENa
zI2vXD2aIhDVJf1lJ86fY6lznz9cdwwScr9ODcCg6Z3mKfZG+OVj1hsdpNSU+VG7
nHl1A1BhUle+WuA9bNQ8LTqXXSC+rvv3kRrazz7FCRZNYeN3YFXz2UgZeWcha7VE
HLwNuz5+NqBQ5fFGPH6OfpbTwM6gEV2YFye37zmtwIGtgXFKXbOYy03M8hK/PF4q
Lfj/J+33gFZNjUB7ltCOESy1a27oXmqaTtemDRnZtCpN1N9loSSB7KnPVTuLEy6j
N2GNMqp5ydiohDTpjJlZju61FpwLJJS1RwRQEeOsp0lqWHy9L0ftm4prWCT7+MzQ
AmWckwVc0YGNA9gYv1ctFhvv6yYhCIS7+OIFWdqVOvMivLzFqjEItVVxQH2Yay91
seAtcDCLLtbHSjnIYrTMJFKqTMebgjQ2i3sK283fxJxS2RDh1ATxdm0uYUq4pjhf
lMzwHygNyyvb5uhAJXLMwk84GYoJQF8vw/+vPUsn+iYVGKYWbL44BoXYAkBgaz0Q
QnGPGovp+LXdg6HmHVRsPCkKAZ9RergmkIwhCMmrZ6Xlard2Bq9/azfA77HKRqNj
1BDk7kBPNcReXWrofMwVmnQU54w1eM5DLbdYSr7ncd443VhPdEe6UrOW/dbLkK7n
7+4sALldhqSX2ND+64YCtZ5IHtqmoMyfLr+OVl9G9WEREdA3Lwn+J1m8rzdboDF8
50LxCyhWaB09uE3fRL+7IsW62lbxb+bCkmzU2crC3+cm4MaB1ik0riLrAY7wy15+
YHkLHI83OrMk/VuRxKV7tx7QOZyc6k/3wr8mXq4gWyOTl4PynEmxMcSl1tTO8CpX
4/LzOnPk2NMsBuRsZD8yd7/1ClAJFNuhgOH2A2p752ksalmriMfLArgFoqND/sHw
ICyobycldGTVD/tDIv9gYtr0CNgPD46+IygS3+6/A90CmGN2UrKQXYpoHNGX1Vww
9KSwHysK5z15GulooXfpKyDVEqM2tOGWA7Lbhi4HEMFRAfhssPt1Q4ddVo8folky
WkZM2drvOsYbj04Vv+zSh9/SWubMM/ecu6gIQeDK7fymws/NmmI82xkJgpQMcee+
OKy4E9Og0i8Yvlcaqtgzx8/nXlWRqjzTPzuoVidry/zlv9Bb6z9VNoxhwmHcjpSD
5cJhShbH1tQCKLR7MKlK0uGTGZ6oupm72cEAW3VolFdVaoV0EEfRoEQz6vYFpWmG
rQ7qJAuP0w5mILEiRC87MOwnb04a4D/vQ2Bi7cRu062C6ysTzeRQII5iUftgPqh6
YXeIYPrSBqsK6i55pTQidM6xnei+01NV8MwsMrPpO/W9B0NRsvIAJq2oOQqVLVWj
HVcTn6FEiyLATAOTUEmANn2nu7cx/yLwry76uLGWBwjUnIuZe7H8O7s1EeFikgQ4
DvFY8RoHYVF3g8MqFJb25wZGOHDht+8vtQVRp4y4WHkixrhJ5NqlI7q0BJBzq4rj
l6k2yfUeUb1FjFRL57GxShvtuxskMjQOlidFk2heOhZWgiYosx32fLUxs8TIx30o
Jz3da2o1t/Z4VFXgQhr4Y4fkPb3jkW5YLYESIZ8/ZQ9JZwa8vacu3Dhr6nMHVL0L
1vnGiWCTIT99Ycp+RJ64WBjVTn2NJLeFOiGBTeNdg5jifL0wKp7BazCb4w2EB6yX
KnmvilDnthI7V0DW+5MzHUx7smXWCF8zt5Rl5kwGHiZNkQmYUT1x4OQzKwN333DO
967BSQy8zyN/Tl+uini6GMBpbdJTs+arvwFv6tCWFe+vIFJ71al8Ue39d5lpXFNu
ITvo1sXaK4/Plh3n/r4BVfMEJrwao4CTptZqik8fxIcJlTb0nYjGbPwzZHUp0DmF
6Vqh7W1LD1GyCqKkVvG5Et4/wwQ5s61KXpV3aRGsrimWeivWA2UMzUuI5xEgH6gR
La98qVYfVPV3v/YnFmRx35NRzgKep4zO2u74zJqZdJR13g2b4jwGd7aUwLLV7edF
gZPCMcddCku0tMuv9Aq/ltYvbUpMgvb9WLGtvVesghBqQj34tAkERvF4tz1RhikV
7kixlri2shEqMj6+fqQoIf61cudlxR925WvWLxdZt2J6zTqbE9bAG7Nd42jRwyzS
J5Z6hydxZWKrcI6/81i/LOo5vIfYZKxjGxMJuW0M231vgk+1sZGSn6IXZ8XwhVkF
f5yFzFkel6aRRMhUVOXMWt1IElu2nw1hx59KRSNgipN990noKckHMKxqp3a34l6S
2dtQag+xtBJVTWWi+OaMh2YQQZmdtHd23ibybH4kdcwc3N7PiKkgFYK66sN7sH44
UHRueW9apGF95okkex1YPAevHSU+k0p4QFzqUgAx3vgep+gg3anfmWjU6w7rxYl7
uzeC1glCze6I6GziEQ5iKG9stkOA1UDX68UPCWIz5Y+ITz1InJZX553AK1nx9cTf
Sslig5F8lVUQsvhZDKwSF75w/wU+ZJ1BcTqe1wzdVs5v5Fj4ybtfEJH7hnTg6RXW
euws+AkhcpGYSHbh2qXBLQ8Z6vUgPeQygz7PNj03/Uyt0CyViNiDQ6ROXTpE4IkL
byu10ccHqJ6422eJayBO6wwqIfE1XSAegFXvQPohVjKqpzwr2qzpjyfUOQhgGqQ2
56/u+KmWLFQk2Sx+XntCo9HF1TpaLgjG9Sa3WtJjhZ4jGDL8JAfJXiwYUy9gkTjL
9dI64ula/1mhjfJAYRnK2RXLn4krxX63Sl81ACXG8bwl7mYTv4krZm+imlNSmNdn
I42HUdmYe3LzAMh4layI5VrWjli/r202eC1pgDthSr9gR0GKGcYIm8cMIj6zpkPt
Uj/8IUteNDNIU+QI+EgKn+79xPyycoM0oLDRX0WvIx9oOHq7gTOq/Pf7Quj0f7S2
IG7wD5odYe619EFyOUdM2W6HFhxXyqF4gP8HcxLlWVN+9m4J5BuN6udJbg3wbLtW
QJXf6vvqFhqxWWdZ/n7rWpb+rMp50HBR41NyHcAyGh2IeGFw9FKvzwRHMiezESUN
983oRkUFmsTqQxLG+fjNuaBz63ZQFUmIsPb9mAzG8vtZyloU+eMBEOEKU5aIEM3/
lH+R8cRGXQavMcP6DruFqs13sZEJ+lLp4NPkJ7rhXaJRuHaN4np3QfBXqYLCwTHf
uKtyA3MQ+Q8zXq41nZImj+vmeavdKOnv941gPtIdK9j1C+yO7zIlqG0hUo1q7fLG
MGs7NJMRRU8rgeCfvqC8scgIRAzXXMnhcamKGndKX74uDfftuG9zh6CM1XSWgZst
wQ6M11T5mhG+qLMWWbcrWshzVzZaC7LjU4vBe61luJPeNvIs96cDhEE74JpZWvme
LkTa863lrbSx+bZe/kYstwdSlRodTKZrMHZ2Pvc9gzeVT7mt+ZruLCf8+/Sr3bBn
jVy1g2IU3RHX1NkdaTu6IQ37oL0IU0l2OHcxx6AlXhNNmv7b8NRjX9PaCZIpX5W/
nRFZYFlSfj5S01UJ9NeIMdXXB3BuO4fTRNVUBvBddQUIoBTvzzubrdzF7hyAE2gv
Q04XRKjZo2jqhUcAF3UJF1VegLegEDOVsr/+p/2aL9RS8uKoNVdfhJt9aGwLhIWw
lWv3SX19uJlkg7coOUbTQ7YJ1TCoJM9HdpcNLEu8ApjYqzsDC1KMgmxpQZmVMqxm
uZjwwVkMTYk8Mr1QZstBfrgp0fAJSyIMsIwl71esTxDG3BUuDD5il9SNbKMfXzbL
8MlmzaREYhTvSlCIdFdBkKt7YcUP6lFPcxlc4nLm3LSax37EmGu4Mtpy1/4xxoQL
A4+DseJSEn1CTJh2Rg/iqDGnBfKCaFDf+YRePxwcOo0AAbmvulzLe2oaRZoJoGpQ
lwG/REjYof/jG2GQdQQfqjY76XZePfR+ysw01xSzxl/38cRVbfProdn+ZOrhj+lQ
Wv7MCTLN0YWrJutpf/XGXCK6FYq1bD0jF7kPqkSndcJcDGnqqbiVjMzdCJSNOJh3
PC09nuFzfx+B+qAJJ+GiBkVCstgMf9RXSJ3n3U258/xGr1tA77lrA+NcapvdTeo1
YYufZxfl4YtSkKT7iATDsRgMQa2/XqQ5z31f6k2BwpMDcX6mY0IndLhmur5UhvSm
a3gDuPEB29GLBEUy6q79V4kc1H2G3ejE0w7hhuSXuvG3H9tIuUhAEkcZhdpIODLN
Tie2E/61Mhb3uDcBZibXaJ/LxwZC1iHwhpsUcqXdgQUsEa5rR2jl1EHraa33yIGf
IuchxQhmsTXNbIszgOlgpJExdTBFYQqcgAK7JktmPlfPTei7sANWgy4kOgcwbecQ
KIPYfwWt8UnKKKbr1gzV7eeqrdD0g89Ktz7SDFubjMAn4xMzTV8UkKLFBagnAODL
IJ8sBj+0McUFQBDICsSupUKVdIeI30Grm9XyjjUD1L2rydHna2pPmAW/CW+3SR97
dy9JYXxbzTo9PZ33582vRnQtEye9mjzUvOUonXfSZMcDq+kXRtMy9qcC4CfUSGN4
YSUtAYHrIhxDFVl9LBTOj2/tgQMdY0XsZ0vhl0V7uWJ8N5tKpAQ9ZgQasRP3p36m
ndxULc34aEz9Kc1Vb/RJMWIAw5SW9LtJGKX3q5BdOCZsLLEkY6al2vbnHQOZSQc/
Ziky4Lj+G2bLw3reQUnv58S/vOd+nYy+2J3CkoiwTmjddKGRTRVAiUzVqV04sVxy
YiC1OGRn2BoeJ6VKdoUPy9PnNNRy1lzXIRfYqF1yVA0LWvxclgFH4JVMVdh9llfh
+2keRUgCyJrDxGH6d0nrxSaAa80l+C1qhJKTHt8lnYWcy1LUCMpq69p95oDFHPuM
xSYcUuZGEQnXhDYytsMSm6kkPQip0lsTOaE44hpQKItZaiNxpaCEYtviB6GPCfHO
iqxQ5M/RhGOBOeUMrA7WpXKfldUBTDTdUuSf27VXCvqfIXHNmL/slyaV4H5K4myr
MUcbzp/KzbFm2dPE0idYTvkGA/0xfQugLYjAgwrcen/Rh6We3mYJdcAnFWnsYHsj
GutAp4G/Tb5Um0wmGaCBlsuvT55dtzww2QqTsk7Asabl9SLcP7px/lpe51NyfiMU
6ODdYF4CZ2tQI6pV306y5/dCt6DsaMMUiHlTAARao1aenuLFaiL+xl8u1Qfx9m3M
SecX7x5B72Z6VOwDAgqKTbgWaKMn/9IhXJZ2TspiKlPWpTYe7KWSYwt8DK7DfWzJ
fcD+kp/oBbaNoU3Q1fPpQVhdozOmR4pOnAud/X9aknSpHUVR0Om6Ei22NLQKVhud
9MAPgxd2Ps+EAGaJIbEsV9DuZKqWBFzxZBE2zHRFo5/rL8a36qFFEog05QZCU1He
ix2lt8hp6sHZtWFD8k34wr70j+45E6IDMEQcVYLrvYerqUE+RnqR9ZFvogeYVSYv
Y12VfiOwI8uVDqFYF13SQ2wlbQDzlHDxnF+ah033Nyw0XeZC83o9OUKnpBUTVe8o
3c7043KTeVcqKft5pErjdtTy+BSiIuIj4lkR8ncZCkaWo1h5rngGDcyBCHDqSZQK
vPf7u5a8LixtzvsS//JbwZeDPfagXBEUtcNA6k1vQBIsLgu+GoVb0pFsfE7x8627
sXY2Y0/tTBghbLHbx2ij1p3+WCzNuAolTMjy8A19TbyHSG8ASWT7lyCUHU1NnnIz
49VM2jqi9aMnuhajQVB3lmpJyhuw0yioc0Vr/99JBre/M3pkZtDqyEsNTWx1omJr
difyNc0qE1KKv2NRlbKuvr57KDzeOtrQenoTH3DgHIL8DBT6d4sqHmgvBbFbzEb3
zlGGYcenlR5Xh2Z3rlAAAcJ49FRBY+FeudpSQHOoU/YHLBZIAZnaoTvB+raqSgCc
HklyNqtmCf0SMnzODGc5JS4jNNXyT0ankmDEslFBfy1IxsA07xBrRzOdo92iAhfm
HL1RE+BlI5KHI5ZaIDu0Es/76nmPd+dgnOluoxusF3xCI7HMaLsh2COZJu61wqsv
92rUyonRdGvWqO47NwixDfIE91u4qSLcz/8KE/P6ttZOX42uq1LOjGpa2mRQy6h/
7zTjJgzXatTpg6gxmHsm7+y0XX2JZ+wUJeOt0hX16Nvncv/Mfbng57wsGbXFLD+u
LQELQr02ZQunpnRFbJRws3/NN8f6DY/QqYxU7GNtyxM2xmW90hsEUu+boaKbvfuX
hdjmGiKMEllVBW6l8Z3cS2bG0BYhFbj7/dNJ61/p9AuUVg5jL3SE9knCUxNOVkzW
7YJXgXclGm3nI+82MlfgCcfmI7gV7YVIVDXq46cGndY1s/8j+IeqRDHjJFrNIAHz
V4BGkRGDxMwHwLZjAQobX4zKdr8vL+KTvAvSnfcKdMwdJOonwuBmDqrzS/o6N9rm
pIAoZWW8dqrdgqi8CMhhJyRsPE/FIbHYQXs146PJ5p0wDAX61kJzQXAA8uLJtq6n
NpuROQ/6QZI59rnZCw1tpbQeVAM4T/n9GvE7UnArGTmbgFcsVDAdr8LhZpfrB7JX
jvC7BkYPqAFqlZEIQYBZOpjSkMx7g9bPnVwKEctyYFxS8nDk5hlRtyLzwPuBQkXH
bt3tL6a63VlTOph4LrUm7s/p2h/tfogf9ZiDj/VU+V9CrupZyvJBKoBSWN4SoO65
h3F2zhR8L3droE51BftF5ysSialWEhAO78grPsTKRv59Hht5Pzd/zeKN2ne9ng0b
WNyNm3eAT2nfyH8r+vzDy9DdElwdVQz4caRz9/S+peLGDdGib4/R1h3rnqByLzys
SYK6J+eXXwTStssupro24u4CfvNBOYq3RbllarXCRCCSkIpT0OIP4DjtDqZOggWP
wPrr8sKMmq6cl17S8TuycMT3RduqZM3Efi0+Zm+iQIjHRa1St/7OMCax2xRfs56D
MasIq3FUBV1ULAhwt32o7qNIexxb8MjnSTstYsorBUY1O/7jYwpOF49DadeoOmrf
taZPH4NOn8fzyFY0RerpzIUchG7IOVJFmjh+0YqPD2FPzQTj9CPs/XEAgomSdlVU
5vYA0alKd8cnTV4nDDftGgdQ29KUHHqkgKmfL4x1ehS/u1zmbimNlHgDHaCBFkx/
sosvYjGK1ZHyEI3VGP0pVAb+c7qZUk0vOeleeoDETNVX5BT5lABR2iQk313ZxnI4
LatMpJf9buCFXMrkSlw2r1Xv2N6wGhzy1yB4X7nzwXQv7m6phgA4MNir4TZYAv/R
SVGesR5qMj7TbRs5Hw61AVQNmMNsoyJlg3D+wbVBSdsj7+zTeqiHcqE0kr2ugiaE
x39YIZbt4CQoA3iQnBXlihDDolvg13eOA9H7XPKYSsuK1zqIpcZ0mO/irmMgk60d
9FATjq3IMwM1MO4ZOsJ4p8LAfY/aReG8QeEEa8m8rbXQR2g4yc1l1EwU145Ys2Cf
X9dij0eOmZHZbH0jz6wQwtT32/GIrmTevu25OhMG+WKJRqrgRRVgytKvvCqX6ktu
bMpJXyF60Gk+VTAKyp616ULPLAjrkv3vnt3SxiyWIPIYgbYKYPx+C75vhG6BVqia
LhBwbA6dPovzXqTI4OKu5pSq/mxq56g2g+3U6k8fF13x8NUc2OmXUzntYNppqD7V
vXNNWVD1+JysyaoKw7rHZT6Y/t6sBZr4dITNXDTO8hsxqv1zKs078OFvysXkDfxD
4a4BMARz8Wx9V0jKgA81G/cttC8FFFXHCKsaa3UlloUtwPEiDQJWWcs4mA+SlWHK
vsmysjJwNkhl0gXR3518StSYIYbOE5T1feY7Y53HEfJY40PiLb75yI8lBGZgvWGK
MAQzANvbvSwP2n9Y9+eECx5EYiNPiKa1IuaG0IZjd2ZJqw0O+Sj5J8IwgXBP/gXK
Jtt0zx31Fgfy9zRkYhqRTZx9cTNFTa2udByvbzlS4xhXC6DPbE27dwzSG9NCOmiM
Q7+fC8caKh/n+347F7Rw0Q4ccA+sydFRo4eZ4gWZsrJcQUm+YyXreKo1Nu82OK9Q
p3SBINlgsitpfqTUc7sIJtGYlvaDvC/in4ICFZbJZroqJFi5+we58vFd5q3FcH0V
eAgXtLP8tZLbFH5aP61ysk4gMKORRe4yPHId6C4G118Mx/yQKQ23GfDbNh2eNe7q
Om9OSlpGcKr1RfGSqeZoAnTgS3vLIdrG+/Y03zfJl30uZp9St8nDNWQEIC0EqMXo
3sd0jBRXizb3dPxGw8SODepSJo3lBiG55gg6hdnXZx+/QxoqyOVhKLJ0LsYOs3rq
rTMmlktFB9fiDVEuhaMmFAEmC2CQlmYM89weX8bM4iBZP68cuphpl/SMAmvNPhhc
Q/FAa9giuxag3wr9k85L79LbvQwSDg9MKrLJadFqixdblSSDzneVhyIlvuhcLFEg
J4D9ZXlJ/gk+WGJBKZ4rTEzM9bHRvHOKfmaEPvwcoZaxxITUwtmmTol6GUMQgQOo
yA205dk5EefMspKDiasLy1VPZn3PyEmQlEO3F7mjDhs3dBaXlJ0vq7OW+S1gJNr4
Q0rrJ1NFtUIW09WvANWQYDrEkaR4zwdOWUveOKoOf+tlGfSYGjIovn+s1wlbq9bb
z5LWzXq7sv/qcQqAXw9uaIa8s0g/7bab4unUNG2e2eSrAarg0T+TZ+cRn3pA6jR/
G3scwC5If8SK9TRtyaM2/OmKDTG7G5Qjd5W76r8AlZFMzaDN0KUqtvfdrRrTMI3W
j1JYldaX7vTFQ+mLDCNEQX30pLsi0qd7JZE7VgKYp1h4n5Kp65y578Od0tSCaQxs
ENr/trhMkqz655e7lVHAKL1lSkBAkC6YBul0ZbF0YK6hycrK7QJB0hBo8HzjoypF
vTT8rFdnP3DhRXqX4Pk3aGnRA4+HG2+By3Jw52CrXV/VmKxLE5fp7YuMq05Lk0dx
IwUMAZYstPgoQ5vzaWQf5kat9TOpQBH72a0jkTMg5IfxutOzZr7l3dPKBzmmFz9B
sVI3qPOghqIeJXMyTnDA0qysQu+1b1xbNBHnwFyIhLqM/Acmay/lSE3gF4pQjbzf
Ox878b6vAOiho4KyGmJoqyt+p2EFsTOymTQ32gUzEUVCysEzpvhKNiZBrZDBGJGE
OnTeGB6uqJvb526mkyO5ams17rpsXCtQqyG6jgpRCrRnw/G22gojg2N+LrUDS9P4
47eeg5rEpCHZny7RQ4UU3wnj2C5gS8ALcLmwfGJJSeqyZYBitSanS+kqMuvY7E7C
UnCmnxEKV6jHCI4MKAKjPvr4rHgrBaipxC0m3o9Bt/vBgAVwB7em3ld7ZroRE1T1
G+8I0kvZ0ALYkhXFKhKqdRQj5jyTrtNXuct38a12NQpONOaj3YfbAwMPe0JKmzSX
AX920fd8315DF0rU66Ie8NwndEFpCc/7e2tSChfGfusAgi4VJXx5/7VJ3cgA5jr2
7LbCiSiKXGEqR51qlSGYrqleToIBzPk3ByrJpia42Q8PQ89NDdniS7LFJkbE5Z9x
+/ToHzMrD3IbDMxMF8kem9Uq2tSUNoXKp0tRukNbcczbJiW1j6wu20iALmDyVORo
yOpx487LK1MxZ5A8VswOg7WB29OjmhQXB+JIeDVg4r/xb1qbln4WCTNRVAjXQFT8
HnZRgVuyNMkFiucJRikBEvcyGBlEnDu4sYa0c1eit85QpvfzihqmnZw94NVLR5PZ
txmcfA07/nJK9gtSaipHgu8kgXrY0I1+YVgH9nxw5iyJB+Kojhue5kFbPeL/aoLp
+nhHDXncbdWfGJs5Dye+64lahEJ2LlPSjbVIDjQ8A/ZPMrU/LSyxlNkqHD7Tr09l
5YUkmdq7rfgIltX4WdfNYdlxAszdCqCSoOGyjpjJGs0IP8iROFrjq8IS7PSxtlYo
ihNnscD83zThqlEp1YqQiijx1C9DGZQi1YVMAo0Ug7OGceBXfMAzw87eRWIP7YLl
ibGwKr65bGXTHQXynAa6PgEqndZRhryiaSAA58yoSfqQaSYH097Hwc4EW66IuiA4
o+ExR2zxr6SDMmpPZEgUCKKmneHDap7+x5OY7BXLRTcIOtezNo1kqMjSyRkITV5D
ni2o/UGJSnr7JuXI64eJzerEEI++til0dgyWiFjAkSJjIfwZ2a+3oD9bAyap3wX8
SkRaUwhB6YMNGBizpaXgjchOk+3cm6WvqOM3S8uWfz+MVYc5vkVkCMWW3fnai7ut
m2wePVbppVjVmfGOPwb8OEqfibGrPqpxJVeGIZ7Bpc+F2VvvKfZfh1+vqg/nbgEu
1HBehkKfnMqctRoKxAzp1IbfqOqnIzqskCFehR/PqcmVuHW4UeRMZNs7JV3n4yIy
a5JRtU/kpREFEGlM2Tnp0vMKd8JE9Es7+wuFxutHUDbyHwOQ23dkCRJRcQwFkp/I
DJDo9+yZfUjuhUnIUesi3IeKSU7M4jbn/WA8asc82/frHKWd5eORnT3X2TPfz3pF
duASLqa+kij5s4AF8PDsNpeBLp8g+SIWStmJ6NFTvZApJyGEl6OzM5peuWFtikyF
JXQ0z/yF7Za2pvSB/yPaPNIkewwC/57k3T6iJpYonP022auO4OSpd8Mrpl3MziXs
/Dbg88IQ4bqWOI5CBFu3dhHPyvKRV9HBM8Sf8yWPpIhR7O0oeJLpEbxl/4ukg6Kt
Z5im+UK2ilnbHmgCja3QgJiqQeGBu+T/ismTQFBH5CAKv3ATkE3MfKFvpGKFuwKP
v89zCuW91+ATRy6MJHAPEDAvKOcclO8Z0yw7zDn98QWIhoSmsmyjTX62EguvjcXd
41up0yQ66x4AilH14cDvYsp4taumbSH+656aLx2LOmhibEdrUkcpoO51v4Jof+bf
K+w/CCi/Q3n6HWB22t6H8Trl4YizkCZPWicM1i8PFPjec1fiQGEuJueE3U2yO5cK
OaCechQxwjfVzM/NAYLidqqjor5/5lrUlngISN6uCI4vhyHTaG0S5MBM3pPAwbvd
hZEPOzcidqDKqdI5+r7uVrHWB4Ot7WgHr0x+ezGnKPpj6342PVk41tOsu6fzwgu/
8IJJG6FZNzg/WR15DNSDRnW/WEp9IF8ygvziYgspKVKWjz9niBrAP+QGLWnVXbrV
I3HIctJtaG9+Qt2VoUP56nDHJYmCMmV5jHtWcnjgb2VlUCiYXRkluHcjk4j3P/C6
CP2ooZ05z5WlX5SvQ8iqUMWo5iQBlYaIJTkpY3bwxwOzkl8XmA6E0RmeteazbB8f
700z8BL6QKOxVI+re2+IUE9aLumizZtvZyAiUSAnrS7MlJjX/W5f2Gbd8JqH1Z24
iRtaGwo2iahkO00BUttCFNGg3Mb/h8mZ8bKAj5gPdFOZC5fyQV/bTKHNEg+JpxtU
EJpXWPYMmlnHS1Tw/+DI/SC8R8tLGeVPrzBbOQk/4NC1yj7P89AIUs7KOxWsiIbx
5uNY9QY6+QsKqumEu2QTqWFiUt1Iv7irwGX/YoDj67OYtnyAGLZad/mRnuue17wS
hOPpO+lcqupp03yuHyZniQMBlZxasrEhKN+9rTnHpAXyXt18FKQb8AUXFXos9I0M
ecH5r9WxTCOn8thiZcud4tZuRel+MLHLAkCsSexKaro5P3BEH2AojaDO//8gv6TK
33vuxNm/Q/8YsD34cAiYrvWcxp6uYE96rU+pKUu2LF8IrM31K1MCatnRqqrZVvAi
UeUKTiMLY1YG1XPewT+ybBc/DgjPmn5uksvGOwZBHWgWAtGVNfm+o8l9lusAvIky
AzfnbBsdkM7/KBWxeJRSvWKy1F7mGv7qEpAggbDWvfKuCJ+o1F95jTebAdbsRgSI
hqAO7i43eNyr52FhA3qyDB031V4+IXMZt49dlOlc4+42wy+30g+Vt2L3M8vRlrDC
siaO6DxOv/N9kK4qF/jquNcwti0qI3/0S/Sej75VoLxF0JTf0zWcTA0k08WMicqY
CTzglZLL4csyaK22fcRk88Ujq2AvcRpos7tH/sbbK71ausa4WujRXjaA3GwPdacl
uVuVoGPKb1LHeNXdyjGuSaZ+058nU5QVvZCiZIE3aeMgwCnuvVUYo6Nmu4ClyzAD
WGrujgxX7Vd4FvVxdgYavTZ8jJKHDCzX2XkOcqTOLjupaSAkDhxbVzAbhi/WTAB/
gLg/GlB20u3Fxr9/RL8BN4xbLJTIfnZ6Ce+zcECRXMVA8X+myvcJxhim2Egerkka
hZSB70NZ3F4oKEJ3ZQkxaOpEshZkRrKjujeqHVzBh8Bj0ios0qQlHFzJI9zat3jJ
i0WfNErrMyvUZkXvwCz6Og9R9nd2pWARbsUM1jlHEpTLXigsqrF30BP1zTv3Bmuc
amMoIvwKGIylE+efXn5BR8HiGGtacJ9gyXwrdaGEtWtZ/AzM+qAqdjOJKn0hYTxT
r5BatEWcY2Xc02nvM1jXou2WcSJTjjGHP4JjuMmqXjH0Bgzn5Op9Ev9iK8fBmzu/
8U+lNPAbyU11cwli/tSa7Uf3Rwk3NvIu0tihEdjsNNrlLKF4QjMM5ar7vFQeDJyK
RMzMDFcibti1xSEwd4JyU/J2hSw6TgkP4znDVEn2yGCPRudglyx9X/pz9/QZPLld
HCpOwKsXzzUOtAM8TqRD4K0hfbO8S7+4t1ChvsDXAO95t/tcxQqIh/OKd471uTdP
8cTNRLh0qPG8jJagVwN3f1lI7hWtSwi7vmwl0d+gzzs3mDB2qeiIcxsaQITqppfA
tLqFCcw2K5R+sNkw4TlZueY7Je8oQg7j/rhO5qghDoLYkDfZUUUFfkwtvQT8qdD3
uS98X2MUJ6lIvQXYncaJ5I4HN1nQfKvrkut+KDqw4cgORCviqlR39GqTiE8aBwyL
aTLhYQzV4tOBBUcI5OBcG/J9VpQ+jC+Heu9OQyWtdIbx4KaAqdWa7NVhJB3NCwes
4KLn8PEQu1XGavN/HS4qapfe7aNeuJ9g5Ajw33Dqkwmz1WcswAO2hxzahzWhIjwy
i8Dk7VS2Nb6y1IQfDDMOqfKgObXR3UgGo00z+o1T47gXnwc4cootEHrFjzt2yhet
bXj1a+MgaW7EwQ0pZK12pNxShYeattvebDDRXhWrQrqt87lMBWvqeP8+k1u7tdzw
TO36RQkCWv18i+ZJfjPY6D5jYGn+LaL3Q4P74zI6d98l1btNp0JdKaHr8yUeP/Q4
WN98DcfzChCzmAIAdvkTqM9ioYVAC4o8LUW47ZM7926z8JMO5uOnFsGdbbyWPEvs
HtNPnovEG/gkQJaBdCw2Ztpu9+Oj4fgcsxa2Jp3KCf1wJulGkkfzRXgLtQO+IbkB
uPdVou+HQSaynDfFUGd5EOujhdC/MUBhzp6aB/9eBtKpMgzyW2T8HmCkjPf00/yk
WK9GpyK6KtqvAI6X9KzLcWRerMtRPhpqLP8luRDFWU3yBRKcFKU5bo1H9GPvSiUZ
ef+9x8jIhI/IXgSgzNmy0RpTVGm+/gvRUY5yZDozCYS0RYkXwoYLz4RimKz2QOUI
pLqDg3/zps2s1LqIojIttwQFuCLoUCMMbFdb50TZ2HntcH/FeawbgwyW8DhdWvAd
FDa4t6lcu7oHoeN7w8BP6VQy4ia7sxx0xclSrNjMBjdkJyiiwX5Qa20mht7Yrx1S
JJ5tqNZbtPzBH1CdpIN0pw687fJE4rHSRFwcGdgtt+0GYnB1xbtdpkpvUltdNVvc
ZaI/RP/sWgkJKBrezAyrmROLGjz/zdB87xrFrPq7typHExojAPXFneDMyDmoJjyi
uL4DYfX7lI+w5YgprMvluJHcJw65F/aJ5JiBobPLQxhdchoA7wsO41QJa5LXM/19
mmd4GESAj7wzFBEWZCA0biJog3y0tTz/4H04nkKjmSoWiUSZb11i2xRelaTamwc/
VJMT/6pLMAV9ZzI4S0KDHgZUXObdVvm9d4gPmPqUl0bLt5KPqj8Fw1fLx6Abx4MX
hVlqgIybAR64+jbcoAQAyxEQ3WVoKe/zFEjdKv1DLmtKKliMbXeqlkeA/sM3MRMh
fMXyPkxeCvUzhYe9lO0xPY829KlgnixCfBqM2RLuCe2EoiKDIq3E1wDINK7o/F0i
Wh2DeXzaKTQaz6c6PWQ/k//2OCa4bBx0HpkKhnsKNE8Bu/zZbZijKx7BNF7QTpCp
che5tdWfvLbFlgyHu9mONujZH/oyHgI42BUJd1BiVIj05Habbdd0o327YkcFTvTT
5Rxbl7UV9kYQm4JhQNTn0GuqwqfkkkrF8+T9j54FqMMRct8Txu/VQDK/ykANtTeM
awJ5hBas5eFHXT5lyHtx1PpdizVWYMftYQFedG7k7tiSrzbyjVKGzHXxk3On7N7D
YoCa1BVylIWCaNQ38RjRFY2hSp9DESyZektRm6zCSzLW2QfTUNxHQeRzyYZfXBXj
DBav1Rq3C8lxrUlN+8j13Hjx0XR2nUoxp/0gafvohCZI/pQSxH/6EOoKCKwBw26f
eHgAozFMBvwX93bKdLIsPdWRzmHRH9L8Skny5u+wErzvvivR+EtkN+0DSG7RPt/K
WbdH8RPS2AvKskScDCYsAZI45mLRLfPqep5HAYLmZJ0qvev8Q8QiOpZoxf9oKjYU
2ZfIrqzIhLyAZFh6SDHw299WZf0RuDyICM59qzGKftmZXt+3x8ipAXFkfCi/nag6
Hfob23vF3MznFHGqPo83rQOupzyEnE+oTICJaKbJhE5GV00oGKWgFL/kId6MzMiU
dYQFlkljoknkitjOMaln7WkdgmqckU7VicpoX2PD06wDoN71jXRjm80yNAJpAa+h
pVT5FwmxftM8Dkxxu387vIE4OkkRlQ72SxGIXinHprED6mthLn9fY+72JL960ci6
n0pTALntMvkxkb2SJaikk5GROyZhTysgIX80SUr1UWPvWDKTXomqoYMGcrcWWvIY
6kWh7msfTzjS4Buj7CRUZ5v1ymGpR1QsBmxp83I5K2s+3osnZFpSkUkt2Dutg2dl
7HAAMuCkR4zF/vEC0ShHulG9VN6sJbRS7oFnxX9GlonYvmSALFSwEZKCbBtwnPrR
H5r8ya234UeejFlpuTKiO27wrzJ5TMzsWoc5fQL9dKgXPRKhNXHE542iF98PbRni
yZUh/tg+QF2faPf3cQO2+05OGGSUvlaePDzwXTVghqhJHMRl1xOgY+goK+vnRJau
fwP9YtAdd06IqzOKXosDDqqM7aeaufpvtUwAQcAl9FzQAGeYZIiEUH6wZyaJlrF/
nFBdSIoMZ6pJxB9RkYVxTkPhe64nCsDFJwBtip2bZ4QZBN096kHz9d6d6Os0XEzD
DDMGsNGQP0RH3LjvHihWICeK/gWhSx7NEgHHtk8qr6RUBKxTpr2O3ivPrkLA00MX
IZ8x0bJnWo+HNRppwLuEuwUvcwRkZBJoOii3PA7Kno+9As4Vbb94YmCM9/w00II7
5PTbaUDDhu0tWnyqj8/xSjuR2MmvLDXMAGrfduXX7wbPDqFSgx+t+w6f/aq5g5eh
PvWd4PNhEtnsfEwFmhmt2FSX+88GErxYAp2kJvKzasaTfwpbOPtpxfB1MEhnHsuD
Ck9jh6wunJzuDPe3O8PgUhiVmQXCYqnwdcujhKtcLdxgabgWRbPVYKs7DY5Nl/xm
0MMjVUUQQulLILn162/bO6wMELrrgXFqU0keFNVqWsSgCD2yOF/1KEcnx0prkTb9
wy5PeJlPsZ5hmjhhwoIEa0lBVc9cx04X9u1kS85DHcHNPYCf4trjSHwpKhCEf9Ya
xuTB6RXCHnpT/9S22LTigLWXiYzQLqu4WA77Q+y7UT+8r6d4lt8MY5VCfTNbgqJ+
VjEJoFO1Ocwcegz189eIlRfbRmTc9m+PShxqApi1iMkOtuRpgWQh7a4xa7f1piRX
kzktzR/lQQLTOaViR6PSaQYsdew5GyoPGZxg6dUISP5q1E7ka0rE4XleSI8M2Lt0
n96UxNEtYMTwo62c8hM9IQ==
`pragma protect end_protected
