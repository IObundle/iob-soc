// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BUTXP+rLS85OXKoPyQ8Fqvr3EhMxehzRTHivRGvJWivljPXXfst8PNNU6qRUW70a
x2G2B84eOcHMCWRUT7qlapRIyWnL72RPzS5ezjQmgaAaqirCg4nLpI7n1YXKpgDN
WJTWjHXrtaF3wxkUpJ0zHwIOg7HNKUdUw4dEEcFyEb0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32832)
yFQOduTlROMVzmROudTanUPJ4bIdgu/6/MiDBsJb6Z+Fz5SFe35l5OxbLJT0HnyA
sTcpqYHDNvb6Tys/NNAAcNB9OSSjTKFdaQZsriStqsEkUAwRa7uHk/DvT5lWp71H
ZCvO7gHoxAAtbcR9cw3t3nj5jR7LpQ5ELQgUGr3mGOg489EX9wTTj6w99JQcLRem
yfdT5d7VxsVqfouC7NMbPITcUpxTTqMDr1ubKjqkvEtjSOVOQ/pV9WlYymirHW2i
nyaQtSm08hQNdV1msPusZ6v8PiuxPkJyLegfVh/hfPZNaWLKUInzG7c/cBCQtIQe
cKRLTSlYvj02MSAdj4GRW+wKmXdiXLqlAz4U7mzcoYdbmfjGaJO7YXz7Gl+4QB+h
ddATkl+v4UsoYvnA5JBfZDbuGUI+J4R3e2J5/bH8P30HsDVwaRpso6So9nE7xIff
L6Qf4xQ/3xYmJZk+JKgXKqJ/6HOaYgT4RFCzT2d6fDQaiyl+RYcOywMKBZNlpgYV
mjFnHdxoGZcWQLU+dhGmV4scXBeJO9vNl7UPwu68lR+87CidbmlaUwlQQFdIuSXi
+ltQlk8K3AqeQfKmuP+AcF4q7wBmOSDt2Sc2UTNW+7yeynYqnHHVbM4WUXXgqWTZ
PNX80Fjn5AoExcBWfbKZzH7QSTsr7yxf7/eL5dgJ12IQSM8Achf3I+4NJvVSlX5S
mBHQfUOIqnSGLVVZVP3+YZbNuXMnJ90YR4lkvD46J0iBwpsKM4PIRM/do6Z6HT4V
5pjCpCNz7/hLMX7mNZMxlGNE7MdhtB5hwJLMfXTroOqrFonSqhmdwAOpxmu86VVv
ZX7ToxllC4piEFUaLk3xb3DaqZ6AdsyIB6inAEayJP40jhgXtJIYQH4qHaQo/WTT
5qhkH2simvAa7/SAm5SnW3Uv4Zkayl6KVEHHfvmY2fgh7nM+hmoJALFkoMSoAXsz
yW1H0wE472Pxi7OADuJZ9Lt0DrmjvX8KAAF/fQQwa5z+m6cRVLBaLZb6RJ6c+WWA
4LXKDrLt8iRnLpOyEps1Aw05xFD/TWbvsuDxArOKPuG5PDstss4QEx6UfZbASjcc
PWZmY/uiDApjXsQNw+1jPccq4sIFLDZJoV1afYoXpQtpJLJXn8DdJ4VNtMMFz87G
xZoOd9+Oi5VfJnX+zwVlwjQdjArjpCwM7roULGD/LUPqYVrvguC1b+ugF0uTvHA9
o9IzTIVOn2uNjoRCI5H9Eyvaz3z7KKwOz9ptSr/pCe1ZrNdDduoWYA2WGUsRWkbc
BGjttZas3EW4o5BJQWlcrHIzUEtxgAWaUnVtqOBwg/ArtuZ/1NAil6EYbb+LKMi0
JW2pRAV1KIHKXPZ9p8FkiWD/HVslk+f/OU1eMM68sXzlHcqnkRsb7I0Z3+/kMhKV
ZZNOvp30pp6jeZdjINXremggCpuV7RrxXoZTzR72H2/GWWiyTFz3edOO7y+2Q58N
9KLCHApulMYrCXM25rumznmv6xJOEkTagPtUACSJpVpwf7ESYqu33x6xZF1W6RPL
qbKB0t1pQSRZBvtAxhAEIySKRdx4e9NzT3+hv0HVMHpLgWHbu8hkzxvsVuXsApFg
0mZH2IE+RQHgenjj+ryYG3tOJXLulQHp3K9XAfTQOgDjLd1Vtwmj6IIea5VJVXvw
Pjw6TqgWukpVdSGBAy4KSVVjqvg8tRz71S5NHOUmHTgdeepawNw4YT45B1HYPqNH
Pc3qghERYaAAVTp3+J+f+Rc2by5tj1dJawEux50jb05/yZ2oQSFHOrT0cJwUB6rD
JV+9CJRcmybgCgoequuUJ2LLBAMj8agvIsiqiZxOukorsvJCHYlar4nXZPZbM+EQ
txvsmJv1F7YjPDB+6xnxpYYPFdMlq5b88C8YswisFNnh7ppleIHWX5w7koRZVwZy
RgFVdOEvUyuaSm5e6A6ZLS1OIgfVsiq1dpyYGCy2Qw8u8Z8a+awDXb/tbyapJvtZ
NBGYNF8I3ZJQ6VHSEcCrjhW+DEx2wqwmdQNzeo/MBVM56rFhV9BvSVmcetPBGw5g
pp9PhEoxtLrtfQOTmhwXY5BF7RZzDrOaKpYjIi4+MRd49Y7pOxrTHFdYBS2wpEkk
8wN64Ml5CX/qdmzmm50/68WY36XYfA9BlVEsp2jrlxPFMyK7/s+cEdExmBXJkCqo
ay+F1t2ub8St6OTGzT6m5Jv7ZxvqB3YY2XUasvM667c5TQkvsnTAMCrPoLUU5++G
zLuDGPW/D1cGNyEQR2yrywQbNtJNyxCsQz9/U50vreIrdZ96l280ahmWuj7mLE/Q
X9Cxqd+kbw+DGSxWpimLCdjqPLFqUk9XV4P/Eg+/pXyBlaTpv6Awu2eeVlfcpZS6
z9TRs1TyK2yiEDZr/VgkDnuc69M29ffFntfch4tRJ5J0IKCXWKmBlAvsyCTsXQ71
bZhj3tdE7Nr86t/t1m+AESH88PhYoL0SKEutAg7+8fEN/MgHtFUcxwCqHum6tX6A
S8cdfyV8QIFLd1K3l2D6aBVb9LGXs+4tfx6JrO681i88EB+3fbEZr3Z1eqywZwgt
thtH7Chu7hZNgzocGqVDoiWKg0VqUGen/QXbOZXye9HIPEsPiUOvhqUM70PUWYHK
VV9X7AqvXF9QyZtJis3Duj3alE1XXSWk3xeHXBZomayAWRgekTna1mXFg+4vjfgK
hs+Ep7CbOo0cooh4jqphgt4LkI0GdMNSUCXSahc9To3nusePCxXdprt24hSIf/6v
diJtWz9OtZTEPoZw5gUZOihiYV7YHORKBXvjnR0NCSr67uNNto3V7G8q3ebMOvps
DaT7lcO2cF6vrh0UDX7AAR7hq0g41hLubPKKOkZt83fWzoNY5idm+H9LlXi2zxF5
rt3HRQijzMa9L2gYTJmv8fjlZUukFytzvCMpxpeP8thZlyWS2iGelftbSdl/YGLa
uWXP/VB6BT8G68RPApYt+cNUI+xGMpi3fwQHpnIqbMr2EB2GI/xbivWscI4Ol38+
nBpAWlUL4c5Uz5C90yrPJqOWq2WIE8Lbok0EJ9up8L7Pf/bH1UUPVC0Ngw8xQd6J
2Y+aYB770jGqMdzUPD+81K4e3jaULgTEN3jywsz7NcoyW1NGiTFGMXOFYLA5tCGl
m8dN9vfkIV+0wWh1jjqguwjZUKTQQ4H9zmBBhOXjdrl/A+v1rCVgX73YDYJVMrtf
9AsMTpMrZuAQMmxCkkyKe1cCxOPgzesIIZnUrd3w2+dlVRHsapZZSOoYAeu19oJk
I1Kntf7wj8pTRhuGTj19tNTsUuTjvQPnlIhnFtVBnqYPdCVkxl1No86cu1DdERML
vj30psZBe6SwhPE7trhoywVv0SmOg11cGJ9CO3dxZFpHzCt5CNz9zNOi1oxqBRV2
P6/SjHf2sk4vhsMOldZTZe9fyhVx5hKLg3As50FPlnbPe4p+lto67XxwacpyRoBY
T77Jy5hMSO8L3Ojzp1xDtqZ9shbdvpqjToYLjGmV3LV4YgZlmt7ts5dqlGCkiexf
bpN2LeT0ww6I1/HzC28TINLGxw3FQCI15ZYtZQu1rmmZ3B43vp9eiYUCSOqxmg9R
TzatwdExT1poWd3jMQIB427YoOc/uDpTLAOsCLlVb94N0V2LNmGoB9PeO9SsogDd
InW7Q1gtfjyQgiMz+DT6mNZw/Ac7YgUmaYWwZxUp1RvsqTgKtSBq6XZG8mk/zH0I
M3NZ+5s7ffSQteoV1VW8qmdlaAh78xheL96yench6nIB1hZlRL5Ee2+p+LCg6rLv
a1E2pIVA2m9KVAR1JCg5Cv684m/E6yaFNNh4cbWi0bBJt6VCkn2VgiHfUUSyCTs2
Fby3QwK5NsnoVxTx13Bl2uJtceTzHEy/XPS97kJkzMCCYOQsC+2arlIgeAkNLTko
Ak81IT625z8MeyrVzi0G0NAwzD2Jqe9dbc1q0gnyw7N00Hmksy2C7aLGSF6yxBJx
Gx1N8laSAsL4aAIU1I8BuRm6V5fSKdSyKB5L3o25wMmd2Ay/77/TTyFGkyjq+Q4L
sNAwdZegW9YaGx+X8Qvx2fBV0ppfxa3GyIbopQA5de9FMtneFzV3J8KwXyjo4Pi3
dLW79LiSPlFYCed9aQm8hW6/TfhdKAsL1XhBfPFKSK54bPbYDEBbDZCgWY9d3Nsc
oOcZKu4COUDjzwK+i0dQJvaCWXyauGLOY/mJiF8G1Mw97FjRNEN7sfHL2xHmBR+f
0hMtwjYXpgt0DSP6gsUhgVOSKeZOWDT/nZxXCQ77uESK7fHUmVY+mJQKiK0pTS+E
SVdAuXtiFociEbulmSDE5m/8gXgSMV8PnVS3j7wJk7KtBIECKQW2RgSOq5oWT9Cj
IkmDkha0VYyj3RQp5c83QwDn75Zlb1vuR2SS//Du2lpsBYS9qty1imEnDUuSSlOd
7LgiQahHnFlI8Xeb4+GUvhyje+HNcxCpxiDIazd04Y1X7FF8IBiA6WgkIKFS3zNN
PyN9svJm1vJ/mTkcqiJBiEig6emPomEx0sphFiOlgDF4z+I8B6wJUvdIXolVYJi8
d/l64xOxn/ctRdAaBXsdQ8rbbM4lfZ+L3RQX7Aw/ig8+20Rdh4UU3V04i6arO+kc
fgLgdlBBiWhDpJvHAcxH09cnzi+Ob0WJtdLlWPmquYt+NH1DKPVM5sLINmRANzlt
qfWhOfmMyHGh1VOqGcpRgxk/gUa5RiMozUSBY5eR7OVUMLG9pt/ZafmPc9iDc12+
+mKzpCRvTj+ynS1AupifLN94xEzESfTy0qpVKhJfSLPdSGXFpDh3hQ4USwSWHqWQ
vIoxiRbCNGesOBAbMGlN+yeDovS3hzsCxLdARb/QNWGhJiyt+pa9K3fOJuZtxLx5
HvFgP7b0eayh5adW6mBx986YqCfebYsqVAVve6xQqohW6qJ8w2h8J55fhBD/cEBJ
cz+YmbzjiIApCD3LfiSBnrXV+FeQFS3Q2a1v6pVljMpFOIfy5BtqhK2LpiqG1RkU
5uaGs1l/1DcfRJ1GVm9dqLCQpzJyCaeZFERaRIdMgbDqgrNqnFFwrbdk7gzbtXmi
hbfSesRgdkq7Qb0cTxVgATQmaRCG+XZO3FyKCzW5HWvzbSaUZPgLpfB2xGqA1CcE
Ev1nUBooKFqVUhJOfeKSCxNwye/15yviQhqlzBaTPyFY5n8c/wXXV75aLu3VCKoO
YwhWNBhjO4+TIKBPvytIq6LGH4mQYuHOJg1iPyV6zghtRTa7kHh1y0HkpkXcgV3t
aT+DXRXHFsnOinnEWGd+HjrnFhst3IxeYZFWVaclXjELZa8EKdoVKugHAUMxiL5k
VLw5rlB2n6oWOhiaqhmsvHL2frj1FHRRnH4nUca+CooM4pDJ0zInEOtCJJL48yCE
Fzy2Penb38GoHu5B6uKKoQgWYXuUS51EcgojlPCw0JZCz+zuwUhMpAX+npuakT1N
/ERmXIbIbx2wGkd8RZFMRGMaPufh/npT82qeXwALm7tGngd82Rvv6XeMROE3orQT
puBqG7Y8uxIOXJkJTJboVusv2KQG59pGMb+Tl1FDR6paSTZLqwZzC/18+W4vYhUz
zHO105mNvz4ArLWc2pDFm+8h065lhXBohmtkET32p5Z1Zjg97KDjSo43d8LtELlW
ZW3NikliqVjJNTeoYBIE1B9YIJLYNF2iOwJCYoy0ScqlJelzpiVCwIwnzE0YRAmc
whvkhFWCUWlGUlmBKzWVGOE0eOKt+xg/sgMCtfYkixEbujclISl7m/vzP2YinbH2
XtnW4tSi//lGIz1chyMR5ZRIUt630ue9R85dlv8bkcDkTdOrLu3goCnwB2ErOq3H
/Yltg6PtzVEU4ralIunxpWZx0ih2RdZEpgD43YZqfHgYG98JGJjHT4tAUVgk7aQn
GmeMIDOHJ936A4f81HjUzstttSHkmJuuPKRns2Q5K7dpI9eK+TvKgEyzwcYjfTZO
Q63k5AcW3ALtojBRckixANf7vgUMBLuK3qLlH9PrHKpouD1FLX/LjjikKaEhjudG
e1xf8wfYbsuteBF4FrjiCxk/rpP991VGHszBYY8OHsFb9dI0sIbjOuWDlw15mQzn
SKvDyl3AyddxW74BDkS5Xq0VBYBqwNnjZ+raDWNqSIwBLFB4xnBc+mkPmR5WtbLm
C47C1noJEMexnWZHPstVH5xSJHzstEIMB0cC0BAK5EBijaA6GdlXozvKKd9bTLpA
VzIcemEbunX7Q/tAEtoUBvBzVL7VGTqPusuAb9w5Y2d8iEWV7PmU0hbn3Exntd/t
GC8G3y5my2nxcYKd6fdzME1f2PUxNIPyWB5ycVqgwuxBNg1c87/eD4CDNjMIUqSO
u1MyiJ6ziKYx+dLBmHbwaV6MiWdPrKX7h7jM2KKUu2P1hNWxoLiyopCYdFJCpbRV
4y1KHdhBjOKhN1WFtJp+02iRNf0Z8Myu6q3/C6h59apk4XYbVKt64DPOsuL6hrYA
HPH7BAer3rTdG/r0fl9ZedisaTqHmOC/W6qu8hEj3KZxyoD7uBbaE9fvDt7xaPAd
hio+HMsfyS8f5HhRtPLX8/9mM1GBTiLvNzMB8oDk++OLc2MqUKsA7Olq28zTnu/A
y/F9guwB7kW2yv+2+UOezuSK8uNXGNJ/4tWekFzpFmc84Xyp2H1+gIHLGfSNkU71
PUX34+J3M71siV3XxfWiZdjRm0vUOy+Dl382wXBhI/wYxNinMbth3xlg3SsiwVau
WHi9N0wEd+GL0GZi5t/Xrdhv+LRwSmcaBaPYt+/gFSmhfHPuTiK6LoIvmyvnjTXr
uUt083zTKLVZdyrnLX0E6h9cwARTQOu8fyNv8bSzmjqK+MZaXpw3t6izqB0+3aOp
7KPaJWHjL7Ftfm0BMU0iG77DV8w66ge42eyc03fAWLPe2I1VfGtAy6R4Fsc2D+iz
lVEdkUp/nzhHD+RW1A/daLOnper7KZfqI/5lAjuxOThGlvrENYCZuzJ+1523lZFq
IO1lfVhiaDKCwMQyATyECefkgT4tbKRSSef8QlHWpgrVMZ9dxJJEsNIdmXS6bRzX
TKs57Wnt0kPF4Q1W1zrP+m5mMkSYlEvlNuVGFgSytDYS2W04jHkbMIp87BdRa+hV
mmdfNgZKiQiFH6qq2v7HQXoHRI7fyAuuVUCU1jRFDRV/Fa5gkoARRhrRaW3+NxVD
eKxpODG/iWs7nib4sJLKvce4AEqDPpXQqx4AnD6x1rdsuW7OoPnQS3IM1CBvhJON
wixzOg2gMK/SQkbvN6i8duvxi4Zx4qjxFXty8XG2cEPM/hQOnxCqDTmIR4LmNn20
9j8TsvTyeltd+UgRABwLvo6lbBJ8UyMXWe112Ab4GJ6SR47eeZCnctidOz6+Ga3s
vK5bV6yqrjiQuXZqAitJYgdLr+MHfXJvGukNh44AmNCB+4+FT9hGvy2eI/nVnqja
Wk5JSnskjZRqu2ZrssOmB4z4ZmgSJJE2a5YacBI7bx10ydK4bCWeQTnT0nxjvAWJ
meZgUxxRWR/vGJtwQ3RTPwP9J/Pewk40mbp9LBU4s3GmIsZzWFAeNlAD1ORfggXm
rYqw246+Jq7a6XGjEcQ7b0tvD2ocpFWTByQJrtnc8dTBS73SrzRe/l4gRds2XoTO
oOonyj2EgK2xt5g/CTofSVWTrkI4EP3zTWSbY4ATlnqOvWhslKu8IWbnUDhcNB11
meASOiG2Cqd1dlSVFaUFb2GMfXqPIfewQlzcWj22+5aN/59jzQKb/gUmcOtbrNEJ
k1AW+NHx+tPjYYMZZebi2QaCgV98O9Cwxyzzubxc0503UP6YuAWPcR9lO6UaZeqn
zGHkDEOcrysgxDUxRPpGD/7GjJId7XLe+UQWT+OOdWu7LWlwhJVZZzeipTgrwqf+
LkmZTVTm5J7MPJ3/gGsc7X//ETcIUOrKqITiCPaWaVAOD4yaaP3EWgzgcNu6bIk2
QttLpK6yP/DoctKNVhnpql/jO+l4lIxmHUzdikzNYEQBb9S5J1rb+BFCBChaNLSc
QoHloa9O08y79GTMJCEi4IsYPv3Jrz/Z46/KV0imCa/6kGYwmr4V+7RjJ1X/KN37
knvAuChcw6vk6pkiwHGzrvdO2VQDsHkZg4bshyG05Cmk84sUASX4016w1+Y9Lg/c
j7h7WqulwYIRDk97eAn6VhUSRTzAdq/QdnSc3izDSz8FBpAdT+Fm84t5U/4/vMcj
OvpAnNr3+M7lof45KS6YGT4mSPBD88B2eTliCErJWz+v+cT8WhB+b99cPa4YQnHr
/hRLLe291N73CU206wSw9KOAcbYpHoKgWL4EvWJ1c0A63tutnhl/Swkdwy15D89k
lgQM/zC574XPVmuQ753319ujLnQ2cxhl+2Pzq7UvcgvQgSR+0OLmFz+6327P7IRP
y/wPo6mj/v0XMTgy2TgBe5tVMeAJTiMAk4AU/Shwr5CN+FV5aGNbLUmm7iPjDZIx
1QaIeyfAZPhlBwMIVAVXceNU9rQtLJeC0dYwdc+CUFeA3FUxsmxsfJZWllm9KBuO
u30uTBqiowOWWY3as5MZF9eKdQnh5stk4ekFwM7hAsnlzdEdA064uv4XEjt1nuR5
GtPe2Gw1BhZjM7Ox13NMTta0JRvqhffL8ivuZ4Ef45zzmeFqUejdS3qAQfJuTFbw
ETKSg86kFNhT5UdZahggijFtOfdQTR3twGkML5w6yNfg4FwA5YR3xxxWFoePIGW5
OZ60bq9r1UTIETsmr+bYDU98YfwMMG52u6FIeffkhM9pPl/xEvt1MIn8d23Vo2tk
7FER7voFVoJWyeQlvGoRXq4bcBAVBN6GYcBKnelOcDbuYnME2nqSqk0BCSInf74I
ltFQ1prIhgn242cYTOsvhDhTxMwdlo3C60dFYM/BLiKJZgNs7U+CPpQePnl67GMC
3zs7yDjvHxp2Yf7011eziniNrtgwf6afUNrPJDbgvrge4xlseKqCavoukUizB+Wr
sv8dte/Cc27pHURygxrDb99WQGsZEDmJQIPkmmImfa7+seyXVRYWHsmQoiUrgAxk
OGM4zyrQmNt6ePR9OZUU2JwscN8qAjGJ2zgMzeW8cuGjz3YP8uc0tNivstp3i6Ra
58LWn+v221B3SVnhig3HbKs3Q3nIoGKWJ5gI8OyhYyY1rYymyt/f2uKiqJ0zWDVZ
aXpE5D6kZT776kUto3D41i1YRvKFwzDMuDEFevP5Lo0A1L2yhi/aKPl1uyS528R9
mR0uL8zMcw4fPeaY5gchXYZB6fcK4Fe+b3OX/rg3PfwpfopKawG3EkYLOq3Pwd9u
wLJRxxjIZy0d1TmzZyz0rNsdebYd1SLoy3vDspXhjrjdcr1fFRnpkDsp1zrtCm6f
R0dOKQrh/M17Qg7QSpSDNxbiw0xRO+A1Eipk7GbjexbX+XjlPyyreEiRZGbAigZx
43n6KsVU3kcFYWdGZQn2advzTK6qfRR2UBF/RjFJ99EREKmHPWMa9HFGAWh9Dujy
2zRDuBrR31L7JOeEN8oSsb8yLirHvNBBTqtwZKfyzNK87hICoI/Ojg+lQSRsy6Az
dR3riLaGirmHyw5aErrCoS6MC8Ylu0FMRkPhG4PQjHCevvxyIBMaYP2POoIo17kT
T0KDFrv8hxwb9YG807l23AR2dwi1cZzOJltb35gWqcH/bFcjz7RnEJjWKEnvaTFx
u6QDgCaSltfyapGuAdSTN/+dH8l7QYwmltgE/U3DwGKKEhh38zIku4lYJlTsgdjE
gc4xyrD3rUOWLHm7Fg5uPuvA7EQ+kr2A4//93Xp6LXiCQqbZqQ9T8ieyMjUXewad
hFx7EEVHFGdOg5nav8wgUHtZxR7MnTTS2RbLmq4NZJ/Wv49y1O2dG+XT8jVQp8zj
2K1I22fkT9AqMlunC6yF09E0jhnCNdzA1xPzu9j1aiR0XcanxMxAMSpJAMwCLkLP
TmUZmCM5K4gdP5rEqZUzHS4r1eKY+ESdeD3ssTlocVkYQTfUrM8HYN/hiQWHYbNW
gC4VZ2GbpglETOuj5McQAJbICNBw+wCt4M6qQpb8cFja7pfBAk2Jge+aYvpeDTP+
w3grQwKvhSqPQZGVStQJRjb8E8k+3iU7Vb0+jPn2gsh684TAJ9wPFJBwy5B6mfU6
PDduyi0KfSNAur/3h5Xo3G87mrkM9+WBYdA5TMyrKdO/BYC213I7iMQ+buxWNKx+
dC5UIgYHp3QU1kplxhafAYHGKGQdqitvp9Bj2TuB9zSPjI7jhxwWp2F4cYKA1T1p
cAX8x7GvPVnCFrTb0OHVqMrufA88EIGzLw8AnsbmI1sdgkuxeofr28KY3Qx5+O9g
7vYmqqbKqmUfPcxvJhhaFMLSZCiH8WrOngL/qn0IDQwK+nq3rfk/MudsVROG3Tib
uPcLoOxYj/tKq8BnNIP5bSOG3xNIUVy7mZ3kmKT7LvZ2ZkKCvycLo+9hTS6mxIeC
GUT5nGHZHAFJIRZIwohBy3UuFBt+3BEqsZZWV5+N2CTKVbaNiMI6oJw95NIqTEa9
3sXwOwzgLoU56nTv5SD5Wvd5ZtrePx3sUbnEKgkYG7Ji8tbGkQq4pk2/1JLmquB6
oMNSRcouo7/9a6fQpzqSj+lmJbJYS3SRABGxQsluT/m5ywNz3ho/tGGzI2EMOSMV
5u3Rzz4bNXNsZtqAR8OM/cYJxb0R7swS0xLQBIFQ2he0ePQNG9QPA2lICDIM/NQV
s/4+W3fqGBwNaMLQ7y+h2Q70DjJOWf7UmHjbo8yTc97lHFeOdJCBqu7nBCiawF5B
JoG/c4+2KDnDeEaupodBG1kF7ryFDpeSCCg1T/wwqO7GGK1RWce830aqBAYAp0HZ
3q3bo6fJv+wDnJWSCfZm4ciYNYqdnkSvMM2X05t2GoOksnuTkK4crrjuEl+keEGc
RwY4y8iUL7OtZ/fAeQQv4/5R2PWte2p+GwHrISE92eugCAApdsjX/M6Qnt0wC7zN
gUTUE9pBJNeLrFP/zZBFm/J14tjND+ja6mNalfEBF0/b4ud8vd4fYscv31Qj0LwL
+4d7cflza+0LBRfY1UchqWu5viHHZwIVNJlijH0QEIail4Twr2UUWoPu4zWJ+2O9
4Vsk5FsTHo7/6nUoMkIb+76ht/wStWi4x2xq3mHKpjTsKBrfTyGJIumnaiK0R4FH
OmQ/c8SekOM6uJVYXhmislY4UWeep3pgL5lwRqShayuqLy1bhuE+MYecuqPXm/Wa
1wlk76xFow4IMuxlldpRpSE627PWrSnv6+4qbmwT+L6/hSqfdmxYfRhh88/O2n46
inL3lVPfsPMKMBtR8DV3JTCGyGtZkz9ZtohRf/rMp8k2Olqi6ZnhTG7ZzmaM2omw
7Wo3gbVpdmeOyroxOttMkmi5nNVGSg+Mf1wTM+mzCOvN94xUPAkUuQpBoLjjfD5n
BLly25yBxmfh7fTkVAo4Ih9IDhhY69pZqSdy4SbNg2bYfmy57/Qif+tetXFzf7cj
0oUuy3ZqtR6LFO9egg6m9/lY9p4tdLp0BwS55fpJZHxjb4qN6rCYaRgimG3Kt0Ku
A7UFXzStpcaAsekITUYzs/hLTqJ8ucoNC/csIUhVxOBMPEwMq8+QLZxxMqZkR1ep
LO3sUwdlwK4xTG7ZP2QyWPxnqTzhe2qFP5+k/FVHtAHfq7uhG+hrGD0AWyAT8YPe
o7dxjF6movv1BNWUNHOUzPyJNFoP1NHAzSqZghf1Dva6YCgjhtNzuITtyqhL8LXq
LLBO8o5qYC6Bwg5ZzaUMdlZB7Q9/KlAtL232RKeZMSWxFQ0xV/wqrBs7dtPsYjMz
fH62d0JJE+Vbk7ue6RrS9oYn6sci/Lk2j01mFhon+czGiR0Q/Mm3Mvjyh2PBbxko
WMfwAc6e/jYFC/L0mYugGVN1INJf36oX5SKEK5QJKpmLXfcHn1UT+YwgZ9V9O8wh
8DMbo1+MHMExCd/ahG2bMsk77NuTrP+OkNDVloRlAj3U3m+pEWQ094GLenE3Ns10
fUdpIFcIM1BuEasN9Udb+CYHmIzmA1psqunTmJhnn905Zr5sSyo8KQ8pRjSA8YTP
fyJy/y6VN/ikNLhcn/asXgHpDvo5SY4CYITn7n1N6wmps1JAVK5tWveXNHcCjnWm
nizVXV1TmvGFK6HriLi2k6IYUoixmtgEWy2RepuIWWvUBeRnqQl7N+cZlCPHpUCa
bWzzbZIJl3wphD9qJxmlpnKf6Os8xIbymr67TQjdLVxM7sKG//ZgRw4LDtF6hp7A
DhczIvmz+Xk+YIJIXuEXcsiKQbaK5k3770YB7cCsPvMZUb5k1UeotIyw4PU8nHV1
cIjBlX+uTv60VQlWlsPyOrVomWUubVOZ1AHPBib3GzOuguOTxTyWYxt6rRJ2uaZR
2ZuIh83ZSrXQnmqTkK1hXrGA79SMFHKJOUsgGMdc2ifKfnbq+FI2fZ2L/q5N8dxP
61drF+OQlNyZ0YTzFQTp3jV8gC+ilG/bOgyzgvkHTCxirTE5i2fmk7HKWGrmRSnp
qF2/8UcWIqPtNx4PC7Tm56e8r9M78qlW6OKD5LMpBsF7LiTKU2bjITw9h7otv7PP
Wg1OsqDmuxNLUqLj/NsnjFVe1k/vgggZQFeeSsh5QptOP/zRFLD/fStgo23xQtvs
7IJf3mQkQZip2opAc3B+JOYGtyuNFCLa1LHeHWTOAdmMhGEfmOP3angu4GVvGAan
f0uofl38P6j+bYSFGvct4+3dzppaKfX3vy18IaAcMNITFjU8UCbPebz7nStiHbI3
vWSddjOu2O0iu65ZaHPh7WO7Je7Jf7azt8BsVcumfwGjouOFs+bFhTj7rblEpIGt
YVUvrW6eavhmBtUPlrzGXb6NHYxoStsuNmKoAvxExxAft+it3lWwrTvpN9UcII6g
6B8MFphzZTgsVrXODcoqmp9KHZgbCrDdNiwuZS/2f2WNrjOkfdA5zDQZQ6vc2o5z
P5wMAQ02VIaRED0Wzc/UEJablf+l/aQVDhg5qgaiGqHPfZmpw+SqMaSuzJcG5NS7
dZicEQV+HWWdAT+B0DAw9v0wBVz52ufch2TCoCN8zUKf6zsbEWT7PlcBtnkergiT
sfic+OrZkpecOmYE75KpZ9jIC1DaDxAvFG7FPH1hlR95CE4FaYR3TCVF5dnAqZrh
8Nk0n+zx6UkdKDShGsTep/4ol2BYKNNLm0Wl/gjGDJHPQFmbzgJm/NR/3t4BPWk1
7MYIJHndj2WZQmYDBSUU8aRehbCbC0RL8aYrr8f0VVRYchj2sJHe/45i3mIBBXDx
RssWeam80mymCYrXeNEImPj7+3J4xZQiw7ClFGh90CaCMq8r6h8vo4VYrTPBIczZ
EPvapR4ROAAQzi1Sbw+2XiUX7IcjEI9g1//ky/1xpLHEBKsLh/9O3TfJviLnbTVo
Fh4uHAJoY+ShVzn/VCv3NVqrPCVSDY5lG0plrw4yQoVtuRQfQ4Z7khJzjMw94Sg8
QwrgKQVpdcJqQUnR7fCjnuXwcMn2Sg1uHTqgHPwy41y5K2MxWev5XblSVZzB4f13
1udxkQ1Gz84/88o9y9PpFAC+M06lvIctIWgo25xIPjzvkQ1sx/Li7vPPjx8ROD7D
vtEo7shuidNFxAN0hDgZ4coYU4E79fgyFHALD5srW4Y7xlP7rR8tIgGoPxdKZhSr
1s4ecnF8A4/rqFVahcfxY2CrFWHcpgwc+berUDdR3Ud5zwHo8t+3qfevFUR4dsuK
JK+3kGR3L0CJeiirze7u+32bsTeeXcwlfejeUiUIMyj+xOtMb/mMOnJYQz/mC3lj
e6qsujWxC4L0tUkn9ylPJdyxO36klg5cQ2ailmB6RnHJ7wXZg0BDHCOtjkPmNipw
dPR/1qioFXzLSvA2FSab+9qi+l8MpQlG4ejOecc5ijrnLSFMkgJ6YnFUmIRpsQON
46I4jFM8kxsOqec9Rbgo+RepasRw45kn/6sp/BRTiayD6Iil7FxT9+4MdOmclHDL
beryju6drJlpF7aleUZsccNzIE6IxgrRtnvw75qaMKC0wp46Q79DqB/k4RThStmK
gBQvK1JdkjaNo+7uRuH17R6Gi+5VQiA/qwv0DjsDyXXW+/fihr35h7/jIly53Hy2
arme1pBh41qFESlpshkWIetREWYErSbifU1zRD9gIPw97YRcBZywKm2BHs5UlZDR
34N+1+UfWiePN5KC7yP+TiFVrDebuhKsB7dxpyESomegpMpXtLeiwMMHlLp+9BJ3
9KrNSGxS52bmyCNcAH3yK20joJzhi97pMDSeYVL1aqywv203mgGA27NDD27jfo2G
WrvvFyA8FwKVnLbbHpzDGds4OMlJAqb7yxNVqO+2cm8Fm39m2lQk2WxqB8u1oBPh
9eUD4oVIJDywa1L0H9SPHR5KV29Zado3yQy+8gDNhsVFQiYPCzWCgeOEbJ5XIsrF
YfTyrh4XuIH1sRrSJ5qz5+XQkfQpd345jfSuYiND+iVnQcKgJTb4YPrcLkbJHTnL
gmqwoHJ3/BNR76XxsoUt3MLDibjnkUNVHcmRreBZP/msnIFylvaYezA1nk8rhmCG
BdS/iHNEDx92X8HWJQAnx51z6Nmpb/TnkRqVdmq0HE7QtlS1PZcTIBLl9eL+VM+p
yxmf80Dh+fdm9b4S7hUjB4Yr8tNwEN/V1ANyQ+KsMsXWSvW9FPEP3qX1+p/18A0M
jYsQo7bp8Frw/29jwyf5YkHji2378GeCSkoD8UxndSHuVruvAKEreARkerNx8CcJ
bTRJhfztTu6dtA1H0QCQkVF1DTQT3ahmaVOduMsMi+k7D5h6nF4fO1tNYebOQK4h
lMnAILzeM+GQb5Mo82Pz2i+HeuUEBHcT5hhjjQgE25+O80OJzLeXQIL3efshDQ2+
gXhSJJJaRCzzQYaWudAfcDQ/ROEYCs4X6vCL8jHt9kP0cJ8blWiHNHyf+oTYoKOL
QVZg/CZr6x6nzRLkcBPGgrWnPVynbuXLN6namC2TU1SMK3H2Vuc5x0kpxQhsfAbO
ZnE7EJlyJpwz9B5nl4GLMa2GnSqGP0mCb9n72S22IHkJ84S0tAgGzpaw7DXa9arN
Yhqxp+d0ac54j5A9ZDsrgowytomhteqMIAfttATpzH+b67JDWOnA06uTmSi3PK5i
BHXzCGpiHIrqNP5spE/WjbBF+Z+sEE8DzPbWHkzI9kkEzrjFs44ZI1n1uoYW15xH
JBl7ypnupJ5UxTUnNhAaWNdworpt/Yor10PYPXxCD7fd6HkJeNgnfrDyRJH2BaB7
lD2f27KOb0u1JEqW5LGZ0yn2AUyA7CNZmxUHrGXlkRKjEhetCKPwUeipRm8fv6J2
Co6azFq2FzLmSw7pNl7IBl3qzIetPYKUXNhNI3UzTBWyqwyGvvU7OOIOn0jsigMn
vUpd92HoaoMd+nO6s+V/fnRy4Dc07NKAoHAv6Lq7UJZF9CWX92eel6dIVf3XVKYN
O+yh1iUGthpFJacKyd7wVHiz1JcNpJ2KqfMiv3DbCWYSvEqFn+raX6BT8F0kmukS
01V/dv/n+kPEocWRwp3RTOQe+uc8+0V29/38/EKVwwoloNhrv6Go/DDWgf9Izn79
h50AuqF64Lp3olKFJf7IwZJaO+9guxQDBkvcAnulsNKnzoOb6q9PcSxiJmCyIbVq
hGzvpmH3im8EPQR07uu+MqY90kOknQiiVqu3ilotgJ8x2QSdtrjaa0OMb4cbqHMc
q5Rx27CeYfrI9N1bUR/AHQycxpkx6NBCuj5+jmh5oj/UrfUFj962OmJGFiD6OuoY
7Y7hO0NKxjITc1Jbysez4XkJ5UHpTHHt7YwYQSqIqt9CSuLUHbJAYRuAtXBR5VYT
MiYrwKKHGTh+BS9dlLhbSQeiJuiUS9Z5eZh94ScqfqHXQvgRJP2l5lcJjXmrY3hh
NKdsOY0Jdw4CCbRK9UZUfjpdoqsqHPDfQUfTBFGOQcprYkxJzE1TF3oRjeTszOcD
ONNNNaFAexPrBFCuOqaHepwe4E7M+wOmgQmnomRXwTP7BWryT1Mdl5CIIzA6HWC8
agsQfKOi/Ujjbrd6n4naHWcAlGQteimkWXhmp8bIIN07Q4zjgemvCFtoZWOztc4J
yrdiU4IDFeKvYD7YSRm+/Ort6rZhpXvpExA+2d5HWmy5c3XKWO8zexU9KbAG+MOn
J/72srrQjtPuNANqE8Dub+82gYEs+6vXEYC7vaBPn/zjdBOYAtLLnMaRHITF4cee
GnNkrRxiePqLL0zoNXjTDLBGDFJfLhvcBkTB+UWcTaDM/Nret1GN21BgeCcZvHT3
gf/u9d0927MOt9zMb186vQL1dHBZgdEs8TLB+a3mYg7w8zamcuMqlpwlRfQvCSHw
i0xahB3zOTf3cqA3m5l2rrkUrB1+BwUDwMtTis72WNy46gm05tMBxd7I9xJX49YO
IIqtcf7uEn0xQlLiKVQlINYrxlOFHQwd440kLMOur/DoNVe0Rcrhk7M8vOszRmkO
wFXd72SjREYtRqNt+/FbPqtlug5XzZuGyRM0MsBRwHhcdzE7FlhiewIkBEDILc8F
5bg2bNe6jZcyI1hWaPX1cAW00lXR0Cvkk6R5KOwKk2SO5Zm38DEwS2nDVfgunhRs
cCAb0SEvhQsUiS09qZ4895sHW15e64ZMScFvmXDk/E+MxTWdNQ2XVUV8PxjME/2O
hDgZpgwX2uE+HJYSBqGIA6YjlY/rn1gBze/qpZRiW02HBx768/gv7kabtgqGs4gQ
ZoSt9SkbSGuiR6VJjGxKZTz3oZ9BspzLISDh98i1NRn994hWTJe3pSmE+EFggBWW
jUEhTZ6G2zmWRhI4GyQeNoqCKhV9YADM1fY/FuyuuLw5VdXkm9ck9Ki3l84Bu1MN
Igqgogl1pZWD7Cj6eiACDAFvqA2TlERPFgIdDeRQ6QGGiF2Wy1d3prRXY3mNQNyf
R+CT30+ywLhCTZiDAdVRPtqXJNmyOLrQAxOB72liQj6uF4PDuMdK4PX2UMrnB8y7
U7NoXXlG5BgOL24m6QTUqMNPe9ZnHk8C8G7VZjOYSq5cWlnvCN0TNIEEy86sN/tt
M1hOnhVFoeyZOtySNEqzZ+KVGb/j2OAZyfzu6i9MBy5WzN/M11JcNRQP7e5ssNd4
PF9nIebVR5JqxLOvC97oq/Eboqh94Rjrxe0ugAmtkpY9D520tlx9BdXPGoZy9jxq
91ckIAEZXA2o4bpqdqjwhDTx4HytV9Jg94TjHhSKZiG3gdbtEV8hSyPeN+6ZMhcz
KoQrESydUd/7lADcLTkT7+EolQVRcKV8FMd+/ySRyBSS3gNih0gi8SzeyNYBk7ko
fAt6JSC/bVDQ+c5y4XHbDDiwJ4zIRe1PO61gJjwjEDC7c7VFY5FxFkJdrGEc4+BK
xbttrXvZNjeo+Z5gVQbql/bmh/K6C2G2a2dPhYzrDVL3PFlqPC54RQspibSuhtj7
Xi/reBOKY9+o4X5/CGn8b8XMv6QeN/xcHGCV+fDIxdNruU0zYVRg9ajsdrXavvQQ
OJYJsIF+ix76aV5nXIqVsq4ZU/HWp9MgmDcC1GVoXfA98XNBqn/XwQao59UU0BNd
NShp4gy35bsaVRTEmKYDBdai8HNwyd+8DirOv4G2fzXb7BNUGBkpbvoR8L8NGEeW
jcs9hzNiz2Dt1bXZSKdkUts7eKjnb1YSzg05qys0nRJUgzd3RJlrE7SfZ4mik1oH
jEn9b0fkzSCCKCsK3bg/bL+Uw2lRnxaaQMHsrcaH8HkIKHVcq9e/90kyqpbDzVNb
XZfiU4Dj1Lf8793NSs6+ofMgrBcXtLf48qOj9iI9MgIfvswOw/IRUCyNmH+caC8Z
/B2hEHxWpK/kjUrVXGN0M/xVHWrsc+1nDgroNFLb7uLqvUD/LLfQvMdtj/Tv9YNv
LlhtAUltq6UTZ2AKLVTM4E+B9kAdy4ULw+oSo4xxjr1IZABRg3ehagLIzObPayo0
wQZOMdcQkRL7QOxQAlTt3gFJB1idFGt9n1HJ3OyHkGOFzqNAYBAUR36xz9aLADh8
dialkpYWfMohkZCx4+hCmB6OGEbYSSeTVNxBibGVw3Jbeyr3DVYWt4Tni0+q+Txu
0T/ZFyx7lVsgiHA7Hl4mmahkEFX+ccU2kdOaUB1C5zrlkx8bGyvK13dbrfjsqFxR
SlSjbuwYanom1oBLHaZ9CSm0cHv5RvCFwfxdzzDPAEyLTOIm87Xr369eqtkQtS6v
n95uwGeP18gEvKxxAgp///LSo2dOoIETn1I/E0n8r5u+pWdJI0tZnlzSdcMsH8RF
fO9xL5e5XDkhi444LMAhBZ6j2JXCTP7wxNW+ficV9AZxfkm580zKzQ/H9C73brOM
qn9kZPWp1XR8IJPsV/V763cdknlb6xvO6B7uVnTMqZ2vlU/lzv9hzYn8ez0CfBMV
YwD3JigJ4iHC4wIpBcAZdwxpCzmMuSpzY9XGv+MBFvfV6LDqI5JaNW33Pho32rSv
Ow7qK0+02fI7hn4MxPLU8eD8qJDCmYSR9U1/EVstquVkNQiagx9GdqS7kXVAgWZp
6zfnIiOopFa2MMEx6bb8jK06LNfkpSNozITH10pak+yGTXY4ZmeEBqcnFDpr6AFm
gok5autu7u5wBRqDemYJW/WXqblEB9tsyOUgKPGXzQ3x3rjbh3cFms9jqRTrJS12
qbMJSEOuGTzMXhvFtD6qdtqNpUx1oICsE0khgGSeMb8bW1neUJL0og/gpxLArg5b
Q0/G2Yu8uU8K55QcA04GdowAziSVF7Zsipa7ZLIe7L8wxT9MZWvdvRhIYo/2e+ui
T+lI8xG7FRA3/uixCeDgUkWUYc33wZciCjZa0+8vk+RBoh2Imb0lP9erhi0BpRNM
0G+F1ZP3Z/GD1e0i86Pq744/CEgr83XD9vp07RoSX/F7EivSZ4XvNG/rTkB1LZ8e
79XFCFb68k6HEsb/nbaOdulcCNJHuD4dK4nGpAKge1g0MW2gqyLUAermzfUUu1AY
4FcSzHKJUfM3TBceGNCae4AThd6AULLcwcxGMNFhXmWOr0k8uLFZXfqZv3Xr62/3
z67KJQkctSoehPYjjyQg9Ese9cxiU1NC67D3kahH+mIOIsRNNzjpmz4viuM/XXo7
uwVnOk+vqrgLbQo9WYSTyvA5LTOXN/s6Ue95E9xkfWjgQjJmSI0+yHPjR/Dg5w/H
xAnJy6gg/1KR59VadfzPStGxvIewca4QWIEDAAWLXWbHzK3cv7AvvKRR/qX7Q4iA
1wr8WyZNGjMtudBG77B/n0vqhrPJ9bVQgmQHV0B8QXDKT8Cv0IcJnkFVblJ1qPqO
t8sFgZ6jNfIL4KtC0rlRYhsGedLQPjfHdEqDc/9wKNLXerznf8tsDpH9WvHq+z44
pBosUt9A3BBfiIgYNPGPajkXIAqTmMPFsHL5vVDWbap7cf8qZp8yVm2zKLAciHDr
NGEOvEwTe7QGf7lP9GRBW8EbgXXUExta2Fi23nL+vrvmp//5KwAptksmSa2RrdUI
RX6tSkn+ov4abSUhQEsAUx2zBIUxq9jo3YbQTgE3mXMn1a/R6zg/MW47aH9/SnEl
DV2pM7PvnbG2yTNQye6LVGzAIyXpbL6wIGIsClY76cqnMWFL+Zqt5WAR1x+nERVr
ixn6A2wfP5SJZOGC28ruAd0eAyJFGoxSa28liT19JheIw6pAKbE/6EVPMQXERffq
pBbsZaGZ5AFOlUQ2qzBBhDOTeH9ZCZKduj7CYIgTPswbu726HWKZoFJIPTEKBPiq
/hnbcOEPfMwZD7dHEeN0OwrBfy8P5NYlyg3tgFTiLi1Dgo+75iaBOXlsZt0BkOYg
ilqZ1F69/GD86bwnI0DI086ffJ7/+W47Wurh00r1Jzakjfne/BwTIjHUBz3tqZNP
J4AhH/abh72ZoanqGLW3XvkL7tIIeu4VuiksiX++q6kCeILPGzhpFuOhPcWUdPvH
8sfyo1a6h1Oo84hXZDNjL2vtI4s5qME9hS3Aa1Ny60NiHqNmiqybO9DY2RANIJPQ
024iObkqrysbUZV7D7kpzv/QcJen9eTt5tEOxvEIvx/O7cmXQya1kH8h0j5YKUHG
nfUKKwo5G9Emw1XVyf7f0LPzdGZhKY0VeSlxcWYc98b8InnhPxKV3YR1r9Yg5Xr7
obpFbIahpydX0GQb1f3U4sjBPrAUlU8LZGKUbFs2RDobA0ndhQsoU0F7iePK0bkM
0sxm9Z2mxK+jzOBE4REZ6aNdShs702GoTqMWVhrKXk8fs61oGwDEaxBEKHAoPW/c
rkmlia9mneRIeMAzXr3MXcSyvqRShnGaszGHshzYQ28eQit8jYFLyu+je5ZfyStH
aPEqMPtZDDVL8tEC6Iqu1GQWXqo8a+E5Zhz6LLCEpSh00vv16B1i0raynfUSCmDM
ufl0EFZNaK/QXbuJYOlMreJTT51l6rqWs0ghJyNav1Of5rlZESXK1MrZTjdCaIf4
o0D4InCstWG1RbLp1Ac0XJme0MOPHci+lZ1sq/HJVV7pqb0yJFjQDm0MgRvuxKQT
W3bbvs2F/PM0+79RysXFBwLiR6CIuwvETPErgYMS7CLfmC3rI+SUQ5rutzrS3Rfq
GoZN4yvpaspDcxXh3/G6paeqme/AMr2Th49YXrqMqd9FDmZsgsHKsKMTrkkbGQ0l
AcRI8UnN1WS07ilxIJSufs+h+yJV9UmM8MllCUpJDlnCIKOeuM4jj/+qPZTprO+z
ojHDroeQWA2rvNuoYj8uSMRPz/6qTERYv6JJ10uFZgL5inuo61RRKJwHCWFYADat
s3pA1OnQpnp9hvh6/eosIV6ovYO1H//boxJPoauyu2AlQRYetzwD1S5Q4PFzoO7F
upGpsA/WhQBLNYBceZOeSaoVwvfsEt4APaXFmUEMpJ8Ac5TOlt9yBxDLZr+x5t/5
mvvrG5H+iNqs1KB4hWECAJiEK996BtUr97QohdbxkRzGOqVpI7ENBvFvG7rh98yJ
V8pn0Cqn+T8C3NNaCh+yGokF6raGjp0L4NHFY/EGrN7ijK1e7GYQ2bgL3MvZHeqN
HBoZztgF1LX3gQtXi/b1QqJnvhvOoHPXyp1rQNl6MNIuD6sqXpGdiGt4+MzGWT+l
UH7MlbLoUATvLT7MBHvfnu5OjnZ1ko72PjcI5P4oSxJpHsuoxyNXE4+UjOwSDis6
2fjRt/vWSX/Jc2AY7dKLz+7tCztAvlU/1/4hbMKnZV3gyRWuQE8lt64IFaHmi/KK
XBxxsVDKqTV5kaLCz80ptYg89SqmwFazKQB/80nxAXqZyyUf303qZXp5lxEIOuLO
8YsIdrSWkUZmwxLsUamYdwH6KjIxxCKMoTJZ3IkSXoCKsagG7gCjsXuMtqQWZ8Yj
L/MWOwNUOPr0csSoQf0BWfXKuIuGTr3yM7xLFpZc5/aqUa49873XoVLOMeqRX5Rw
kTJ5UQwN4c8MDsHNuwEglqkEoLe82G/ATg8HCoe1ozCEaI2cDOeH/2/CqJMCRKus
skadwzYVfiRMWytM9euMHBEAKufhlTx3pyQalwfZ/KbbLh0DvuLlRz1GuiQvo7H7
085E1wU0ENJNOChTk/nPVgjsEUgr9oclZOp0lak8Wd9kUm4Ruwf25mhWh4k/Y+K6
CFNzV9I8sxoF9co8Aevf8Xs0qIEml5Wdvc8EoOEO+fV5WU4P+rSbWaGf97E4wTbE
zNVvC8z5ARWvRGEyxrTsM5Sz0fkC0lc/yBmG0zvXndNJZvim/+zpvyX/dOj5n2sE
Nf60PIUffsi5uoDyfF2BJzc0GEalbIWN1Fxs5Z6MAqDelNC1RWHDfSx46ewW32jQ
xSQWgXHlyR3PCBR9Ni2TaVgaOfrjZlex+Q5wdCpktwvwol432cDPpgu/L1F7YLP7
AhWhCnwGa8ZN/8781aoMvOzDyA5fsZg6aoffXLHLtTIVmvkPpdvqJVyCROCMyk2U
1cVpOonS//Chz6ZuOSe3N98bwSxHBaiZgMoBzQ4tbI/FnfHA/+8l4aLSBazUJf4k
BmDfGIxVdTaWSGzutd1BwN/tMfkOBvWHH6YoMG+qm17/paEeRZ8Q3oRBHgAnpM0r
9LCdCWShXRkF06b98Cy8ijzHX182sWSQto0fEPsoUyF2SVUxxl4uHoVlXCWTeSlM
6QKzqK72bW6QQ7bL6cEV9OABjQhRSwY5VEArbStbX52ISJpKBAk5d8kviP7/X//n
z7yov2ZnWxj31FvPQYTe3gaS2CDfYxF8mvMhyRUDpNWEymHU5FtHP8SQGnwWV/sc
XCKl+DEvkfiYmeCyCXnt2tcJrvvgxq+eNyplYd+mxXRujL35/Rb/Aa8raLC5Baq8
KWKJUvDcWQ7SYZ46DyU5so2s3q2j8nnm1McpGlWMWmAj4rdngySIQtOTuMDkv9dg
scWkdCCuNXFeZ5tiz+uZ5Df+D5XGkh+8Y3W+h8Oe9xKf4zrunfIk38cQI7pyjamd
cyvbiJRbyBig23ddM1SPY8rKSMJh5sDSOVwBoahqDnQHqlfBzWAZRYmDVLLQ8TE0
Cxr/CouWH/arRsr4PgN3jga6ZkYDPTHkH68qUs7J+cbCyPYiQOvco3TTsvom6i2q
fi4rpm2iq5D6Yn4/FLbecleI7lIACakfOltdFSA3TvC7b67mN7hYdiiH6W5Tk+sz
sRoMJw+4fmM51GCYPmtPcflP6Tw/7TeiOIfhKqCnvpKmcjkFwFVu6k+2699qFDio
It0+Blj4CWono1Zup4OOpLlAkuXIsqyCQf+HjIx0f+yKlphaDn4t+3pe5dl1X952
KIFvRlzmtAE1fH9PZPhvtk76ngRcwcT3qy7YwazQ7LnQXhHYUam+OB/xCw+3W8F+
AyVU9TnsLEYQfg7gVLrCc1pZqAbHMxqj+zw0VnYLF2GESPzxVvHOJfbscmSLu+f9
oJv5GczuTyf1MyfnlhmSHZojJNPsqI3HGPAKrMLGNM0fXgCBiX9WWRp9QmC2hjod
nCh5pLFi5wvnep8bfIqiHoTFW60SDc6Jf2DX8ftylKLT8VtmcL2M/9lqeTu6DzdE
hDXHzKn9iM4VMXOlxlWljDRCn49M3oSkuIopZjmEKYX6v6Bf9RfWgCkLpJ0FZDB0
+/+0bY+hN4iaqjcjY1rQjl2nlMUJLITwWgL2eOn9g/A3GYfw8AWOmFAlf+BOsp3Y
+0RGn1nGZkOtrofGakifNn1dMwR1qCRGBeCroKefo7C/7nYjL38FKYvzwkVOxPaW
S048ftUQGYJojh39dhcQZwyDZ6zdAYy5Bk4jseHLekYkDa1fvlizCIZqukA0isNV
wnNq2tuEHXhOKnJCMBiieZsV+lo87Gy9cwJmJnXxbTKEATFENZPtBroZbxJQzXzd
p2DzPDcyoQmbP7lh7qvIWonFOQWMX1RxT8exBteQcMkOQJhGBeNX0X9qy/cXq2t8
kHlkeDxv3SsZAfZAjoyi5XH0O6OTGzyyLzhVDuNM20ENeEfIvmFYmqWX7poelf8L
whpmw4homPNIyyd2ZI54D42mdiqmzseidXzn5b7yrpAcDAB6QBW8srS4fyqutmjx
Yl5nNBo4OJmbB7RUcuUKkEiItEyCJZ4LnPkR5mo01Nu+04WUlHQAjYtJg+Gy4BzS
pJwMaVYrSfCedc5JsiOzmsiwFSQz6RAYdn85q/Wcpg7x72yRYExF+nE7XxJoGgBr
WbAbomRPJ1M5plyDE7l0x2g3TJAMjuzT0kKO3SLqANtjAxp+exuL/Q0z7sEYY40c
FKJ3260hG24fAYad9CsjnjSVbgfUO0ynMESwI4FVTZE0iSe6VIrj5zF9HPELP0U1
JTR1ots2L/7N2zhtv/VUtlx9pFeEy5hPUJdpCK3MAtp0jdSiHeoLVeU/dNo+579Q
25LTKaoQ8ZXzt9fUDOR+NfvR4S0prpbKgjN0YmeJ/bhCt8rgkUNkB+hGFaU4Pez8
o0hwQ3tCAOit5OjaSRkhk5JPFZDDxmO/qPXQz6ZRf4VqCJaVcJZrQUihsLzSCrwv
dHxd2EwYQhIbGa0YNHPMmFwCxLaAWiUSZi1yORMFVBPldhcpFzvuwyn/qbQ0G2t5
XsfOhS4n6icFyC3NHIKwAtPOUdjDiPm8upqA3eMZpvGqr6DYURXKFxG7HuRwbgSJ
JUOLYTbXGdA7aPFzDwYMuGpJlivmz3U4Z6PcLDgyhlWvomx0w8Ib+x6J0AaWORhX
90B8UNF53aG4ick3K/nQ/inJqV8aQxV1tqtw1La3I/vXIfznfzcjyLXb1uPAgeEJ
QN7mu477YTs8geGC1Y4k6thGWJ4g37CuGKDUne0xbNWCNffjiYTEAJlCnjiuWeHf
T0Fs8lzEvlHHvFIuIXRyLcVnir1b+twE/FD92ALGO7oDKtsataIGWOvAU58bV2HP
fTSP9XLeunoVJ65T7GO9xGVbslTPHQ0PE4S2/tC7jrT16jVWrqIhxs+bgBkkV1U6
OOKB6pTHl1lvIL/cUI5xsRF9DpPlmoJloVu3ZL3j79jbZmaMrPSx5xjfZjHvoeRZ
5NQLEzAonqdCvvMz3qPSnBU/yHeSHZ5blQgo16KvVvTjHdosPAStqGyRaCmvijh8
D8f6Bcu6Rzo6NHY90UG1q5tfljqfe7t/zGarNYvT7xipBTWd3DZkvULD1lrpsPPO
uT6Q71IDX8r9sjphIcYmBwVnZ+73zUpH+z6bePxhgALOmWceoXkOK4Q9KwTqqsD0
vHQBgvgTKGZcbqf1MtMhS76LTVlIIatb+NCgyck9gtgsF+iLYa7hqufA8b7IE1g3
eq75ji2S7csw3ZAJ4w9dS6IoFkl5MqAWQqXDpDPgh+altBRMi+PbxkWYLmFLcFya
rDAR9w2vZF5mcnBeJPksaS8Q/pWbAtpSX9tgf/xDA6IMCDF4zkn9QUPwiusq7pab
crieuFtJVfS8/FDxQDSoYNwwtgCY0nyc0GJ5+ZoTOM7EAvCqvLbOv/eFcbqMBXSA
iYRRpvCMTr7FI2v8kmHj4gvuBMW4MBQsg9B00rA8zqmfmV/VRsHdufaggj1JusLU
3mMcP+LMEKBQk6ZgwIqjBYMxfwtCFcfxZNMAnEIYxVorJycFkZdxRfEE85/UBfQO
GwgyG4WICO5FQFeIuzE0SCY9A1ZctVsHbgWdXn1X+gxLbkOGDqdja5kFbkRIcAo5
OzUgBenmUV+CcZbyr4GNEEhDSj0gVF0ycWEDI7/4lT4EgkuxKwSDy8poBMn+IgEi
tfqfULJSYMOfYi/n2suGf5xF6tgqxnbvYKtjzrkhF+fFFYpw7C8WT90Zef218RV/
QD0skA92cW3JcK9TJF5/YI4s16ZR1Im1Hl+Q6esXy/BZeyIg2bxlf8ZaqpJVG0p+
vdELHzfMIzxSiyy+QrVkayliTQOSvflUrWNbLM6cyAxOWo0XmuV+FofhJOenRON4
OgpGEs6KP1J004vZWwxrvr/j8owjHY2OsPQR+sY6q7Z5hlc6tF8DEGKJp1oYFhKa
81EWcK9MCIJ0bHCCnO30kiRw1WHahBrJE4g8RVCUXZPnrMX6qPt8Au7jZIWTJFnX
vYDJbqvBxw4Ag0xLedPoy4tui+SFBOdJf2U5J4YMg42DXBiSozu/Jd9/WeJQbeuj
oMjU4P8yDGuKrSFl4fVcC11PNt9Cz+7bZMKJkxUsO7ed+/fIPtV/pKQfCFbtsyj/
TkKb2SNKsMyJ0ejtT2O46DAgS+CznkgMjUGaFngDPeb4MkjON2XFV3r0lssTZLo1
/TQwv9414joxX0HeiLRHTmXI9i03C8R7RwLrCoYDktBuNF+wjLfoeUwwn0qNniaf
E3MgbiznWx9vhUKvCfiYTf3RaipWOHk/l66kyga1ZINhdviOka/gt3Jj8iaafm4G
0G5gEvF2/pHtDEEdyy4rd7vG5y9h8oJ/IUiUj4/SEnxgfuYN90Y3qZ1YeFFXBwIn
IMq8fooByHwDvcC/Tbzcka5NTyJ0Gna/OvY8i32fuX2XjQh1MTilA+CUuVQAieje
PKgzuAsOwPTDf5AtFG0Lk0k4IQBoPrG/rtdvMSYOC74UInWqxWjA2yQ6ILg0l2Y5
25oHY0V9VqdOp+05DfrPUlQZ2Sp6sa7SrDAzCuxtHIvWJRonAMVVIh4uoJeT6UBp
74t0uDNB0AvBOV7/hhtMXMUJ/fknMY6dYQn72OqRNobHkPuJr/zUrruGzzoOATq7
ROtQVLPitS4vpXuK72IHnN47lb0K3xPxZ5YBUYR1NoL8EJePXn0b9uLB59OFIbkz
WO6Kor9wJuBOmH2Gr/YY7W1e596RDrDtsoRQpZ05/mF7VO+hpCHU154J7Ksq+Vxu
SaxVZLjkieEA3vTqBZ7oFvAssXt6itEB7r2ASLXnoaKD78WFVWEOgWxb6JIjzh5l
6c4xu4BksoLhGXyY82kdIY0CLXINRofAlLkQnr2zkaZtJO85IGqHWh5QFnJ7T8g7
QPf4RUeW6NS40AW/8gWPGhdAK+0sDvE5OyxUc++9eMmcKMUheeMap33/47TT7RXH
SlnXBrNRTGC7gnkiTsPG4AwOJSsdAJSP3DpitO6lGbkJHeE/DckhyQAybYjeDIr5
cu3RnDdwERMYX1SXcXxDDxiRPlDd/3Rfb2sBqxA/jobCy0gIBiZD/ADg5ey1hSCb
ZdqgtkKQ1FgnQPX8TDYWTwXlHoFdrS+pqXaHsj6HtkGvN2XL2Q3ll6SZipIfFXWE
hnPvw2IVfrctmdTKjXGW7Y88YJwW8eekgS2jiDUae9l33KqhyQk1cHXnudtZAI9Y
bMaP2WbNHHwD+TF4bMzt+wD/tOx1mIIDcjLUWAH6y+XL1EWxiYXPF9x8l44sv6TH
LTVneEp52bxLpGJTilqPGSldr3aOapyc241WOryxzrR40OPTdg4+hKCbUBcR9M1X
k3rM4yHq0qU1sQofVQWR5vwjCU1yjc/5e0dgF6P2V16LbaRvXjyek7CDY0PEWtD+
tGjgU4IAhZs/xVCZKIw2OFuwtdx1PKxfnY2kcd8MpIJ7zWOw/G8URdxdICvXtZiG
mOSqTvMMe+p1x+vXGZvtyp8I3XsY802Gwb+VTP6JFWyyoA8j0Hp6gSQ73tRxTP3s
/wlt31P6OPdTD2e3LW4JUhHDfwkJW9TMyTVFXDwz4YhEe5VJ8hH0bwmzE+pfxL/X
ua6KnKiyHO318UzuP5W3rve3kfpVVgFp7dKWLOUw9nKnuD9NfoknJ33954Mu9FR6
RuZYhAChM0+Q4pP+4FxFLCA3I8osBNV25nuzYZ7GPUVR7pctdqR+Fy2OCoR+03FY
oKSog1rFdVTTQ9Y/7lxuEKY4kmLNEhoMpVUY6hEFtoCV0HYmuBeoMGZ234w1Q/Z2
gapytbnYxz0Lt+uC5cxydZyYu30TkPwu/LdZERdN3z1E25vJ7Tl8ZCyxCjge6fid
Vnvbzn3N6SHqJ5pzp+LDprmFk5Dp7cXyEpel1YnhdD96G+sYzAIQ4vZsOtkVoCq1
V5PnuhC1eyUAiHCiIdfc09KO8ZOclRYfmXwE2WkmmjbXbKJDGWsqTucgWrZPLHtg
dF+nLWhX014YsTnv0rLYa09EmLjoeNnccrbh+qUNfXvDbhIJQ4rqM1ETs88eAPD8
H5yRcGYowtuZujSXEBYXXOyNke4jotjWwKPEduW5VUgjnnFRbmcj396TrJgo6WNa
gS0B/hMylkxzOnkSMrzce8ncK3+LQBkiYeB97fMPqE2xNGdRepxFZpinPnzPXA2I
KLgxUYdguKvjo6UzZSs1QBC4RDzRCHLeZh00qso62A6ARz2LDaA5XVj3XLuSgHYs
7B+Lk1w8UxatpwMH3cGO4QPWO8W/7mlTh3B9CMawpDj6ierFYE3QojiVdW3PHATb
+v4PfDTwjxyTRkm2omffZp9kQO7TU5YsTrKxmN5OyBIBFmlf3S2uG/Cy+79ONqAS
vpgfl0eKBqhkAOMXcmAlYAW2K4XEX9ch+1QqKG6A2pLq1ReBBGhgBfe/CVXDpGjb
fDzkuhTe/quYtkQaIddhWwJ0QCxR5C1RqhSVqRKiz7tcbWAmaOR2k5S7xi8+POiA
McrGGGyYGalcmm35wqx28ilLIpjMh2o72H9IEHJ3X8ZxdAdcNaw3+8/M41A8X1Oy
oKKN/QLD4fmrVIfmPIwP2nfa5CEcJnBEAp6PUNWpEGI58z8Z09JqYoiSBqQVGtIm
RxW2yhzJLZAUteL9gTHp4ymyy/UbmsgGSNC+xCfqLwnsV9IzqzEipwDofM98aTIR
9kmoZ93bujgV2SYI1vJ81R+BCwoP2jLf0WztvrkK8Hf2Iws86vzmazqpIiVCT2QR
Ujgqz8XW4afjG09aOxM6juXjYbx9kxQJgtZ/13V4GqdmAJ7/caRnT9xR2y7Go3Rv
A08vNjsQNBeLuWufh0319Kl9QpTsVTNBoPRVBFbSy/9gbfIp0leW3t9yC00kA8n8
LwdaO+PlYg/AoBHxifsvNJBGIVNHWGOlJmTOAIemssf6DJthyBgNj48/n2/AT5pe
ANIl6KJRugh/nfx1Fcve3viskKUoiA6jSXrNcBwL5e1lfNKm5YRqR0OdXtQ65gn2
N/S59KOXiwcDVToN69b5pOlUs9noW//JaOabFMuYO6uAjBrxqk8vw8A8wrwoXe1U
JgIL5Nz6lFx/K1V/URf9SfldFCvrHskAfGF9As47wpfe7bW9AQHdH9PDZNjOOlQ3
zMxlpGvNSXqfp70Byt2vVBhHgQOjHL+EWEGkJrA4IbIoMWnUd4X+2EwJk55Mfavz
q8knABVWhRolgsKe0cZaiCatCJw4Fk6jlcrl4CutMqkEYSoGzFU9Z3xsbFQH1aqG
tDufIk5vRsFiRAgFiBGjFVP+okiOodH5kWmvJARrYXmZgvMqMVRWpEqgvpsPRsLW
yL/EAZasFp3pOd4oEKFW6hgNK0KskKMGU4+ehobhHIDX4rSMnyD/q30IMQxdQ5gK
yumvPWpu9Bt1Ac2cYo1dYAW27LcnnJX4QT3+4WEd/nMG72JgemNP/ki6dntHzRh9
c364yjNIzjJ7rV+ZazoZ2wBdDWXLxtRe8RPHrwpK4EbAR2FntcxMSIeX9mpAAYIK
ImhQGrJVIurrOKn5s3HayQyJIZ5ZrAs7F3HdjFgkNg62AB5u46KSiDoJnZZ2lOc5
jv1wQtW5dKsADeB0r2o1wP9SnnNBOK58wptrF2o67/uPruedjNl8iDJKFy7jNt/1
2eH1x5bbfMtVsXBOXrotY1vmxYK99sbPiobkmE7LFIbwxElz6y2ugtOz8Ph7lCdK
IbPxO2yZMSYQksJLYVEnrfRcvIsVB/Ro1pIweqBVdsnPXgVl0VulKPMVUWJx5btd
3GGHMBc3XLjDj0G/zXyayFTQT4SfL5LCr+7rfbf2B78D5V2AOi13HCXpM95MDD/k
R281IxJBvC63EJnaLfJZBP2XFuOd8ydm6AmePg4dz3V/LXk/fsqutNbv45tc/Fa4
zoqbMzZPlMf8G7s/dIiirbNcQnKXHNpEd1HbITjG2Z9yCjs3Js6B2dpY+FeiqOTj
xh84Htn1jJYeyC6MPU7RW99Y19hpboX6Kd4hnwbpgiNpxZp7/7gBhw2WSc9VaLAw
Iw5EG9WjVb2lpG6GIUmTSXo08qxarpDV5HXt1R16FrSUBOG8XpXB/YdP8pFmc0oU
XqyzVCNqyxtrcIZjI4V47oAqhSPwhSOfg3tI9YgefIfN4+3cNWUvQaBQ/2HmCG0T
v0HubweOGBjCrit6wUUVTNAZCW8BR9yfyoD2AzOpFPYnsFUVqWryD6RwfOHnIciZ
Lpa3NlpP8Fz0JlSBb6JuVgqEOZsEd/qduZa4Vtic4G6eQn4OYtQrhn8MA8/Guo+7
nUsaui8ZzR+CSLMxQyMiUyIlbMLY2whRWkzXBI+yz7lXzmzOYMzlfDMZR0zH2tWx
+odSokPm3qlkdESPoeYzHMKaLGfWxdoltisAuwxFU3paw06MucLN8BApC0h2PZif
ZMYDm5TW+hr+jJLCh39KOYgL78veXB+EygazMTrwIrpDhqCcbS5uDQ1spz0pk0p1
mxUToCDkbT3lMwqBpJ+N5XI7Wo5Xg/hj0sYvUV9KS3ZHTXhbT4+vcsPyAW4wDhIK
5R5ODuq0RGTw5FyiBhF8rZj0xuNv7KoSZAgIaVlokDFMI0GUuPzGb58ur+vzzlkV
8cVsynAGBeyZFdnqtynLq/IorxKbV40AZCgjEu1E03LmhJ5MRy5kA46GlLt/ZCpU
quvDFJ+9Wk+wLWWSqjZQzw8ZKzv2RbvV0QaMbNQhqFwUxl6q8g1osH6A1LXK3+Kp
XD706U0RY52aBkD8rLOoqMeamcyxqXw6vRk8L0YiloupJVWNF52jlJ8rJK1WgMtX
h1WOH2h48B99h/rU1p7TDS8qkKRpqJ423/uWwPwtcxUF9xsZOWXIS6/IDaTuoZm1
0G0Q/0rcB1nQHHz+iaUOWAc9BIq4aR0BkaQ3PwV/80DpBlP+CDBPGwivtgfmVfBO
qie8T7u3ZjZKqMbDMGx8tp/xvx/M0a6C+xK/bWe6lThIz7DCsS5cPkUAUGVFSYle
Q8VHw0MlM9agQqcq+V/WLaa1Qlh6h9P72VsOMJi+rpJvuBjoCVZ2oXkgFSTQA7zI
c6YKLiAasn1Eswz6FJnOA2LM+sLKgM/UovC8k5MuFEww54xU4G503wXLZWlV0TiI
6vTupZgwasPbEZizuSfbWV30w7pzh9Y1e/vCU8jRVQyptkPAIeUlAnJVZScf/geA
NWF6qX5xlOVOe4YH+MMArNFx9O1e3Et61K6r9kFU8aYC5FX5XotsRlUKTOvljeRX
DvAHMN8v6hteLNddkDt5X/ceLFU/jP4Wdn6IG1icRpikXU3+E/K0YCjDofaKiJT1
bBgllxy+zMQ0/NIrexLKBVh9u6UsoAEX8aMRRnBxuvxfGAO4FF/bRVQwnKo+LpVU
4gSWopdIuvK1Avb7Jvr5DkPHc72xrilOtVAGBeh7q5ggp3UeyCZR+PF74U+aPZI6
4cFldSO6dHyFb5eSUZxLtbHwkxVlk1g4tfYy6PB4lI3OQUNpRXbc0O/RUovSL0Qq
lcYj4O24Xr0O6nqXPQNXeLlLbiKUq1dZzquPPoe4zMqnaktoUfH6urV04TdfnX3/
c0poBg9uqnL8QsJUoVMVLj9geE3Gf7M5XaCFmSWzHml6X2fDcTN/tj8v5a0VAyyi
UE8JZrXDHgJmoMT8DdYafhjcv5SZXtg02RF2uO1ZEzR5hk44S5T8ztNL6y3+O1/y
Ia7cQJFFPpPoRdew0bBBtvv40BQDVdxcB8FEN/kGzulenX/9aDMAfNinZ49krKAq
riu4aOK7vEpcPZMAIjP4U1h8esNC0peaqEj9BsflDs2ZZY3tWJhJoB9Snf0rgR1d
ESDnHTIQ9aLdZ2d2QVm8SIBLAQraN71NjLGT30dvofg32jEx5hczE4YV8BPGNQmH
lG75QDnveXQW3FpjH6ncoIYd0v/dZE+5cO/xLKyhFB/wJESQ3NN/rLn9KDrMsIRb
lNdfewvPTMPYAgyOyY/ygWFKWeXdM47LAG+s48F4DknJmGrfhd+ZANwXNb32s8le
rlQrLwaMccKv+NTyT5Ofpc4EQkG0bWpTQM9M/AP/2eO/rmRlCMqmHrvSJBOhxZfI
V9Ygy5+nqdVZrvif+8b61+nbp2pWz9SQUr9jYW1bF22wRXPBDTiUHq0PeU6KXQVi
7ng5C0OszX4XBu0e5oxrnm6rLAwniuc9s2h99Y0HGGAsvu0/ArJTqNqYBKrn0H/F
WVNMP3j68VWY9mD2k9K1lmxFUkMGrQGWJQXEX//pf6EoGzcAeSmB2cN5PoHeR3DI
gGyWayBOAEfMh8hakl6jeo4LS0Rm7IJ3LuxqOKU30yM3qP+f98Rii5cMww9mIEGV
VgCixlHs/eG5qb5RNExNq+6DCFQpUfLkQzLMzC77+fISwFhFz+/hGQU/JUCzdl5W
mfZGlBWUO8sud5Gx+3MLpjXlNRzR8sg5pRlsOq71YwWihRXmaNd32CzQhvkECGoV
HxOFMXSy+CkejpZ9ZZ1pLJ8VCRh4Ee0rZhGU30+Uqg4IAQ+uB1a8LhGMvVSqQOyK
UTdt+RkZQiP25A7rik9Kn/iZtpVNCRvCpqcnt1OgTcI/e+UimfqC6UxW3nSc8c9t
QHVRBF8lJPC+6REDqr68KJvt0u8HNelXr/9A9csw25syArOxctnPUGdH4ZaWRj+D
X9BieaQht68Hx+goRaWagW8YOqozxCrRTQZ2iGT4Cf6LcXgNein91upokfuaVwtY
rnFIkrjYPyFbch1hPS9DXhpLGa8wXSMZucHxT7rbnXex1iLlyRDyFAhoWQfNu1Po
kLaIg5eGF3eM7ThPB2uiHsP90c7DcBQVqK4N8UrJ0R/bGPTHitmk+loUAbaOkHgq
lcDkGt316C+MRTwTpWpCtXDUjv9e44iQi0KQKo/tS+SOiDklO6hwuuYiKqB2eUjg
bVqztR51z9n3BwjX73EWkmOkwLaFLWJV+g6CKMe+uy5SQQxmNPamGe3gCHZsY5EW
1M66uX8GApXoaeZeX6Obo8EZkvV/IhYT2qo3rRE0EMij1Y7aauTb1xuBUNjtFMkU
1p2UiPDVB6rPj2kOBGIqgYYsztjMQ/oRDo6XJwG1JXRqLcgeHNwwcSfIg3SE3djo
zj1yc+0fdX9nfoW3sSmFqRme7NUovtNMYQHZpJfhRcDxqb/t/BRWvixq1bZl/Oql
FzXeUIuK1MhamcJ6Aq7eN/vLFMKn/3evuSUy5zADxpI7zvK+2sK8csqruaP8or7K
qtUV/NtpuILpPlhpiqmWpGpxUlshSvOp74Siuust0y6LGwBnOlJqQ5BzH/MOdSO7
jCTVyHIndnDm2A7JYfLLbIc6IBRe1F8iZZmj1lzpK0i7nv44/827ADGeSJGFfvkp
Cwvy4esru/zsPYlttR/CEYVUev/6qt0K8x/g73Cxef9A1LlNkEeJUK81EAMq8Es6
2ePnfOL7OfSkF4rGY9ebqv5DvlZHOyTmpx7bBceDRlp+s3eiGvdK68T97XFCt9X0
gW9IbW6DR4cXcB14cWVQUcHJPRK94hd+41EV5lcBuvnZKx5Q5U+kfWQP3z6YTEgn
QIJw2+LQa2Vh5/KMDIrXiwJHZzezr5Pm0GuqMaT5sdR4T1DDu7yFtf/c9vNkoKLS
NV00whf08lvlLXnU2qA289u0XbCsQXhYK0Vu5TxTOXQOi4kivwV7S8RbSTWkcwoq
xfKwoyRFZbADqxiSzDt8d23JfvSFiE2AG0XrchHYC3JwOfAccwx++5SzffzAXQ0O
nMn5FVHtDEa0x6b1eX/jZMnOgjC4xQNv73wOcICB8o4XYaUamWOGOppWS4ZBDpJM
TEqkedKquJrUT91vrTOaoGNQW/A6b9lT0+EM+xGcAkeJoOncRe85WNnpll35sBZQ
UhwFS0h9u1twkKTqT67T2KWEF6oCWUtDeNxAKzvYTQkwSFqCheWp8Xni5Etl5MF1
UOlfNc281AJ8JU1khvsKzqE+PqszysbreNIYlJZWZbrUPdAPMvqUeidOpnAOHiMT
HObXCBuEZtXtaIZWafJvaQE/dmYb3vX2MxoscYCr2N9V2em/EB38LxvxGRYkdF7g
SGgVyxbymlGSi9j7gvt7MNaDfnrCa5RVx4EnWPyKtqeWfzsVS+IrlautiLlAT6GV
JSBZNNZb5Ibdu4jSUNzk4QqPCIrQJL5u1b+GrDAsmDBnGyOyXvGNVtvfqj/lZNIx
npKkhVsTkM0ftDHH70y5I2j2QnvVl79JOGwFgOEcqftnpIVSqAe0sNRcOIwvUQRg
kHAfVExBnmLfhR9VIkz3B4Tc0+D2EOmdfDRON4bnX38/LB0sfefDyzxrAxPrKPUH
1KYvfXgMWmr5smjAXiTJoMQ4R7Xho2MUvcR9PqYEMti8OxOwyAjibjTNfPI4+uL3
0xs5lOuDRF0DgFx7oNDdtSVUSnt1NPrFhqBL3wo/BsRjeaVLc5UDy2JWrCJFPn58
Xqakla021ttDTchJSJBCprThBM2tbKXbrhKAZfb5TB3jRbPj3rXKWoI7WSlSzLF0
XCVwaU91Ny1igk83S2lV75lNGizVMLA12GVCibAdOkhmQSDy9Hmr901A9stlqx/n
DA61FLdU+LlDFiH7f9Nhj6B/zOD4wt3xD/NXWk0tKksmZmAMAhlx8IFq0g45wIaw
KkYqyzsQauR+tW68MmHhAVNtTNI50IVLkAO5aILC9x2XO0dDvnhUKGrFGKGpUuH5
sLuzY7Msu1WQGG0CPAFelDURNwk5Ai/xn/kU2NCsHgq2ey7VEzRv+Jwuf2fHGeka
0EkcqXkrw+o5LUY2b0cMVtB0YIJwdKbZ5M9Lcj8C0SgkZYjZ+gNN4vZTHLMTKQzJ
9jy0VyuLUAxO3PE+mSAPSb+LApxmQ/slG9xAfaF9MO4liSgcjKm7gCOSmm7VM3kb
pBpxB44EMASueMojgWEg/izXxH6rjzDfD3WUVoAL/7IElKQ21jW8iJMMXTxk72KN
HEywIFnaH4XirDckRif7IE7qGKpfNpUVxyJBjSHNBv7ipQRh+EdWcULHekd7UKVf
WyxLkZ2A5NEUg8fT0ZyM5sq7VhLZpL9Sfk49ddyQZQKZkaNg5ZNhK3BsQQwcWk3r
3OnqR5tscPuW6gAoRQFzQjEtmcVu+ezXxv95E+wekGqo0R7G2/BnpGCZ4NrpR4uq
fREWyAcsDw6Vm0vckAl7sBfI88CxnDCTRX2Lac1U5FtBmwdcq3PatMlVN4Og15S4
K43bZ8ySeyzNNl7MVqHu6Kt0mr1ipkkmEd9pLc5c9z+ALn3b/Ogm0H0pZ08MaBUK
1InDeL2KDFoIDLabaR1lXqbnhB9SdAbz8MgA1Kqr0QLwdWgDrltKfyIbkJs+9cv1
c4Gisk5zg6lJ9zA3K46Bb5gPrePi5saBNwq9KjRU8tlAbLFGr2EWvjNrXlRlreJZ
PGoyu7mZFZEByWarDHkPyz2qhNETGs4AoCXnMpFiL63PD9VZYcWma2xIVm7guPhm
FYEXDkx6kpofPLeYFs+iV+e9hvvFd6J/k9S4QysXCDjGH+eh7wg3essCIEhweRjv
FX7hU8PTJasWY/KB1O3efg1AeVqaoaPQtAcfCMVUvnahde746dNw5Gwb6Xe4L15l
XAEvwwMLS9pFuDSWmuBFYvUMxrCYc4WNjxYhtxPnifj2J7/7uzMGGzgRoCG5MXUL
/ERZKkidpLkXmg17M4qH++sUh27XVmfFS/riRXG5Mn99ieuZB/AwnRCakEqsK6d8
CKth3QeYuDCR3dkOnRshO5JbaXpLVN0SX3puN93c1E0AtiXaJBeggfgvRravOEQe
SbZ+qwBHuqT2+Dgak/WHdIx9/PpvFJ6fIgeySnrF5hzQUVd9f4SVVof1iGy44GcY
I0TM9yqacuzdTVmFCOJo5y4AcIAuL1FQQLL2h5DLQUZRHN2U5BRXXjxe6h7peL+2
5caioY2cpsO3+/fuXDA3eaGWmJmGBGD7YiyufMw89/gsDYd8My7nhpYoo826TQ24
7pf3srvWkvrVAzkvHwEUeR8x6Dj0JF7WfwtwV3JMx0UaG9OMn0fHyvYbQK9lvuPA
m6XswNKWz+QoDj6gv2gbOO2caGynqygn9W9d3KD/W6ZxTP+1Dpmb9o6RgSGqBdEj
2PwYaugwuCOaAJjy1poKbFD8Z3MXJz4Bg91TGJ7ahj6Ws+X4XjZjc3C/D8imngaA
cMFcQKM89/LBWG+us3gS84n3e0NH7pLWPq9Hd4JdHkY7FBSvv0BeVNt/eznRJd0I
rA0YnCnyuB6D3BNFQRm9+wbFkuDrqWtnnMmTUdWEQ40RiyWx6/HVX2LwOedZiMB9
KpoYH6qClGoazyMGsIZ8kAKjBWTXaaQnymY5Y4xR9E7x7HhM6TxPUFRCF4JG3nSB
/WyHFygd0UKHFpRCmADaM+4FBm+/56VNhD1q4Iyi9FAQgHO9+4p0XYkkbjG3nl4/
6jQHp9h8hhTgGlWZ+1TuLc854TmfvhihY0Ws6fYv4jEzRb49om9x8Dnu+6jmWjGq
NivGkP0ly6NIVbShqAye4T4v+CT2BftAMlfoTDIHzECO+uFVuVabJkbX9oNTGkDg
2dUkw98LBJNbOG8XZhmrThshQzeU+Zf4ejTlocTrnTVaIW49DAfciPryvdv5JWny
NUuiU+r83Qd3mlIhHp18apzYApSYxsCRRJqLjvy20D4h/5OOg938wF6InYUzdhAL
a6GFvW5mwHivmZYMt2mSa5KfckGckRpbLREcJeuJuKT/aG/hz93gnOYZSbp+qs45
Xh0VHS6FWciv5dJu1ujuWMGPcdqx2MOdUfKjD2XlwBAP/9UWB24oW6QG1e0WoK+p
tcWFm2M+jyk1IrOdpjnQUj5ZbUEcJ3znWp4GyuLGRqsF+6JscIduBUiWZJUOoJW/
UAzIdF+sJTYOc6maas6B7gV/tM+ibIFKElumJT/CFlQsCfmmYXa3sTDcf6dERdZb
2cKTh37O/S7wUNl/xHNkhq7vDZc5206gA10Dx4b6L0wBv+0HjlzhRITnO0RUOPeX
+I7qJbFVDYUXkdS+z5/p/L1bO3e1mSHrMK01fIS3B4KZQNzDYeNW+NX7Uh9eZkYS
hTCbZHb2x79t0VEyoyIf+CRWnYzh33JuqD18cbzIZdR47DCM2tjeNBWNPZrhYOLk
9u7rOGw00n5OzhMWSO4leR8USEt6/RBvBi2XYz8fdFbH6sX8AMRw4Sec+a11mEMp
gcFnXUfk8oQyIRGtV6cKL7DDxF59G+xqNOZ7FsTMe3MYSwRPKNh5wzuW/1k+mLr6
Ou5oQ8d0DD5fXlDatti6mnr+StQPlzMg7YgZiT111MzBGekksD+STsqcsrU17NDR
jIzdTEjRi00mHEw1uVc695cD+tX+QXK0WPjMxvg0C5O14iN9Vm+J0RCySinqo3bt
ydB/wyZFv+aNH6NrqZtywuP4LK/VJmDJz16P986wJYGUPTQL1f7MDh/EOMBCYz+k
MhlS98V+iOqTttjPOy7GNYT5IfEhBmhlzLtt3PwunyZ0OqnPF/ptKIFZwdCG7SEn
4dE/PfosAKeUiUhJ7vDoOA1JXPcjix9pRbaZfg2Sor8IsKloYfh3+0SZy9YKQ2i8
F/8zXHGdYv5iSw7JTa0Y35XNdv35BDXazKyc4WyJZS8cPlsu9X/fl+/uYspFBvTY
GYs6XLvijLiAft29xq5DovpOaajgFzL48h5LJ7DcpAinJ1SboXUIn3+4N6ThnNvM
qklTRNPfRbQ+qtPjrVoWJXdiYJjEm+7Z60spIxlMqKebXV11M8zLyaNo9C5xRZ4X
zusVodnwN1YgtkL29koOJ3lMSFs8R4v3VHQaKNbrMyQkiP8IdOe4xg4g/Io5moNJ
OvSmf/pXispVjq14TKgoVofGYN/ufp0QSPActqlHS36k4JsgyFDtfjqo7A6ioGOi
Etp83vvgiyukf2NXsTKIHxWetdEEln5r6oGDaOADUqqW4ME2DM17ZqS9DHEOR3yT
7m04NV/W4/o4nGddG/4lDB4/B0oe8IFhdZ3XC9BT84jK3Ggzkl9PFbRhjxrIVOEV
izfgjQPpcFuvRDQYPVs6mHAsnyMw7n/XZMx2Wlbj/QAUC/tpyW8A+9rq7m3ZjHPG
Bv+KNgxI+SMUfj+Fpaqxnd+LdngHpVVT1Ax/Q9X3GeoAghuTy1qy/xbBjQp1GPm+
lYsMvoiPqFiDmTSnYzObSf6F4EcDndkhazapHGmV0K6Xpj/GkEgatvz0pCcqrP3r
rMP6iOim3TaPLMQI0GwPTGNArL212GdKxP5OCCaNuz5egdZFck4JgfkCDlN4eGrI
gemjp4d/C+9mOe9JX3E84oZfqcRIm9OpcCUNOF/ogrLC2CzOupCnCEUq7OIMyqr+
71kzr3KWJeL4WicAIx3/OujkdAABU4fQ4OwdPFF5oV01RqBu5tGj+hlsqtWp3Iz4
I6EitxeffJaRtzVi+VL9ecasZJ+6UIp6U0u4/K+J5zR8GChe76R2g2po3d1CHHIJ
fbIi4IJ1tWflctqrJjU+27l1OM9ffg1vEl9Bdi81f+ovaQghsuOyEkjti8GpyD8r
xz5Xcs3YqdqtuqFWUsU4xB/+CxMlT1DHxK57+g/2j6HwASiqZZAuHfp6/i6Zz51I
S6CxO6q9lZQs4rQM0ynaAOU0C8B+Zhn50ql0YeawnJO74L0N4mSb1v792L2zDJqW
uIqH3irCAFRmp8YCQxqQiI7vn7WZ8bakoST2Wy9RamNmxi1/Pp4Vn2vYECpCLFAo
1LQDSWdjleSsIixCV4crHvfoqxJ/Sx48VOplOkSfODgC9v124hGdO3S0JXmRUVEP
1l288p4SsCCzt3+2Wl0piVoufzG2PJgUsNWHDvHsTC6uLnPhDmCPfai9y756gJSp
Fa4cHKriQtfYHKzHedxQhvYw60GFtaRkOfwzamARMuoF20yXBpwT3EQmAT4Vhs81
wTX4sm+gex9RC9QBdE2Q8ciFJBV241F41ze3aJsGKTvT4kQMFtwxjS+X35rQS3hG
ZSk64HDY0gj9JIvQsVqNVNd1bemwL9B/58OssX3ARX6mmqH61IIsx8VXarj+DF1O
LxiMZ2TGm5CEKmX7E58sCON7mfdLfTi/GbtMTlul5ZucGzV9eW+2wIW8MaRqwxTz
J74F/az+J2ScsMwZZMOJMvc/WpK+utzG43rzYPhbp49LJd77HQ3iHMBu1RoxEU37
mcVg+0W7DKlf+2cVPr9G2un5+t/0oiCSEhVpyqYc8Lr9bq94FSabj6y84tXBtXme
WEe7rO8WnpTRppCM1UQzA5JC6r1Nk4GPW+/epKEyn0FDeBwdpHCubwo05vRLnouc
7usxX+eNbWbQ37Cb7ZUsHrYz6YkQK6eiCmN3uYSQ1TtqFJyHvw7D8Oy/OZkjbijw
vzrq0j+VDmOUYilmAwgAA5J0GIJgIKyptg3rbWAV17kJOFVgHYWlhPahyhqKLZsn
LkESA1blNBRhmGM2lBNJsB9zu64/BZ7J0bL7jhGdAhWEpWNXKnEYi+Xm3WhIijj/
5OrWwnxdEPXm9drEpGVNuoTRlHTR5Sq/KJOJmr3HvvMNlbbaLim+PGPtDezFkXoj
2HeKl04f+eZgt1vVebmaCgrDH338r4S89TXoJ60OfOluYT46L2jAAaKNK7attvj6
4c+qqcfRENBxM9cCP1ig5aaPrxZ6OV7l6P5K16FiXT5GdRXmIDVyT7csNGmLaAAG
AN4I8N9ymiZ0WbB9EZaC/UzdI+CX69imtdSRKfNmJ4qDKbc8N3WOll9kMvG0wPTR
DNHhtypriE7e3O+VpdNhLcGQY82TgSqWnaJZK8CyMfk0HbUKUpyL1BHDA0DkTxPt
AfvhslkJmnMBhfPfT34FeWk34ZxFzIz7MVbEzMPsU23uXdiSFfnkP6nvG6IBVO4W
yRJLTdeCACCfod72tUAG5IVAV+KWbgY92ehuGSRZ3UinUXPkuGivHAba4B7t6reW
TRm4x/efkR8M26bUtFkIVSqcVdd3A41s5NADcWmcMgDzcrpzpbTKHQBTmlKC9ioY
nD2qvDExie3FL25Mc9Ke8F30KS0ENjYEewG8th+HJNQK4Uheqg3FwJ3AiVR7zNKO
jitlPXtqs9KFqm/tFn5qY8siOg2GTHLri8psophGKzW8ypKg25KNJFsJPUt0qhwz
HafvwEHI6aSkVjA+hCD0xi+KI+IyskBQgY5XPHgIEujwpQU1fAPI/skxXrjNLxkW
3DFxurhUuywrOFTVX51JcoIPGsWkl4H4XzZfUulCU75uB8L3WymVfMoH6UZbGCzY
LAYOzPcYCE87dGANVEloKoC/mS20JrRzvO5vRfaPwRSpZzbjyQXfPtJM3odv542M
ET97M2yVrE5hnMy6DpZemVJd7LZsfJLLWEMdJm34UtC9vXzP/gVXZ4tTY1ybCEWK
Az1zAruCVAmGG0/7eSBzN6nkFFUdOV4mFdYmei2PEUPs0Mq995aG/k7aCgXNJBKt
uoPBZQ+Ombl9VKpXJbk8/lLs3x/hhRV7vKFiYfsNGHLy+NcjAvVGEHHwblfSfhZ4
O7lzNyq5drQ+VEW6P27dL2MZ3sz2+0FG2iJbhwiPKtF9fKE//f8QoqTg7TwSAuEg
hcth8UFB8+oKT093uJRV8XVxB4GK78fWGY+Vk5gNmAX5vputcIIVIWZIqbn2kF+f
VX9ZSVuhY53w96xnyF/PDpY7F+mf3/F0VbvJAArZHZ9/UHiUwrmC5frzV6Y6/ZAj
SgbDu3HLAX7S6r+WobbtCDwHgcl9UNz7wslRYcIzFZVsExaBLSnm72b85KBDMmcs
1UFH22zehuFsbcHpJNwbplPs3VZhisMiT3GDNCytiEMnHqMwf1Otawk1JJfBgO3f
L8bdCVooDvT0C8fn6u9QOTbtO23+2Gi3eBKB8uHGT+x3RF/u8ZG3LsknPfexJtPW
XrPSqDirCLCsveNkQfsPtXKMOP/6SzritVW4yoCYHp2HddgoKsuMWFsCugWauLjI
3ZYZ0Rlv+O/I70BB+k3Q7eC82ThHOySmOcO9azKw4oJZ0CUjoIRrofCEMaBsmdKv
vfOZqXTbK1dPSZ3yYlFd6RKRXEMSwqYFuChczpH59DZJTzZZF9drmS32xv/n2tQk
esjw9cMYx4Lhra+DwevFr0uwcY8Np7ieAXp9Foe94AA5KZsdX3tXl1JLEHSpgMs5
wwuCHOiZ6Qwe6JA3LIolArq3jELGyKRpAzuW8CBYc/8yY/Y7J2nm2/9db+af/UnK
Xr79i4/xKqr1FaEjw51CfKvNRaaX64ObKDWQmMnE2QoxAfeflC1wHEsSTa1RMMv1
yO2qIaAWbYWBKjKeCxMjVF3W6C5H3B4BYdFwSgzoG9OJYTzWh6B9kphlBrGiyI2C
RUDy4pP0LCnsaFEvQhd5CLqFeuP9L/T7u0l2XULm+z255El5mtVznJCDJiKzZr/c
W1TMS2d78gGUd1lYcHlT3Ay21ilZHDPOTuiRVCWrrPlgT3oUdGzN1qa5NwM4084/
EbOIOPnDhhfhfSuBU74H6iYpK+8bYG5SXcuwSDbxm+Y5hkp7TXxM7mLfobVilIqZ
cM+jPqW0VHoPKHPZF8Np3q14BPULnG/Qs6pk8KkNEOfNqu6qYLUP2PbqmXbJuBzZ
jQT7Jv2fHSv0XkowS4prpwpHnJbnpov965ryS2GnJYHDSNV5FN57MD4bkMjADpYb
vP1Fer99Ekebrrd96aEZZ9ts/mqj7TOk8GzF5YCDP+hL8RkSu+FC4ZofgX3//Lf5
r45as+zAvFh/6ceniBp3CY8tyZkm0929b/zGXYdQ6hRWihZn8KwkgdE/2cBKtIu4
DVsUKqA3n09NTMwMgddVuKo5PaSZNHjgs/MhAM39Lq3iO2d8JOMkV9X0mi0OrhpQ
NpbSpq5I9XUoP5UQD+++YMTq+opu3qZD6Ie5tHN37cN7wiFIZUwCg7kehoH4BKNP
ZMqYtUQej5WuHljGyjQDGp0JbHpUDABVLWK/OWCG4CBjydsIBP+DTLj405S5Zbc1
KBGm5giOOIFv4jYCDTAaq7kaf1TJcuGRWNRDQq5MZ0p9t5VWzLr6MI6ZlpFmQKH9
lkOyUTbBFVff5E5ZHPbG43A0ypJpfVlpfD7jOQBylq1yQcR8LDExxpQQJVTt7yj/
EJ3JA7Jw/IYpWwXUtOAA0t9ELuch3d5Pp+qae3TGc3jANn/7L2exfjtEeWJW8frC
ItmGOg3vyjFygY24DBxnqBDCBCWyZT9rA+ocPmo6sYQ/Lw7PtvdkeoG6Lk7gjdIA
v8ZLfbRjMHe2/6+PzzWnMYbMBKOIngFd482SWwDI/Mjp/sjUZ4KCUqtcZNRHDH9z
H8aQCb4Uxt7uZqA/YAqLFsB6XtQpcyJCcqstWiNnQRfL9znfLbG0ey0sLkhNGJvN
EozHUQZ3Gzy3SnMgZF5WMDfSpn5A1o4VRtco1QFnQ6Tj+vcDFwGXyJTxfUWIWKeP
rIj9EF2PfVZaJTFFFTWOt/0ualF2zJXtX2SFXN4ooOusdt8aeMwbZrF2xrbnv5Gv
eM8egTSR5sVgt14TVf1CSHbCVftSlg4U44tjiujBKJdzGlQfgPswBjzhdj1AeEDi
r7TYrS9R8juoaWaPrbq3wKlE1hfgvMPAyxqYNaavRAzfWpTjVyQ295RbxA+z2SZa
MTFoXYJ9uYSaao0jzjzjE7FtJ9vLWfGk7sWV2p0ZF5AR3mu9/SfzOGK9Kh+IvBuU
7dI+CORYcIXa1d7s9poeFvr0npRmHKTQmbMB64ASVauUOje6tL7pqGIQswBz+Ysm
YySAyliC9RsHBBcFw/gIJnkCNhkdBKJ/WK70hTPTLBcsm7cFfC1uyibhKZZvdoJz
dCm3KodvnC04tKAzJ6kp+dfvi8W0jOT35/bq7tnSVxx4+/jXIgESqZBGPSpFuYik
u3dIhQNwjE2k24zeawQNAMhI8cKO8BwPxNVzxJtYKHFElHgUcUU664rS3JU7ooKX
0XLmV2bZbO17Tiy/CXMCGVim1IXkX8gEF9ttyM0gWLBDkKQvhRARtWLuP2SDuMkz
inYmJB3Q9mW0hisu0lFlgKleooy/CnfHHomCCCfRqMUpUccVWcjkOn6ZaGwoSzl5
VyMXUgysNu2nmL16JaiLvujBWq3Uwfe22EXz998LLSVvjwGqAPTTtNjww4HixM/j
rjmO8SO3+H62t0ehaGQqVKIkDLYA08LnRn+AYUDXfhW7DSDv/z6YeiEQNKVgM/HU
Kqis+s5QLj1thhV+tWffq8AnOelIF3dXa0+KLtg+9OaKPorPt+48NFKSVMXgZ9/Y
ciRxeXFGszP64tuz1SVNJ4PZro55fo/50aitdblQ9IL9t/VIsGl0oCRnQxSzpGRH
coSM7SCHpY2lnhj0Nmff09mOIAWc3Jh9PLWr4RIzfGr9GZeoO9KMFXWmrneGdjOO
6OMWFUdRvq3fLo9sJwecLaz+pTLxfku+APXVz6U4LbDZHgB97aJdBk2kjlqy89Yy
AJagxmK5sLMDXnP6K2UwGxeLDpptZcqiwpT2cy8T5K+JOSLkJo5z3IEbm2WlfXvR
GbK4jVk1qqfvH87VsyF4fssSaZtkLGRpcAN4Ig97XNma5odTus3wF+c6jWp9ROuz
aXhlobjs+EnD6VCfUErylzFpihIxGPaCWNE2o6kuPJgyolalO4S3527FXhyLr2Rx
C/3AK1V18g8nGFvGDlMj6rIs3t3MkNzSgJU3X4BIStii5UhAcIv8SBVs2MukyCmq
EH+078s9l6uHOkXr1Pm/4iPhkyV+9CnqYM0bZ+CXlxU9mLWVoeW9SSoHDsB6SWy4
BokIl0tYTsNRkT7p83iK/MVRSAps0Je+TB39EsJb5aPFKsTgUQ7omN1rqUEDJsr4
JvwY4Tv0JWIRxbaUElTGHWDEizs85KcG+Qba+ndPla2SaF24sbYqimIpAFuGfYGW
dd5+4YvIioohRL7N1z8/+HKMUq4F0HlhlDteAVP/2jwsnz1Jdq58hsbHBRTRJeU2
XupZo+KWrK6VqXnR7b7nx+Pm/pSAalNOc4Am6dvuDHpfxRarwT405364ogfzGEPw
ptULTn6HFAdIY20XOyWUHupznwwA14mTwftCW6xThJlKg3Zacms/8MxMG5eshmzw
KU/XJJaZtJN5OLWH3JtZiE7HNin6owG9YOxGFxT+FgFlkMPJVeFAnU9nsgrg8cg3
BrZ8vEavmzRQPbSgwxbC3RifrSIw3BWLcdMTIHcUXUPrP0gF21NQ2NWwrqmQnblJ
Jj1Heo5LY84RzYLkgpD29vMvAm32chuvGtUdqwUpQ5DqYVgW3atBs7bV3OpRUKRj
`pragma protect end_protected
