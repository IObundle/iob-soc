// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:39:48 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KL6TgjwBX7R/9z6Lrpn7kq8NlBhPu81JPNcMwN+b+/7cKH+8JSkS+N991fOLrEdo
F3ugjph0fUF7dxK2xym+/DXfxotUAw7mjkEXDq6ANL1BenST6Pt51IRP0clrW97u
Q0PZ0MvHpBILYUmDP56WtTaiop0Kp0Llr6IjoYqO1WQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25104)
wgY5jD79o6RsWeLDRVzx4f9yBeZTXywbhW6CGWSGMbVqFXYHckDaPK8kLRvnNU+e
CBV5GJMEwyWC8Uget7MwdXRTHRaslWz54bDAaVLRYlrKys+2pDes1NR0x0A6VlPc
LLoNzX+aHnB86esL6vtOYmBn1qAMJ/L0hMKFLYf6CBZqekuWVvFnt0Lun9TpcVxA
z43oX/NsH4lRzMe5fEgsQ8UgkEO5MOpVNCuw9doYO8ldPzQLB1QvgQAduMUVqOwe
08/lfSJxVIey7kVoFEhrWPFz05OJQ5HKFNlqTNJvyx7xPJH8HpbQWk56IrgUKh2l
gkloD7KgG4+DlMMHiStpa39sc1vTYFxSReK7ZNXftwMBwrz+U3pURmPfqE5HM9WX
uJAQxX69AzgqVyCC7LGHGWZ7upR8fJxeanoKAL6Cj0OTaw+ljaw40KQbInHdJwMT
DdkMBvwFwf8MaG+1i7IVEZqum2cc7atDyc4OmS5K9hkSOM33tj7WjZprmBrF55ZT
mGvHSmsHq1Puyirh7/6U1WwEAQG7T2M54Oac/f9vR4OJ78KAYVN9V+75FjgyEe+b
aaGa8pRhKlz4RoBk5zbplfVvkPZgJ0rUqaBX57x91kDu62qdBrjKAMsGDpvrJP/2
RKxyE5YRGghv/PitbWu+O/Iwy+x1DOzd2zMB0QSaVxbWfMGNo7yd4Ba39pxJ6gYs
JiyucJesZiSmwrvkA7K0ilKUhI0kE2IQjpO8zAki2Dlolxumz4uzrKG8Ioj093RZ
m1n1ZuWxkQ71d3biyWmN9cilI4cJEL6vF0iiC6ih2YWETc5MzXB5pMA2qscaEd1d
gGEzIuM+nDfaca12MidxVs+WxTplru4/At79pKeNUbmcsavbruC86Z4uzJWwGy3M
RWkTcFRH3n/GGUdvStjbwpYENSDItVZgPQNI3WsmqlHvSXzxp5BAX8oxF9eP6cHp
Sbg0zu1N5V2ta6Jvruadxdnh3OMj6HeJsU1N+JUCaVPe6f/6wqpiihYcKbyu5ofZ
sElE5vf/n6cxUAhPhbyzFKtTZlkkT3chN8gOeP76f3DZX7tqsMk1WbXWzQ3Fg2p7
fI6L0V3DG2vGc/pwnGznbNwCvcamjm6FXCOktaDQP0gvOpiEHyFN6HbamTQ+yEIw
Kh1vvF6YDmDsc8IsIH/2YuqqG7fgwSnz2UjcpCU4bOijQFT+MgUjVL0waRc9bk6B
WS3cSEPu3nQiHo5kH83OW+Xo0rWjfpOIYeZLezr751/Y62swXD9V0Q31KO++6Ku1
Bjngodr1NOatIhbIEshsK7Z+IiOF+1WQW7Rm1feakFrKlo+j0gS+9WSliFnoznls
SVw7iDShFRjBALS5E98+UQw9nH2w55AHtAhh1JqBOBmDhguCWSkqm+fxKP3xLFH4
lUbBE4swwwkD0tooAG23zmANhwuaFLwfZaHHhM9D/cf3TchLGxGDW/UVk3Vyq1+G
jdX1e/4/smUkjjG0srsIrnZ2B9hIK0T+m7CE86epdiBFotBdIfuShCWSoyNj/ZRq
Ny7IKzgyUZwGTkJ08nd4BNf4IDbSHZX+US0ogNWe+jVuiM0IcImEppTz+++UL+4w
htUkp0FnDtpi1Rrdhj0MLe/+HCD8Ne0jEmxOMvOOcA4dTDBl/QrTUxt2+oLiWCb2
TvLqisX1LeqasfcLtBAizZ14BZ0u1+aISdDenAisdhS5eRtmhoPIQgA6l98VUd1A
gMPKtrf9EG1TCBCrqQ+G0FkzW0MmyWmDmQbUCL5erU0+j7EpwQ8FGrGWCZ+Qdixc
Bgn1EHq02XgFdqlf2iQWzSSENcKrOePWCnmcJXGJZ2tV+eLUQKkKWCaMEE9l8mHI
Zjej0dY4/zonjMsXqnHfcp01FrHGuEPahkI/zR/zpQPXCpWKWps0X800n44uLP3K
eoU5z5PjJL6wuVRPTxJK4hAmQupjB0WMtKc2uZ6pT2uM4WchbAOPInVdY/jhCDUC
4vNJFCMjNMjZ7j47FaxQmd7V/CNY0GZVi4nqHDQEAJmHGXEJLSqUHhtv/lnZD2eP
+VP63N8nFGMsvtsRvyamtrQScZjxxu3SxpFQS6Hbzfdn0GJbEOHOFFZwkH7ep2Qz
PAAcNGSugEkAeuoVjLEzBTNBf9EEU+pRRmKmCV3pfUMbQnddnmrU1/Jhb2P7ZK0d
WeH2rLP+4/GKqX3dXQ9IHiEY9s6DhBIjM6gCbG+P/HX31F0ZA6REurk3F7+WAQmo
mfZhEw6kGqKqIc46WPVPiNSIx5Cd1QXnnUet9LL983EsqivBsUwsbfuawdDxp3hs
Ws785LOlCOV3n/dEHxy2vmsy8bQnnJ+FZ4WN3epmX3H1yIuXPojyMHskwd1ZwYAL
FvoiemtfElTwEOJXToLEosZ/VCUNNlueKrZX81Q+DIcopL3FcyyraZeiVsOq2DSs
USzuo9AMjM0GSzjdIPlaD+neKSD/LoYZ8/0TOKd0YVaM4XrK+3ixFu3G8B/0ZB1u
RSrGX28DbVkGWujk41157Qt7p2ROYDmJFzNLUU+Dv5jQ2XUfK8dtja4oW15cpCfq
Lcx9vJs548NwHYZQn1i0rQvkNNnlW+Qk4rn0DqrHJ/7ulrmAnqP1S+Cb6MTkbh/M
FvAUuLvatIFjqE9tNUcUZPkrL01n21pV2RI93qFR4d+Hvhhzc0GG9uEisdeQG5a8
/aErYYKurL+Emd/2dHG47LmU9NAxboTV/E1CFy0Kem1MRpTpdt2RXltqH8isKdWs
pK+VvpmXq25rxAZq6FVSO8vmvI2pEYI/QOMsXHlha0yPPaXu9HI+pDJazplxsvsI
oqZV16I2KmgnKJKbhEsaJA26C4FLm9UBe/JiOaaMv8AsqzKPCSxK3J/RU5nsX3QZ
KJoE6UkCT0uUsxK47uDNf5DOSETALkkSPoXdjWvIIsWfJW2Cz974b0Jfj6yxIOm2
U5+5fl1i/LHZu5I+EzuwliUmsHDNym3NOhCKN0ZESGK33VqZwmn0kyTBmjURq5xV
MbKWlCcAS57wI5CkaTnww21ja/dLQ8JJOz7+rYtSS4GWHfPaWeqWa8tsNAdpMBmu
pdpKkFbPbAkLFJw4M/JuaLEZuwxSzFMEzPQzjm1/fG1zHLdZueB3RlQTqYC2Zzgv
CTJDx9dX2yvSzyj2rmNLoP/3Wa18nTUR3J0CSDsyUDL376wtbiKNU80GfI0iXYZE
gfVIRhhbN4HP5AkcNr4XDeG3jEzsoJuHiJC0j4wTPi0rYUsxNPdoy+p7KBGbvZaS
AQRhNEw0KceouNPxnt7QbKQKdoC5PtjSIGMcfaOMHDueyVAsS1KON3d9a7+ERggF
1gXxiGaDB5jmLGRHvEDsYLMqU89aZbe4U+xT8zOSEkid2w2yerN57KPBO+5SxNfM
rlr/tmOQ5B87fgvSlgfzK0Pqo9IvXHNIAhJvJWD03AUcCQHL9VFlnzoRRnWtL7wj
RbstfkuDepcY8W1R9oAbfOp8p56unr4+0XnB+L1UHK2parWUEjzIsWyOBsvtA0pv
jBgY5XvgPG1QUEzDsRGV5lJOteOtYVCsvzvKstXT5+TjAsGkxUQ0b6Zzv+FoCfdg
f1AN7XWjU74T9wmAm8sSWiOktSeKW9CSKRQ9MpjFnpNO0gQIjKGSRMHjiPMvmEw/
dJNwUZdC9HQcHmATBnVGyw9aBefYFne+wQsLlXe9hYfRBP4yARJeXSG1RUkaY1PW
cCVuNXJFDkJCU8AgeXeo/3sJNzCndh/Cz2ItoQRrxp8StoEfXSI53D1M2tx6PX0+
SpZbVX00Re28TaoTVQHai39QXZsospxbwmm+y18MTtwhknQwATc8jWkW1526NG5R
/gm0tnx4H6QAWHntmNz1r5mw0FE5I02KKM3WCCCJqEvYwzkuLrCt8AcyF7lxxGXt
QnuP3SWGCmkU89Z33yBXcDBRY6pFR+cYy5G9V1EVn1wp/Xb47hKx+kJYhc7sn+iy
m6oLiHb9T+I9H4+AAnlkzKBiD8mneLmhAX1HuOrdyCY8ZkTznSyt7FCPR80tY+bU
n1O+co2bBFW3wdZaXcUq33U/pT2FHlhxY0H9SL+ism1gzNJYHOxW6muBkoSd8Z8F
ieGz6NqnempfDaCgu8u0KcDAkMBlylUObDkFvxWkNk5lb2BkEpu1k4t5Ow785MuR
0MmJ8kOF+Xpb6jYwJBcqjgoDqi7xqBM9hrwQiIiygDdC9BmeZVgo53t51geRS06H
pimWRMqmngtO0fjY3zcs6Hhi0hoM0xp1RoIqEn0MxPCd+jl8uY8Hm//8UE+H2YDq
RBwGarsS+oUqUurPCbqsuHr2Us3OY4Ia586k+YuWWOxzBpfpo6BnebG32o00XeIO
u4kQ2/vjtUS7NhbAcRbxeWfASU+JVq2mxbct3NEqq7X1fg8VhqVNfAn/vW7Z+SBI
KSNGxUfAlYgyXYxTIFgrYiX5vMKM3hJjqj6q8s/p/evmRE6scEJL3Q6VVL1KRy0k
MB1FPUyt4EZFten2ukLd2UETjcU7L+OjVQQqqYNOFYoShQYTj3cgnqQfh7F7oQ7i
Ve3dvtniLbQSUkW16HPTxffsk1DfJ5rAStxjNKfvXBBXNAeEsarv7jcCO+GP4rQs
Ls6GOCYbbM/ZqBvmg1BN+77hhQcXjInQgtgRNcIjmcqcAmcqE9iBdzAlIOLOIaAO
lxXShrWgNxQ4r7f1saAEY1mA4Nooln3AjtZ5dyYv8iYDxJWYk/CL3+qPc+hJIevW
pAVG2WKygcaTJgDRvsJeGWX8w8vx3D4pkUnD4vp76iT+6ODxMuSGd3Ixqo1nw/dG
8AsFBntjDx4aMpr7kmqlBjRJIiWtxThFeV7ICHJrUzX9qlS4WrCFy/wb9U7sqiJj
BCGfaR03yWNO+A79Kr2Lk4o8mr1QymS9JP4hyWwtVDqimMhFrrWLWU7BvnesspiV
CKty1FROrxwsQCuF/YitKPubvn26H0EIqgiEKkAETdj2RFWC3TEEvtOqifFl85hf
QwYBpmVZHO4VXQk/uvvU317Udr6jviDLzC9C8tDsgyM1urw1pbsHjZ1sluqyza0l
KsLp2UFXAaylOZq5wRvM+oXaCG6lkSw3eUDaRbCOms943QMcQrUxHHK1Y06v/4bb
HyPX+I9WdIBK7Ypm//eP3/8bNgsNykMVOob3ncrSU11E0s3qKTne0h/YwEdK1Fbh
4CIb1x8LtKaDHJGo4CpmBZ8dcXPd2x1yMNT1sdbdBPvdgvsOg0uUsBiG80QHOdvC
IrttwAWJ0vQKxgedl1FIhcjHQ5oUjbko3q4jmQhhu8DLhcOSGKCFReASSYTc1Ye5
zTdYHh6/9JIS550P8eek3Albwyd+XttxA3DDPr04SiVpiKM99IGvna1qQeaibtoS
wlJrK7Ary2OoAnMH3nDXp6rbXvPmPO5icuRyK4w82r8nZ7sAUlOPLWSSi9Q48RbF
Wx+C647nRrDQ6py0HWu8jtAmbMsgFNvA75zwP4f7jRXaYKv0Es/wozQaURb0i/Wx
/N7U7l2ddL3bKHlLx3iuBc1fqju3dPF9b+HRmxV0dWojSr+eINXQcPweWwVsUxYK
XGTVfwYaFvYM9/kd8fm8lZtRJeYuZxpJssc2oCqZuCfb19TpxNxvY7ysLlSIMvqt
jStB88n+/C666Ly0lz+vYiCg9fBrez1EJft3XbMcZW320OaIfex7nsQzOVXCQS4b
JAl+EIZzAWPrTj/XuHx/k/dOYCF+uzq2bEioDXOmjFFXE2DC+Y4rmydxOrv0/CsJ
Eu1rGQaPPxpj6tPBK+N/aq/TW2hFGmWuJ7jLM+xhKUz+SE7RbpwGsgp49p9gSlFd
LfVXV6zUqLSTDamLjctlxdPuvcApYCEJ0+ibw1TISMdMvYqhIT1/SnWbpSx5L/Gc
ZeBJYA7zm/474HKtTc6FnYQ//HP282IJ7TMxiq6zewEGFBj5J7U7Ql1cmwyGlemM
QDRkyiZGo48WkwA21n1EWBTF+tyjx+M7ucio0qLvSl9GKs18k3i6GnnUQ/SuQvYn
nUNpxUdo4QSvGpmgTeBRFq9AIxXjooHbX/QQL/TXWuW6WTQzUz3PjqJ1kbrCuuqg
zoVX7l9Di/LmOGxa4G7UJ7mQuWzPA2clCNIfnqXNiZbz9uqLTDaSJCL+iWak+b9a
Z/BmIUfkYM/iMO+OheTIWTxNV0Ag8mWwZMtNZffsVgUhuJyNEwGsDjTUj/ciOwrr
6LzNt7KgAq9GLZSAO8gu+Y4986z7xbE/qUBYPoWmB/+bx3gdh7BJqQ0zUFtyjQV6
Agoi3d9YwecnnynQ9XxXA8IXfvZS8pqDCem/8/RrZkLMNZ6D+3mAcpnhET+F3NJu
dHOvttcyB79kMuuI/djTWJyBnr79EQNeFpPAa/LFed8HPoYMje7zlxPGCez2iU9n
EHp3tSXYGaRGsXx1RgwR9U2T4gc0rHwED8df6rbkK8fRWuoI454/0jvQJKbNzJtP
+daEHaC7yYMWitO6TRS0RLx5hwg7L8YpaJqMMWsBbxHJPem0po69tC4TOrE0D1Cd
yClITcoAUn2WEMwQyF2XgIzSSq7FbdyksxViiifkuxUTOh6zJgQHr8iVVIQZ7iPQ
0R8UvZplmX8wnADmneWLobUoMEidmih5TzeorPzVJHBDgF27UHgL8eu1SKo1ZSkR
va2OOFcrWEWa2J+aojvmlAbW41Xl0BTuWFWrIgMfXYMy5VGLV9l8o3TibDMIlVUA
d93Xh8meW/+5uTiEajeId8Ht9Srj9wQDwH9GG8KqaGAA8WCe27/02JMvYOCQP53p
S3RLrBB9MivW+nPE4Og7cy6wPm77eCaLAvuyKuZJRU3pbTJCOBqTIbhb8d5WpMAw
+2yx7LudGUfiddXFHepAXr2+Rop1EuisTt0nuT6uCGPshyCVvA0rBDYeyNBCUS7A
ib9v1WRNhpTvbZhSm4SiSrzxRgoELXCALpQs0Jeq+EBWp1sbI27R9wWyYtORiE97
+7EPX21hMxK3Aq2VIyPcXfL/lnWr9b8YDxYNjVQiPimbhX/4Z+NbAXSfrRTesFCb
7lYHpz0fOeYXUh3P5CCVDlpwRCiKuJyIXpOpDnYWD6TLTbWjtRgW/6HpN3sVDYeE
xCSD2FVi8UJjpbKFoJ6AKTI6H6r+/y1oliIeh4JINKuOD6biC5YIgX72np+3NgR8
u29AL9QyFNVEYNg2oD1PScJ8ijHbMzZ5j5lf98Z/sl3VBZJS0pwlT22zV3Nnoncb
H6rCz+lA7yO2BFHYdSayC2C7TUEokOs5dohtYDdrmbgELPCFW7bbyz97HvPCn4hI
mATsikG6163pPWiohOEW0qYedmqF9IUcTW3LY33/57XNFf8Q9LMEXTIxgB03tZFA
84wS2F4NcKyaLvic05MyzFX3KL1xCg2gqmA0/rR1unyIE94oJR/yTGYQMFJp/FQ8
oR7uSBKoaKTBw0p628hYSrSHOuLf2ekjP1EF6/87SGKc63kmD21nqQvAjJRgv7IC
VGNFijhmKJuIopcOISeA4Y/PVghtZYGQTnKb9V2pqZp0jh2P9Z/3YpzkD1k7HO2H
gRl7wQQ/1IS9rMx+CCAIJzoqgVoc/d0f0PKtbLtnlgTzs3zcDwAlBK6SL+edEbpp
4oEuSu/w+5UGOtEt+bNxjzSzMGTrmWf7E/2N6Nx095Tdglbpc10QqB5L5naW6V65
V3+XS6b/WBHFM0+KRWmhetgp8FVy+CVyYHQlV5oTtWyxom3KBfvCjwayhX6tufoq
XKTDSSTSwjTyn2yYlaygEMaJxfiWpcoyqLTiY8hy9AJMN3s0XN8I86ikkCdgr7d4
AASixIQUvyWIPzbDvyYGeRgCHitsgPbE55cUZ4R1IRTYabepIO76/JmPFWmDR2NS
Ee+S2RtVuBoCGOQ4kIcnESn+v0w4fDL5MKQEHATyTNNUO9b5TiRm09o39QwNRf1V
sEABvZeGEcgJeVs91AGlf1BP34bmwL7/JewPBo33a0+eSJ0/+i8Ro85a4YBq/g8Y
R6PwEW0tPdLNmRrQkuTwjwxCMpF7NRn5s0AB4vJUF+SxXx8KaplniRFfK+163oIN
NKXixtT3MSu5WmiVJwpBfWo1pocd0DUw2Q6ELYmH/UxwgixVoaJ3+0Uz4S94i1aN
gwJvUOBoyYIszEc/gVbdYxVqyW77+YlGUIMe1GTeMNN5U2gk82C319xeuExBYKDi
E2zD8x+GcpuhgtS8pAmwz6nVg1C9aY/397cayuWuCLSCYpEoK0uIOuqmecvZNFGP
s2y8T1K3gOgbI3iAydXlNH4q+I1TD8LtjIM3mKnXXRmS58vXF1oP260bJB4UZhjO
mGZfRhYKl2byeOPoKwhrkXI6EV2cBf7J8jEb3VcJk55No22YbRbOs6dSL0tYpFFd
GRfe8CIqqb17SZWoje+xrMHiUS2bzw9qARGuKETb0fkcIdT9IqqNTAQm14dFEmDL
aIUMH4M4gywfIzYvF4Lels4tHq5odj+jayOv87pfd1T64ytLUkA3OTi6vXlGUw57
3ks/dm2xB16njC6o70kCmZTyBzj+UUMRqoehkwpcUIFDs5g4KfNc5WuVWdUNikra
lSxaiKR9cjt9AtuYwj7QKTQB8aN30BOTGaIkICMAi/N85/0cgRrp3NWsRtKJ/woO
a11fVDR7O39Q6rEsl/9Jw7VC1w+VwcuyWiwVqOHlKLOBdDrugDsAPwBtduA42aYN
xP+8Gwwa01kQz+vfZdVnaeCl1FzmeKrojT6DlyP7Rp3EKRbajRAMOHfOn+X9BY3k
TpCPlTmneM60sYQeRsBEJO0QG0XtyWw+J0kZMdmujlNoTRtH5vLWRa/0/GV13OaZ
8KAwz5Zl6XocawZA7rgZh0F4/D7bfm6uL0ot3pItSJRPwCsRP3UgZGEeNsbjKb2y
WFzV6/GGbNgK5diztLJoUTu2rMVqe+NAmnEWXl+6frTK9y6rrDO0C+h45Fwb7vM5
25Psw7sWKfooVmJAyr8tMDF/M0GPszilmgRQLH7XE0q55TWzMrZiZTps3FTsVXMk
iWyN6Od/YqefBzIsJr1Qjq0JGXlMHmRHeA9w3a/yFJt8Z7I4ryVpyZ0kwhKmdEsk
Qem5xhkDIrFAJ2dIbxGsxr6tCApjipF9XX1F6QbQ6B/U3oNRYYajFsDod7Grf9NJ
36z+EqWbgBOVrxRpH5jIwHlQzmJ4bI9s5eaS9QV8gQgzfVhBxdsh7UvJ1Zjw5FPg
QFMoZXT67kLlFlT/GGzWd2CjmECEz05VWNlhDLDXdFqS+4E4EWC+N82RHIHDru0P
pD6YcoRDnqCDzdJCHO0t18OfsYRsQHqAn+PvU30M9Arbls4COYTcO3RkqdolOLg/
9edYN7VAghyNDFqj6T55K4GwcavVh6+6U3njNHIirlO1x3qU1ytKutcN8NS853i9
SfYuYQ2cxC7VtlOqSJ8GmSVmSrzoyY9QLXo6onOjh50Hcm57hdr8QWUW92sZjgwI
tqp0ZaNiREHBnissEQZegV+RWUJApPMiNnkvmIxLG7LLkv3KMNNEeavG29dr3NJp
dniTvRJhubIO5Qc8t/x8RkQLAUZv4QcpH8HEEFmYWXrWK4oS7zGYqGlVhdqubUHL
8XxCaYhKavYVx3b9F6NeSNtKWmt7ap5sd6qGRNno4tV8itA3U1I4lMiIm0oNo1Jr
RSefIKnGkHVPTyuUtuyMRlyZyJBncrW2xzB9HgV+fMFv19ZTWkoVypGd7XNPQx0v
DhE+BUuYuL1PpKVcm0moSOQcvxbcoYJ7N791z4Ynk/U/HiScJsSWyDEs7Ji9tqYS
yc3x0rNgg8/Ma65p1FsUKj9tRWj4DbVrG1/jZJXuJB/uerxAJOs2uz0//DVpD1sE
4n+4NNWvXf95BOQdCe2LngR7KovRp/3chsRlIqWZTpJrSPofInGl5ABEhDSCAGuP
ED/bNQmj2O4PQ27weslE0N7hE4j340uLxuSynK2M5AkJqs+ZkFq+jihmZ3P+8nE/
9Jjmc7lQ/IcfnKOs3vhE6r8a6Y/ABwXoqyhjUueB5krRuTkVrSqovgsBcUYAoWc9
44urr5ZLNEtjyNNgSqfCxgCYq1qtrvZxdI98VIMPqOKDqsxuo8ZRGzFM0FMhZpa1
u95zxmq34UTw+mUyHfj9QJgIYny6IlgoMv2csFGJNJgtxBguuiQd9omC/lEFs4OH
nxfCe/JvMnixmEJTBO60Ah2TYMuB/x2TSRyZIq0cMRGCwbyETnXlZsT0WXn4MUeS
vyhmGBd7XU2K7pFt1ts31H/bSR2zsL65CXjDvgr+fwOYDqlqjuc2ANJGMW2Z45fK
/G5CtlZjQ/NavA7MQudBAK1NmDp2TniJGQDa9dndHtP9SEHqpvswSYSHz6HkBWLz
iHUByvaJDTznNKUCJmyOn1qF43D5Ie7Ip7S3Vm6Ljo2axCa6JQKyh96utl/a4gLS
P4fEhW0rW/bCinaY9PVIWZrUIsOGfrOMkTGzVGexGaJMcAYowuUTbMbNBet3EN/o
IEtnz9h626L/TP2Ok0a2E05A6dzObaHbZJlB42PCLdLxQaf1hk4ssIIPW6W1Av43
kdnlf4SsIr3YxcloZRjcDonRm/4jOrFrHMLNT5zantZPD38vf+e9zmz6yOpYmmiq
dTZNcUP1iN629PIhES+WSn8wYg9wBc6Bo4xAI8qM2RuVNRlkRqnIsc11draix1LU
YSRfZJs9HSyxTLH+Mt/KDUCUiqFPFPoOlIFUVQFT/d4Hbkqk5J3mW4tFAi83H+tq
RS6FD607CPAcf7PejaNUHQ/PNzNZRGKY/IXGdY7CotR5aq1YISiAdPcnUX4QCj4S
UH/fOZFGwJFYEhieHQxSPuElWFQuSBXzRWmvax8Piz5w9tPgwr/MZPzjl9YFq+jS
sCXup7PBtUmn9ZTkxeBcmF06OAqm+b9NDwuZkfElizeB1Z+X8vOnTta+OGmxwTW0
auGjRSve4dwEVIpZ9l4vBZLzyUaGsAZu4i5s75wmjk9k4M7VyvwySBqMvGBhKpf5
qSHgmJGcelZFeyThCuWIK13DcBN0+AL9egYWQSLOCrhF/Qq74/0x2mvHn/2bbzII
riV6wna72OXmje7BQ4plc+sAD0A2WczE/aGLqEnWKUczYgSxFj37MQ7QZjcuieth
/J2+PXc6J8UQDuB7L3iN6OF0IkZM5d+13RR7gA8WB8LTnVLBJjwhHV7zhaDtKEMH
Gec2qGlE9Wwho0DBnICFrwKrFdVq9Ewa2UYPC/wvEe1PlS4C4wdDaBwi2YcOUmQ7
vvY39aYJU+zay/v+9RET0GeZzqkKZLrxu2sYo7DUggsLSq5qwWBXzxWqxfBFXU6P
w/ZbmO1v7s7SJwUgpKZFg6QtkM43unuKIgf8+hwnyUDsULve+aY24F2BnCI8/9ao
rNnLInGTtOPBjAZFDOYsq3X8k9BZYF3YWj0J5cNXRY4N/XqpWiEI8N0INZ1HHF5s
5iyFajlwsPFA80mrldSzJgnOEtxhD1gZ6v2Eg10cxgr2HFCQOG7YbVhld9MxdNn3
qIJ1aGNlSFumHc3Ge4NCKijvlzuPBuOEokxK1kHktFOO86FIa3nV9u3klPsRYKoD
llxVHdiqnuZw9Xiwy94Uj375/j5fIKUKyhgRCW7tgcjuS1nn2eEIWIvp6wXGj3bP
HD8cCCHZ2MNAsolh0xpJKtuQaznasW3ep5y3qdTSmbqW0urWuFieXaqWmyPghHa7
HRBu+8KBpqo16jVNYNfvDeiwIOuWOe5g/6861CCf/SRdNUc40y8NyS/DF8pRbDlI
NOg4iWhLQxe38z11a5mTD1QYe5N3MM1KBXeqMz+KjB31zmkfWeWscYx1Ec1egVFE
O5EAPBAoOf6NG3csb10iCsAVhB94EHgBYRpTzcC3TXQgjMDcyw0X+jt9FONc2CGc
IAByQ7w9R2VU9cZzBnzRXFuApDufGrGiUHQ8XiE/yfgciCUOCSiftOD7/HZeCHGk
7XCJza4SLEFZZQkLWqRaft54hZLZ1cBTJCgqyKlzS2JBmB86N2Q25itqfxC69DZD
89I335RLGl3lr7emDPXQWo+CW76vMSl8zH/ySvt05agnRazY3JJKp5qXHyyN4IEl
mH9yRfYkXK4LjVdgP/hH23J1kOymxLbXqSgHiap10g7L1FGSi7sGuC88iqTd5ziY
T7xEKA+e1dS98sUQSemuL75YLg7BrwlPjnNQk8hLnwM+Vs9mg6BhQHlVTHyc4SSu
5SLObllBXqMPxFPgD6XfOrpboFf8fiwNGHoqukehcLfV0qnOM4+cqCeXoys6LXs/
vbwF9RZ57q7V1QrhyUeKGuoBPA2voa8w9zR0/uVgKKmf2WbZ0hNUXy1DzN5EqtRN
laLqPOSHKQ9JBuq2HWVDThNcOub2yE3BHmnGZEKIVRRvMd4C7sbI+ycnVSrHbEm4
bse+NL8zET5A6xlXz1Z0R8WsSHHjDsTUSikeTFWjEUQgnjsOt5/JquzMy6Cw8D1C
3LyyanPiUR2ED/YltNrEVys+argUm8jchASA/W5KDykEdWv3yP5SzExiw6NXo2xb
yeDR+NjHy3Yc650VfuU0z5Um5KuPNlRZNXaa87zC+ZOR2O798/7sZAlqNtVVT1kl
G6avjo4WW1ZwtL7/SX+CGFR6jvPn5TDyfEvR0EpLoORlCpEr6TpmL2gdn9qkzw+V
IF0H1SY+7tQ2pRHzzRLeEyv1teeos85oUCTtdXR1+nPXo2ZBDHrh5vzISOdTq7lQ
k1JWcMHZlq5HAZ2HI976SSh+lNEgS4v9zfnGE632zuH8C0w3COprM4zp4sb6RXMC
kmVOV7mMyHVc7Th7kqYby64wPK9aJbF3cFdeNGx9vHCBvvrMY57IAKS2W4My4Ifb
NOgsBZ8EbTSaLgCxhr5PoM52mr3L404NFi0p6Qauc9iKLFlce9PaPrsrC7hcB9/i
PC5i7R/OL8kYxzL9zgQoKEpFY81KBdAyztU4s7tRq8gVNuww6U/QvqSPNat4DqFd
OgMf0ExGpw7MFFykVTONyMb2g2zashqtsdaBP9foXNiXh2nsHHSjGDgWIuhNMKp6
wZW3qZjoW75sX5sA7G/Gbw9fgOZz44KXhCSiuDfSd//DQOYsLbHFJtRumhIe2YA/
QkZrtj98mutLdgBxzArUS3hligI+Qw39rZhDMDYHrPZkHAoxN+rgxi7eGot9R3IQ
fRIAnQEUVXgjZCPlAJnKq2XZhpe1MM8Qe7Yzf+xNrUz2kiVe+ilx/HgKrsF+9KDi
TbxdvKeudwTuZKmG/vdWgYQhG2QtHkpYqKtTu0XIwAJ/ErReQUqI8DtIwO7v2FsQ
cQwbPqbD9LuI8auSUNcB4HOlbFE6xAAKRdHJmrOAmtbltxSb+5U8+U63Jj+UG/6t
lMt3lPuygPvCZU54iJWVDf3CGUQHFVuw8mph49H117Eq4wa4+NuIg2EopFqZQqaw
oXuhflcziyJ7P+GACcoocUAc+YdsdfALLl5zVa66LC3ICOD5Cy8jTFdv0sqrMgZd
zGgxov6imdsAjIjmF/S7VgzzcXZICCDNlg2+1OaWba7cVZnNwx+Re1luaMKV5ARF
AqJkG9SAHBEkEefpEz+VCGNE4HeVy0Eg1gZ5AE+uAeX5AW9usuVtIihAv++aZx98
tydGdxS1LK13E9P2JuQcyrOY0tyRBxZSYt/qO4VVDTbGsenkQqgRE5A+ghstHdZC
BWWVlMhIRFARwzE+FU8Yo0y39VhSCAhIliyR9DGnMbiA3PLhffTCeGi8H8ALhiBF
qKjoTdZfKzv2DN9LHbmHLJmkDmOZ0IxnoZa961ZcuLUUwlsjYFi7cf+hhlWOZweH
wgDZs00la3WIGUOHAdd42YBFBBT0uJ6Jnz+40oP/7IqQzsedFjy2X47Yj6qlCybw
iciBD6UOgu2u06f+MOOZ6nx6JRAISdKQTB9YBREWyjCwCwJMO5Kz+BFBYKHjf1kL
e9CaBtJGKwbjRPE0nfH4R3p6p+yNgEL0sC9HS4K9x6sd75eIhFOiEvcXcqp5HW7t
vzXywVK7l9lAA8rqM5GX6ETVJ9zvdm2eE1PoVeLaj6SGogu3UGm7lhrn2+iCHnDG
Pdgm7PqsW/niKnia4mQTGErTBsXT83Yb5YLi+kBfX0NX7F/mO0cW1z5HYg84pAIo
9lUeB/zpxxfP8FwoRV8zcZ3qAn1qtH1mVTRHccxOoW1a1lp3Vqzs6tY1CpzQMWeO
odDSAWg/7+Y7G36S5XHGwnK0Z/rhrrwGJt7zWk6D2/6jWyIp7j6feSo73PJuUms0
clr5qrQU0vsPXCQAxFLczPLwm8UujFE4ANwve0yJOKgA19zoMX3QbpNasNg1ee7H
YK65MH1QTiPY6CTL6U0cjsLv96tpCuloO4K7Tn7r5mTiRvcZQMW+2tL9O2XwLiTS
EOXLljRsnTI9ewABmtKHkk1gvG9gB8QMu36kW//aZqc0NUvqZTEx8qKC39mp1hkM
dhtzCN9nOZPOErDQ1eVXw5deN2cEIHmv/k/usKecDN1hvODKZpRvgR/9Y6ONa5i4
/8dHfRcdY3zDjv0qssGRhEftTIIrVJltWBH782noe5nDDK9cbWyzlgEheRh4Wzsn
gsuCj18CqWfv5IgcKObuFwYXA8NghNYb3BUqn5G2QzyafOwDtaUdnct+CoO+pSwK
RmUN+knihSKJe/gf0IoUam73gPCX5AjcITLnBsKR/8VVU5tAAyC/QmuqisdIbxCA
d1SOY/jiBzFzbWpN7SITsKLmVarfC5LM91NTbAViscUmJz0hotR+pA4deaUIhhvO
YoqxlxagH3YDFIqIJENtvBW3PH1NW44h72Z2oEvHG8NzofMvEOqwfj2ygjhlxs92
5R/cYnZGeQk8ogppiThAkRL5OrljuOEYhsmohoMeHAFL8DYTFt+2TKe1H0Jkd0S6
ijF5FFqUBgkZgcODZUkABaNqBLj+PZrzV/dGpJIirYrf247gbMKsC6IaAfbe5ow9
UwklawGAY6eVRRydtt+JS2BxlTYD6ARwKZTCniK71TTuwjP4wGzZcj/eoa+rZux5
bR5BBjP2AjguEsc39RYbCVQ4wMPbQa+v08MYj3DCR8W0HDUZsga0S0aetbuE7Z4n
6YIUD3NmFhiKsURRR3VHAQWFyP4gybhvIYVU+RDc3o8k5k1V2Ir9MeunuCNnPciW
b780yxxy36rdhE+JyQITtudPCT/0PV3PvBVoAVnM5BPUlrgkTKmx+uXEQI7lBKRI
zReL7wubpRuGV5RPydjysWfuChhUr5V97lT7HKDlY7jj/3ul8G48omf6LY1jl6D6
YfMmgKu0wTIsWCamgz+gmYptLQY+akQb3zXzycUp3ifXs4YTrSzwIo6Ef5vFYcCA
7faLCr3rFALCWfCHC5iM6LT93hDIHOTeG59jB48bVmdAX399RR1b9fTfmdOwzHPc
NgWOSxzC+fqmu+mC3v2v0aTounP/NB0L2VOEZF8MjUAfOk3wIZ7SSB9S+YWsZf+8
y9Catlfn3b0TiCrgGngrhMcN8MRMomtvdgYSFtvpACJPuG3pK3yVY6P/t2/JyAF6
oyKCA1rzy36vL7oXbd7wOuF2jktfNSB/CPsQQBL769HMgerDBPl3RLlj/pYKGsFB
FHgM06u+bkQcX3LoWY+wG5QtYcMb9IFMIUunmd7dNVEjDIiH+J97IfSi+PuqQCg9
ADnZfiDzwZvAMq58puUfEIh+OGm7re2n8k2FDn7WR3kDC9rdPuu5CUyd23N2RyQH
UkJ/QVhsoa8AuyMo+coZBpmwPFlwcgLaw+n+r7mdzVkHbn3EmQT6VVkcfrDSEtWc
icwbAmoM1jx3fpS0pVqJbuiG5a1RUcjWLRow9LhYm4SQYyKB6mXXEO3RDSkmhPsn
coD9mBk0FlJQGOTFR+CVHXp0EOQQtCRpUKy6h3YLHO4GIAtIcer//6Ikr7+cNbJR
EfOjD0LvHQAqxkp7tDOAiTfAE8QYwaZ6Y39ASiNGvZfDP2LE2y5Gbq8fyNRbnbtn
uX0QbVNMlpkoC3UpuvpuqBAKwYWk+KUQA8RWROYQIJ5481xkaFv3G6qAp9paMEaJ
Mt/UI9zvmpyVJgG9/PB1geomvNHqYeHitXS1iS0tDa2z8jTJWGFT9rem6uzHR4uf
30u09AsFHS9nYy4Rc8e3qAQ8mtm0mZePXTc5nG4tW4cyhpqnwveg+FUiXQm+7Yyj
CVY7+XwVTCmu8FvOP/KP39uGyN98iMv+cdC04UhqKUZgYnq+oLXhn2+SXEXTnyIB
vnlNEeX1UQQOF1qMX6JpdYnPU/4kpI5T/lum1vps8Ifvr9XzTJjty1p0GGCifhMo
uqSd1FSO8pqf/Rv5TupjSUXxzS6gZm6eWEo/QoZFjHPerF96G+LStls1vHq2wCqL
Xj6YsWhu6XFH4iGidP2gZ8ybTFP+aj3gkS3KT21q7ef2/hVOMhvU5lJIQQ+GqXrk
KZE3q4vqQzT4M1no76wnQajqQvjk1H2HsCyUnNkDTTLBz/N3/LFytGjtrvZzuSMD
P/z+bT4hBQMA9WWegm9RLFsE5fhTLv25XaRri19niKZIJBVF3CzPxiZ0BQi1tzNS
tw61WtBnyiJtkwJkcagc79fsR7aVFJYULEyL9Klw6tfTq1tke6kjC6ZnKb0eumcl
SsKdUwND3JeVojJ52sI722EO8OKdEjQVyRzBIRhe+gCFkA3WDDwybhpjrDHyRXCI
B6UdgpnaPMwIIz5M9ilVfU2TmXIpiTIXEe25+XhIzV4Q+MyRPddH2wiTAzivToSn
CGhbILhnNQZY0CIMv3wQQCnZ8IDJxX09xdbKYsAByhNyqtC9todKNlvBaY7CELRu
qDS724mTZDmXAEDi2Rafc4uJV/ENEbShIpyL2gilLl9ftB9aAPTZbqGu/jwxALCf
SDljRgDzbUuZct3WrNrNNk9N8yJ1FvbRVYGM8CJNPAtJGX6dKcDuFSUwxOEsFW/K
tcL58i6fEw4MTBsDRxmmnVqpokPbaiYpYo+jgkXAbkStmH2KFCZO4jqTsPKHnkQE
Fb4hROCWoUDFPOA/HEGwYkoRJ3XeOhD/CDluZ+zPEBx6j2u5BiQwA+iSpOFLGbgV
orufcuNru9hJNAi3ktlhIQJrYwGNfo60J7RewR16sLRZPMq3+QHuJQQl+RF/MNTf
6qAub/kAsYei80O6A6mqqIf3AYyJxNu+bamsVw9yRH9or5F/52rPW0rL+zJALL/g
ewaOFT6ZI/aUo4OGklac77AgPLZc3QBCDwqEcZblgsULc8UrXuy5pZ4M2d3c1z4O
ePRQuuLG/FxkaUpoq7Hz3rPEj7hw8PUzpR9m0RVMcsRXtYLK7vJa0MiLp3qSuoqt
9vC/Wb4AUdpTTXS8ATwvsN6RkI4BbyLuD+HwszBPXVsFZ4d42pMq1TVSZvwxb+Si
jrYrwQKvnSzaecuQxaMvHBEOaOGYtphnCnFLh5GEe8pLGeiZ/6xfrLlS2i1yGejj
lNVHKveHi2mKwUepCMEc3X9CZ5XtfiX2BWqmDzPII6sQuS0SsY8I5tdYakkH2Gjs
IDW5zH3PMwv1MqF/FZF8AQM41DWRrCY1+y2qeU5qrdmKsC5maYJvCwnjz3GYM3LM
DLCMK9ONhTK9QgNN7fPuoD2Q9v1o3o6P7f7pKpuKuM7FVagBeHhoJGrWlAn3VJT/
yC5Y89ZOp6QrtcbMO2+GjaCcgjgfkywqP1/N2rxpJt/8KfJ+TWNOkmSevx7rvQXF
/DZK+G7l/7LMDXQCkc8b7SDTuruPmGSVh09FhvuSYhahBCyDIAUclH5PM8MB0e8I
hvQakW5Pip/HFyaMDprG4czDPB4+kSoqy+Pna/8xETuNJhoCgwohXyXiE4AsqQfV
Ya6SoxY6bfvyavX/7YPoplK9BdfiYyw7kDg6M8E1IG8qMw9tnCz5SyDuRH439E2S
ikzjxRWTAlxo9ODhyVs0R/YuhNE8/Qsi+V349pdiqv1y8tF2Ay0zevj3Wp1FAffk
asZwg//26kbWWUjXVkIWUczip5KZRH/ENAwX2vYFm6ZU3hYy5hxf7R277XrOIVZV
hSgaaaRXXC72GxkRuQeR6b9ZqpMnPfVHVRpshvhprvd+Y12c02GMpTkpD/Sntvfk
bBWSTaoprGPP1pDvdAZHAkTt6vwpAG/QWsdgoYn+QuyrAHSbk+ITr7cOAr17uwLR
Vfwqg1uqueAlK/TN3a/ExDjjSbm3gdXofd3WRMjWCbXuZvH9An4PKPpYyT17dH5Y
OpZ6hfFZxbFMO/JlL16djcgoSHp1E41os4mCK01mVEU2fv8xK8CakpcvmqzOSx2h
v5h8LskpHisKm+jhBJvEYbPDbL+lvCeF4qZ0xeSA7827KIMoxhFBfgdSq5jfzH3o
IXlJpkmS0KU9iaMt63LoTJ1NMnuzv7jZ/tE8gNfENNjLzUCTaIPM+GMduYFQYBy6
Tom+K9PSg7Ih4fkMkx5FGv52GCszLqkBAUUSv68Z1u5V5BAZsFpB2gemiTb/ZGb/
8tlpPNKpFbglbTw5mv1B/OjInxqok50fISFWbZDlWTgCwbxf1yp5BQc1BQ5usB6l
6dj3RpOEVFtVCBbxJRxus/84jayRx3k9WxUTukco/UM0/is0stKIWqJ42lKFFT5v
IAdoz8t5R7t2p8wFTwja2fP4RsMNC0F+Yq5bmNUBF/ZTYlhis62c/TiSMs2K6Xlm
y2+6qaHce6lONW2+RB+JdmPbJfHJxNf8mICNVlhi91uJiLT7MAGa63OiWletgOqd
RC/FzUxcuz/U/c9AbT3OvJFqgjYGTdRBvtWy4A8f0O6RQd8YaP12xERybIEEiFqS
Dfhr55hQ5qugBugEhw75kGLR6XLqU6xDqs77TN8OC1QlZyWvCbM9QfKNH5E+a8sB
d5sJi1KqfFdZ8y/vdAsjOSuNlKfKLeVXXT0Lju8279vzARwGwFNxsIcLDo9vq5Pf
+rm/yomAWTPU9hJ85bsXONwK61DWuW1UZkFYowsAnyeUnudTBIws8HfgDT7UfQWg
UPjQYIi+YhpPvuzRZh9RAuL3dhNyp+FNZJPz++a9m+rvSrDDM0x0YrGt95e8B9wI
Ow+MgIsgMaP5rz8qYIDboN5ECTi4J/0JNhswlMhT3yQQy7KCyVyw2Ik7YeaXjxx9
16yCj8KW3HwXYZ1tAcCj8Z2YFxtxJceUyDHUaUF5i1yKOxCgxEJVjiyqQM8vugZj
uF/JTwC9Lp//7qj0/RcGM38MVaCHKe6g/U0WZucp4+zIakTsmlWpeDHrRlOojIto
dB40M8XKW2b6MpjV97g05bfMeWprE8NZL612UqJ2B5Aply7kdEAICv/g2aNFO5uv
DLQtu4sPYub3XJS0zPWakySRzlGeBIpuvIic5MvZGcSndlq8B+snxCeQJcrSquCd
YotRONe+M0nZ0SF3HP7bZkuTND04m0R96iUdIYGANUer3WDcrHcbqJ3QwzpXy5ZL
F0Dt/o0retqpH1xZtMESrVKTgiFxnFZKfJWRoJPPF8p2ouauAWZX7FOVZthDCSL+
tvYv+gEREaRBuK+5vnKctS20NV7pq9jaQmx0xFDvSLVt6LgbPYP8YEjwWG0g0g7m
dGPzNhip5BG7sBK6phHq3WBgLfn8ehCudOiqE9vs2+c7WGyMHjWHATpFF8eM8rtc
b79RbbPQ7r5ZV+AXRAC36HLWO9td1UkJXjm+Gykg+9iWj5fksB2v+5+T1qDgKcFG
3btQq+f5GDcaJCnvwhbJ7dd0NGX8OYtLD4E31V4+Wy5ZMxjjBMJgG5JX+vL6usaM
AhlQAo6m+qVoc8TouMr6pTci7yl7QhmiPCnUIbap/vpBnBYqYjaBdVGRygXTbWdN
ZV8bTl2VjGaVzH+EInrxQqyNUMm6zdrR4ovqEEsZsmP4LnYEdvoMbk8pT4JS4zq5
iFKvRePFBp3pjpFG3cLPXpiawCd/kvMIfAWR3cG3YEF9DEqDH3T6ZwkKOmMzEeDy
LJkWHdvcUPHRvEs08LwhIy3wAKStJbLpmqJhqafMgJVEpZkZ6LQi8PTzu1QukDmX
HdgLv5w8QBwQsta21v4zoPIhpmKSJEuSGCA0b6aT1c6scZiEIF3BcZ0CeU3F6erD
wqprgmyALB7Pe13hQxOWguGig+Z4LO0DYZRCufQn+cn/HVjSuEx6lEeL/Hoqal2w
ZJvu6cii4OOl8vjRlyNvCogtbRU51cA83qBijRvGW45kkW3A3Tc9L6TUIuQDVoAe
aiKgHLJeqm0Ag3nH15NGtgRk4NM7Sn5Tx2VWYy/B//fkhQYr2VNz5aILn24YQBjK
3z0/x+SzBOphrHKWDj536WwTAa9oMMeSoNv9YGdcUfc3Mki1bkN74cI8uIkjcBKc
vvtCbWWamzzIHt5pHK3cIHu/CaJmb9Dm9bIm5i2N82vA6BgKCdCq8EjtY+NbE+D5
II5FkU+z7LG1YhOlPY9rnNOetnm5a11VQF2oxwT/hBUimYmSqfXFM1Oce+B4Pytl
NROO0p7Ds5aooc+SGExGelmMJsHjLtnL5OjkJFcYE06QqdcQ7lrU0iOghnXQH9Uz
dsHFcHiusKOgpARp+aGSIGy2gzTKodBwf9VczyQknnmU3NlQhhbaSc10Dzv7gaPF
xybYKhDexxdOR0M2uyNIP0iKOETnD+vPwDL6mgxN6iLCyvflYqegMzu72U9kC3ec
GW8+sRRZCyhVIp0fCXrVXFf8qdjgP/skVYtO+IIhwdHdqGK79MTkB4zUT4YEEwwv
ZIN/C+YF3BSxztt3wslNYL2PHkNfCi9eoQxrUC8iy8KtOJAHcIzcAepn+o9DHwp3
T7FEELA3r0tDl7qXyJIIgX/plcn0pN/o7BQkKNThTt4Jo8JGfoSoLI3D6kLLONB5
FmC9srdRUb/+hYFAWTbXFOCCcu1X/sEMPo2C5L90YITY+A9jl4TQyVndhAnMFyBA
Gr6kM4GtaGkbpzp5f4d7qYpI+GyNOAmCaXYtfPSuNEn2iJO8EbRmzLwCC5LfztLZ
WbHCCLgUmMdtwFfZyJk6hhfsSB4k5XfZXWBo4fdWhQh/UgBqqzkoAddhAnUyivHD
cEs2qfyyIXv6SSyVw5IShl5ldYUE/9kVi25y2uVqXgDnMJkeJOQXefHQ30uKE/8I
JjBzO8NnSDzO/0EEHg51SEBYrjRlK7+hgCX0vokMnOofAvHWaWk/Qq78p60rChES
C7qj/6ehnqYSPVfQregeXgOS3ZmQIqf25XqdPxTZ2QZSxAEPm1ka79G9gJj5Ymjt
CNq79J2qTiSHcURsAqOeClGBNwBy0s1An1ZJnhXvjrdMy0SjbqWlO9x/L6BoJd6l
TBNzZ2B0NMkcwIOfIeKcxMbBR/U0OhIKuO+2J7qN9mFT3r9pRxsoL/CH1UrzVV++
40x1wG41ADJz7FEwWrjy+mnl3VB4BB+WrJ4a7YpwL5Uk5Gm6s29iZHKDnRajrTGt
SpDEaOcwhuQGIuKYaHn/FulC3EYDsK2uS6Q6ACBhwUbFfOhb4E2WHop8KTfqGMcK
acEUP89wMu/SYy49GEPa0RAE/dE9iLjKgUanrEZ2GkNMmCJdC0NAAOi/t3/JdVES
eMw4Is8r3e1b3irxMFAxsdWjTgey6zuqtaYFnuq+M7JYb0coXKehMECRtvSKda44
jLn2wbRCRhzPyAzPNvIiCMmcQhDacw2JwhUY3eM4/VgOvyBm/z74Bhi8bZJpky4C
tBa74DgmAUG+VsvJElC4CaHPDm0F7K70hurFG2sa/VWr2kgJIboMW+ZwbYv3h9Dx
QRvZ3iF6XYVCk5AL/7Ku7VBL2KM0IOkYi4hC+rH3nmC18sJyfwaA3WYov7rc+0Hv
hOJBAo2R1AH1Z3nAa1NJC0N8YFeHfeC4MLuXJBXfeGrE4sqro4MTrvWkhNF7CQPc
laJxpJhkId4cBY5xxO2H6XJWD5CLWAVbDKZ3dq7uAdPgFdBZjNx2HDrVSF5Rze5U
4CtvjbxD2ZGAeFswDunJ281VUFP8YIaR+EbTpEECgoz6DQKcsVO9/wFBmBU73A87
V2WwhOQsmcVRpUSJyC5+d1NqxGpT2gaNHhfFRvjj7sPqCWHClXwVtmxx+2LPLMZx
cZLt+8vAxqU/FBYmuus36wYlFUjbi7j338yBbOOLRQo6VZ9ctrASP2yZ7TYscCzv
N0QHPZgSHaqh6aDmK1719cXjzuo+wvs1lOj7p5614tjR0G6KI5tLCJyC/ERP66DJ
S8N4S36CyLMJzSMECWTMIZIfjSe4IuiEBIOxHDqEENI0qfOY8uo5gRHYf2VI4XF9
gAliJ2mlHDAifevxSUXjjhp4AExH9ATugJh7G0aGP4QkWwPbIm9U78BqVytWO2ni
8rEVhU8mGy6zJ/FY3xqyLTNNMiovjnAxZS0aiW2D759YJPxCrkrzd8MLe+CkUivo
F14zDe9DWpXjRD6u6wNaX9RrRNKF1/6ceQkkYonFDpDQvp3S+46jp/G+ysYJUBh6
NggXT60SHBAgAVwIqu+xVcxZlcRhPK9oOXlzbcKQkSSj7w0xc8RCFpvGxHZJDros
08rMzSwUxpvhU8IF/X3aDgYCdLj8ueyWM82nvKR8qt2W4owI/j9Q4d2a0EoUcalb
IHQljEQT/1E1S8lT+S2fd/9E7FslWCqp5LUPIO1rtcNVvEbPewCuxYCL9D/ZdWGO
YxQWOtJel2Hn13trGxdQ8eirpe0w6+zFM7GGT9iJxdqPFi+NnTnRQxKUbhgX2dJD
Ws4peZYYoY5+1x12RIUAhGmIBwAzkdUEaH6/wiy9hHIpuS9++oZPQHUGLHixZHfv
jNKkSYSn5Dt8d+mPUf/VKuqJw93hKZUU1IlUW3wTzqGiCGwiBwKk1h2Bue+a1BC/
VJNy19TRrAx2YWUZAxWd2Q7gSMcoVRkv01lYQMcNyp14oS7NoPqRbcmvnRM52RYK
V6ttBZMPRExXKFBElhcOyRIc8eyzccYuNQ4LcXTI6v990ez82yG2S7WDQobjDiFk
muK1ZOljYFwtzemDWdNr1O0xq5poql0IRefv+RVeJYz4uG8jrwyFfGfg/ZGOxW6L
kPckX12tinZASGq9PFh1ZmDdg4usfdaAJIGLwf4/JQZvmz+rR9g+BZQaQSDeI5kH
cqHP1KNlCbMix/kKceT28vM19/j0g8XaUUhIjZTfUlQpfafMYnf28MRFoAwOpbSW
b5HNZgNuJYsiKBOLDl2/RdgCMuE7JJ7ODHufj/hWJcwdfnfA/6yQlVJyWTWVVmQM
WeAb8tyG6KSMnZHThzDMisnIm4gC24gygbDsMhBt+XLEFBt+eOgcKaSFp5hCq7hJ
TrTs+aq68GojhuYiYp8krQPABbweWrRbXqTVujGizZntJ+1HuFNQbpimPsFikEYH
Z3Vi1LZToTXgqxP42OdXqLqSzY5h/BCGaEPPtWeNEe/S9g/AybxPUXtOgxDwT4bx
CHvZfw43MkuKquMeWdOdUFewLXvb+DFgyKV0rJ9lZZ+BY1NGUlM2Dt3v4d4yRaqo
ulmytIJOfeA30NTma6JzXCVmlLzfZeA9muXN01H7YwMNao0wyKpr+LDa/7K/zMx0
pU29sjqk12btBGdmAcZJG87kTawzR4IE7rwChE3lhwnGuGqrL3z0/NQDEeuHxruU
VqcSLXqa8PL3kUcqM+1iNbLoyg7u6TyvzxFtQHn39nH7DP2AOWKeLtt6yfEVwzjd
zvAdkRGp9kzwde2D9BansZfmJSKmkZ7jDWBrgBw5SZEXp788LJpg2Y36YlhEWrz3
2hCGgpRV1eLoi7J9oW6cYCO8hpFb3cuVp6f0N3kM4GS3jT9Bf7PLMhJGfbtiqLLN
wWN9sIpxuPQwR/qnddLdBjoOnE9gKTlNDj3BbfL2khQd1KQCzm56cYNms3GSdpFr
a3gfW7cePwZNQrenO7mruR2bQktDZ+GJJoBswrSXKNGXBlMVhUEu6mfQ6NY4YfSC
wrY71h53sReELHcprkV47w9EiIw2l6Pg0YKjcx0Bm7smFZ1alvQTEFP8CQMcwnMI
vz/095yv8nslmkUpyCmQQNdJkgqsI0lBS1iJ9yGv010LtZzeWhJDsIr56fQiGKSv
mc/lgrycbbw35W50NzMg7yPJybKiLs4VwDJhELqvftuinV2YJ0Re0DaVQzrEzOiH
1e3gk3w6MHND4fP9N5m/wzNGKVI64x/i7qfh/A3ra50m7FcwkeKzFpPDEB/PzvrW
m8VSSbLQ2DSet8PT2+pCD4nQidPdq12r99MLgH9hfMu4gnWx4d+HkSSM49YTQECF
Effx215zQr46VDErxHesjDFkYVWFKl+ibzYvMswwoERTOSG5USAFDAWZi9HUJB6G
GvdXYiE2y2U3rJjA7vqWLG2/lNKC6kYqWXz2I7XZl9out1lezmqQnesFqYxP7dcn
bB8VQDJXyBsQ4XXqevNKs+OMkx32aoWEW8A6FiZfT+/ETItPm1M+CNWU9vI1W23D
TN/qLpl1vZTySrRGuivORZaeEuDnMG7ls42CPtmAjrNRNTvS5Q+faY62KN5sjM4B
kPnWwn20XIWyN4hZQO+WchUTpgu+AdX8hoK1wQSdTbUjwHnTBG06CGlAtz0cQXHX
M25aNnEYpc7c2fDbi9fb5IlFToH0vinSiDQQREOK+0W18s7YS7YD0vyaG2JmCL2M
HTMa/GDghofm18A1xAAP1xmmTn/+8o/dDbbQxRGCNTwdHsAb7DNotR+m++R8NWg9
WdvF9e3qxIjwFaUX3uj9ta/6KqUUfy02Wq5mbZrrPVWM4Y49pFXWiwUku1Qqvhft
yY/K62RqcIc7jIX9+UC2xx/vLttgue8EGgqeA6mbA12LORG8xwmWVentFNL9MmVk
7BoT7N21srVWo6rkKUrM6Jt5yqV1N3LUQLCUo7VxDrCHLhCxVDijgO0X7jI/tWSJ
I0+S5nhBnHUDI39Gj8yhV3KWCX0AszuC+ODb5iSCOc5XJ0ToB6szxe1XUPSzKlzd
fKfnF9R8KttLcA2mvo74Zwqi+YxywY7BUB2r+VZMaH8lQ9TSob0oyE7jsYq1xJm6
SbLzw0t+pxf+uKx37rynk2dGmqkutX901Df1hzfuOHGQFk6QNVe26vkXc1bwpBig
HIO9LGLy3iTWq6JQVsTdQtgW4gex8bC6Kbu4YwSxw6PpSyTwV4vTStM/bXbP09OW
g2/YCIeKToNbtz0+kKb3xEtg4Dkx7bvnSCqWyteIkG9w94EbbSS3xJlk9JlZhMYA
Ai2Nhw7jiSNPF8K1jGsdX9nEoEFKKYWQJaEJgzwklkIcptxWatm5t2u9YSOBj3tP
HUITfeqeE+AAH2kWjeFZnTf5g8maWhq9Y7M5f+L5rZh6GrtZiwqQhvML/yfazEmk
YdSXPGHr1xeGMFxApu6t6WkvrjghIJRV73lLxb211/TwJWkylxXW1NYXKiipuOiX
scB3JNqv4Cggk40FTm9Z+EJWSQepgaOvU/IZDqVbwELDS7lqx5E+OY9yTEqyHeJ4
6PE4dmTJ0GGt7GpHYHUNrHbFU1fQg9EiAGs+3uiFK+bJRvMwx6YXqE7wM23Bey6U
tspCo9PzgRLpRHIRLK4prqs0vl1VmiLaz92Kzp19EMDgJc1slZgKzAUfYsIX92LI
agWktCbmUvmPMV2WJ9/Xi+JrSBECeH/VBUIZ7Pr9bpAKfQJ6P1eQ5GBYUtMIp+c2
KcVaKWFB6x2Z823bkdjd3owdpuLoCRUIV8tIKIGtvQW0hLZrX9btyDvz43W8ZexB
EEH3qV0FyzAK+HJ9vOQb30mbiUNNai99e4h6+nTnj/XM1pXCArgR528pjgIx4iVf
z8fCuTMknyBCZhSk8Vh4VZJY6NBWjUXAkLqXIWQWSnPJ4Xn02tUnhFB/kp3J+8lI
T20MmwxBu1OwdSaW83wSSGHllZe8zXe6W7HVW9FqlgajE5zKSQxh0O92sZJssGkK
VE4/AMz4Y/7MPplRTTs+vgvqF7j2qTdpYQI9rpN67TEYW2tKfIEcU6GOOStItoEc
3gO4jzqYij93pgPJAi5DEzml/JAv3AJ7bxaIjNV80+OMf0QxVIHPE/zA1gzTkG3b
CvmqsbkGdm2NIUY1dOyB8n8SF0d8gSgbV2a3t1mNPNUQl9OC9HHZgemvapQeN80p
wT2ie/0Oxc74fKwfNSQDRf8kGqN1zUsdndwaqOWE6kGsf6VtLruw7lDRJZhGZD0B
t8CnG/EBqJmOEemC8k2aKFKSBd4ag/lttR+LBNHnE0SPg9Z95tFaAk69/e4xIbE7
lZcdUYsXFnM4dNtPeEyFPscDdDZKrc5uC9NwRIFauuA7bW5CdH0l2xPYm0L2LKXi
2H/BwcQ09mE8DZ4RjP9qUUCEGHCYPCh06BWtPzama9RDL1gpd20IgkIKc3nxWxAB
2hgQDZE54BEykjUPCfwwkvdlacSPOSlmsJq1pv3U8/YPxXLyVzKVcSrbyRNsgM3j
rvkTixDqsdlb6qWC8EE5d3mg3IVPqaU1vJLh9UO1dr1B5DdimhbuE+xMIdvvbHDh
U/ldvb1Blyo1nOocPY6IF+1krBNUrdRNclL7gh6XsW3IJwcmHRhnqsrUDJ5tLaGX
PSWyKWtuudhba/nAX+Ky0gFgLwVV8oDfm0TOgG612bV0h3AY3mT7bnazkUpIuIG1
iBHm2EfU81cORZoLcrdZmkFUqY4oHKlqSSqeUvffNZM0atH0qR/TysPJZsklIvKr
BZz6Xgu0a8xi+P5331BePAmZxu6dSWq78MTfYa+hhz3e6GL5CIg6OVIYdXa7AHRc
i7LR8Pv1zKwS40pMVXIT9BkJlt8tuG8LnxktG8tU15U1DTMI5QQrMqYIWlf+vLx0
0RccvbskOo9hEdW3cMKrqCJDFRrmKg/0Uh2cuOHJEK1GJ0pfyTOHElvOuWlGOyK3
F4hOzN579NCrHHG3sNcdwAwizgCG6AoWGaChwKwC1s2IzV1G2E3KSZaTKrqWEJ20
7XKXFWw5x3AiJBer0Q3KaRbRC58wjoa1Hz+wPKxrQZSPYOeTN8QoTsqZyjlvkgEl
a0em4TcaMQqpYME9doH3j3qmW5B7CkYQ0HjN1KE6xpU/iZ/oRd6Nmw09BBq28j86
FJbdMLKYqnFQFEcEtKdQYGMYDTZze4/oGXy0uGEVnYdOeNRBvRYqQOJnFjSTOl10
7ECDakh7pRVWcn1XNbPImadAIGMRVQ0schs7Roc+CZZxMcP6uBv37riLsTK+1F+F
y9VkGCkpZQsdPzY+vLQxciNxGykURX2/bbHiBCiH2zK6fOLGg6TOXLFCNF3eqFMZ
HXezseJmNY66ast1dnBn1rguOrabRWcti+q9t2PbJDkl2NVdvQxaeyLCsm0VmPmX
YBwKBiQO1m6RqCITImPjf81V37jQky8pa47r+7lF7wSvy1O+yx7t3Wshdf47m+tV
bFjbhKm+I5xWcngEz+UzG908MD1Eok7xCjhWk9/aAeSrQ6oTs14g0KW37z5due1h
7RuplrM5G72THRroLhHOHyiTpIDRNZI5hINEholtpEeX21ZqS3JYUzCZbo8ibhjK
ciqDZV+fYLGmOFt0eyxvQyHk6o64zvtLd+Rgc6FOBr18NOtB9UXm/apHNzuyYAie
ByA6HmRYe5k3TjsKFnXWrH7lcqWvdYV++9MRLafWkJ4OEW03M1xR7Cf5/3VgwCYc
554ABmfRrt65yLFn2leDkjplJcpmDB13I42Y4WalEbZDGK/5OuXNxrJ5HdGHkF9r
3LbHzRX3wlVpRSD1gtbWOp0vfi3PoYlQz4jfUF0Ht25rBI4mERd5LR37lQ7GV2Hc
tgIKNfbAvvY6to3lDpRMgfS8lEoi0NACpmMIa0bQRuCtVXjiWczkpI+kBcw8c+9y
eBFffAYF2cJofzsg+9mp2uygdwkQLwW8VLm/enAbbue5m2CRcfsG0WF/wDacOqPD
IdjsEY2fYWQOJLrqyyR456UxUo0LmXXXadpPP3wHdh+iyzOKU2oxW1WN3YzaQLJN
hlXcj7q9EbAswthuRu74IpBC9m7a4kWNqSwv+wwXIcFtb5ZRumjLy/DWv2Y097eX
WJWkl0sfrIBcyzmFrvWZCtahQVwKM35deUY76u5abS9HVwmcJDKJMELBIA5DQSQr
Fs74/Bc2OJ2Th18Y7lqD+jQ8Yg3nLWhnABHRi689JUKq64vvFI+HN/e1P++mlNYj
UVYZOX0wnV9KQB7jKeqCvhBgG5oECmy9Lms/dK7wf7hb2zwPDEJrybkCJcGLM7QB
0+Lc6p6YsQvHHRUwIfThIKlBoTSR32CO3Qh0M0wzfty281E0yoPAlY/cKyDJD0bE
vkjSUd8GenjliNISx9nWmwm3P6Pj+YUjDqrKUdwEgWqUgcdU6mIZV8GTPmX4nh8i
7MdcKT3DcODQBmMEq9zgAYEtInDtR3+xz/+FKa+dCR72PIfNHRha0rWtFrGaSi7I
An1WR04FE0Y3zpqHJfImir0RpI1JZ00QdpzhNx0QE5aiaQPE72xBmIJ9ZHMtgeOc
/UbcNwQxnudSB+cfLERsTU8oxoa+NDlHfWxlDhvMW3zpQI4s0TFLnHnhfmQLoYo0
4pJVhZxIgHbUW7u/CM5/LSJj/mQkAc5jYUfkEUjnnTRjbnFD86TkFCByK7vr4llr
4M5leZ24ymGFjOEUBYGMuuYhdyuEUzAPUVC70o0icZjYzO4SVvhOJbfzEqoXSacH
cbCRhawT/XcsTqMU3tLfyc62mbsw43UyhkUm2WXVwRL5Xg7/Ga/g0CN+is/6I6vR
9u7mrXri0PTymX/4ZgyT1NLHqJseSIBDSnKMza1F2vgrjJaQNRjP7IaXNCfCxUto
aHCGNaLITb+ccEVF/gyTR6b/JuIhSxTPZbmrt8BRdQ3YJzRvT5vn8XUbPpXnXBDM
Rn1a1YfKuzg8g1TGqHANieDhUjHEIZU/BFSedJSlUhmDR1IB+uxj2xAexciypIiI
WGZWK1UG27hBPa7FwZ5D502YZ7goqq0/Xr/Dl6QsBjK1aImqjSEFsER2NKagZ2zT
7fpgPQQ1xgM7B4oiOGtQ2aLlqUbhA3qUQjOEyD3kiOPCrdbp19sGjXzEDLohlAIM
byBNqnXY+RgJUMpSRxPlJUfyQnSJycycaytr44zKLW0HPUrStECAwAqcAdj7v5Mh
snBmPsVbOUzHpL4KUIxeuq3S37/Mj1CapLXpbxabK76myVoWrH6u6iC98dATRITk
XVaiI23aBNK/USydtiWmP65MsrL0sNnk9RvPSdWBhLgEh1azBH9q6XS5ZnB7fgnl
NnV2HxyKTKnGT6AGyiLsethi8s0mwEVOEja6DWVR3yQYT09rZqpCg4qzqhlFwU6I
aKHi2wU3YHdhBGmA7FNIuz47pa7RMcR1KjHgWUcdOZ8QBaDdcehDhOTzfIinf31A
d7MfuAyMu6EetE7KHQcrUkt5sPYjGOIdJkrSAHIqq5wZub1Sfq4cUZ/HSipDof+l
mCEgY9lvlYrPlBoTLg/Q5LDS8tyrEmnJTGRDLnodEM8CiWnKaRZIhCd4K+Y3B4bg
y83TQzIZH4D1GBVIQ0EGjCbX0O41ujJVJYfuCoenK5NF+qcx2t6RO/Mo2ofccQfk
Rh4G10AJ+W1aWgs3E6qiwcOnq77i4L+YW6j7OPkVoGmsh8xzKAS8vvQg2i8V3ZqS
270B0WpThnn4eNug6TU19g7/hY0vZ6Qhtv1UMpVwDCvA6igBvkCsuVFTMpK3eNSD
lg3ndCKwCiZIah/AB1dU6wLW4jg7ZKRq5g/ByBeMQ1PPF62UM4EEwkv+kMTkYjaJ
asJRRB4Tu1oh4TodUnPuYjfftQtsmp2YDEJkRWi9UFK5IiAC+1I88114rPgZhzNc
9qG9IHtL+7SDX/HBmAGy7j6m8Hu+D/VGDcGw+0h6r+g1YoRRv/gCi37MBTsqYzYV
P+y6aNjjSeqmg2+WzrwqKC2tW/2EI3xh/9t78XnLJKh9Uyah+iS78vCnb/4nO87e
lz+GaZFrWJu2GdkZTlcAfPbzdf/5TXOJ0nQVgXnlzQ5qyjcNyAZ2cdRkt34zXxrU
hqynsjeG7SaXMpVe7ueKdfTV7oBVt67lt8YOpgYQZv+0qWRTvIy2GdsTvAgxXtQG
lH9/f3eHvxw9cU9znnCxYqN4F0MxlbbieGZKER6P+lFuvH8hPf7ohpy5ax/iJbgh
eFkn8ssYOZsAGGz94TyTs5Htnj0cttE1eDahtlsD3fsu+SbRnEy3r7VrXxb0ZtRM
UYiD7ExVc8KxsLRvKKHG1v4thVwMFu7MQp5kNwxEL6ZxYIXxpP6XswOrmlDXAcwL
jos+/ytmdQSgIlwSE1dLD6HBH9LKET9yN/EZvyh1lWPSTObOZCP9FBYTTeuegTa7
GbwrVjRg9x1frxlPIhsxXjbZTe/Py2UO80HhN6pM44eCPCkOUkvTNCb3sSRRwB4R
8c6XiAD/Yj4PJuG859kADlN2KYJWYZNIv08RyzuDcoFrxElcanx0Wi9KKOjhSeA+
0a0zlOvArWznFvCLrd7vJdkuSLa/DcdodD27AZUBOWWZtHy7Gq3wC8d1DW3mlHmh
dcLWT6int+i+CJqmxYAqDZDd93Mwqy5SZ9UFmQ42NXzU9877KRxQW6z+uGLEbztR
934lSOqORn2ocILLyToGA0IBoBwhEylWS9JX8XmEHrHZ+3k+D+2hpOAypLolla4u
+Y4TVOvVUG64fZm2dJTw1/6VZ+Q1siLdGzkFzAsEdlaRJHhyd9hMfykxpgR4qJwU
noVQ4Elbn2ch4C5JXwu9GesyiZhMUWBvgV1m8VpGAhIqGyGIGj2OghiCWTLoBuyJ
G8IPWlmjef3zUeo0/tOXvluKvUQ0XiXtFC4043xBjRkIh+KPeb4zkFEA93si3FSj
/jnbOv+dyJRoNs1lSIdJBRIn0zj+yvd0KSwMVUNLK41LRzMs5Uux47bA/kEs30Fk
r7wS4WR5HRMzW+yty+U1TabYVSCLtRzeqUIw9zqXjP7hSptlDNKRee9BAibMFg7X
WXgtWMqfM8gdxWaeU1rvc215umGDmOfRyFobeUnYjehFvmJwGsBmAD/djyk3u9kn
IUB8okpiUXMdFs4CUw42U+ljZ3sxkmjFwUShmZg/GUbSSQXaB3PAX+ut/TEX6P49
Fgyq+FpwLcHS5eRYynfigpKaJxFbBHIOJcf0ZTYIC05vpeizzg/KeBMx2Z6/rteU
1vLr//tt1kGn+67uWBHcoe5Cew9GH8zOculmZTZNofqTwp5frAn6LvB+nOdH/an8
4doq3512Rgmdnjy/vXsjlS10Rkc7CtipFhCtEk27yEfaVZn0Bin5WXJ+w9swX02X
sSR69BkImqtA/14X1Xd6oX8bsc5t4U3YuLtKJvb/wT+XMSz76r+wG1BIsJG8A6f5
HQhHqdbtLupvwBITgHDZ6iui82ofSjcKGKV7J7BKd5JEckeiJYD9uW7rdPQR7XVz
rY88GycDGnC8i8u02h8NRpER1hkWdQ6yRqp/K06MO0YRH0GGE1lNE+bgVz4CNPOi
ZicOisRgc99dDYg5xKPFYmlGVtWd+7CAFUNsV0AW8ws9mVbahddhdj7wpnoRHuFt
ZLPS2d5bcrRB3spy17aAiYfIjqjwWhILKRu6zknUO07oJZ84jdV1Ln+yJfMKhOzf
UBXLwlKz/kqdMKBouqgItaRnouXm5lgSqts7veLzuFtUvvmpm560QIaifp8UKEPZ
B5lsbYdwXhg/DWkpBZmIzZCNIAxpicJ7S7kUyZDJfnZiZTMzrjUFlwWKn7wHLC9Q
ELbHEoglbCc382imEGp1hpKLGK+F1NKgVqjbR6Eh+hczobJDqFH/Pa/HZK1haCQL
KsAe/h8eEZvO63eRv1UE0GxDpZ3IZMbE4NEtmaqK7MEfHnB5VHihb/dfcS00DoOf
GIicl2Mv2H61hjf+oA4PSdj9bDB96AEKs03zJig5ZZ9zKcb9FnY4YROumUeGUmSy
fe12C6XIEYgPrMu7LkXSP49S7MFpla14x79nKrXSj6viSWj3jF206pgmedMN+6Xr
Wjt+pMGC5SEmaW/LbhJzs5Y7icYtKyXfGqsuuiw22mmBJcMwX5GXTejkspYtrVwZ
piSbDLY2Clty4FL1G+utKFESNEuNTu7hTjHHYY97GGXqiegNP8lsKw29/KRZO8Jz
/rGRMRvMmYo1H/lJaEesKK/mLOD1H/XDVl+BX34/rZssOzsYWqCwdWx2fvKzZKGw
4bI1nCEMecn2iE7pSVwH1VY2FkMPkG/da1cvklQcNrxQfbglyN72pCRavl0t3I29
VbzBFoj9x6nfKlFIYw3DaAwZ1HBUpVmyfoln1DqkFogTjdG23Xoz+g9mgCSUGwfy
mJepScBixfS7g1dlogsvjRfcJ/zxINlyvVdOI3Fv0iP3FrpjhuwQ6PtJ96XpPwbT
MDBadf1oxwzuQMMFa3ivxqlhvrdNj9LvGyb8lEHeU6CcDgG4ZTld+QVhAz+NHGGv
d6UaJRPFotUzoN1tbwB5wVKZwn5ZjjpevyNW4ZjCO7jftCSE+pHnsedmIX2vECCL
LqFvzVKY/tv3jh2Gyf3lRxXDYQWJIkysBOry8Z6KKgaTHf+UVjos2cw5IqzkhjeK
R/EtSL1YuWw0WDgXsNkpa+o2SxeL56P9KCCjeRqig+LMBekJn/iMVTmvRd6bwwn5
Egw0mt/YElycCFKCErur94ubjjqWmOfqsgCS22fZhhqtW0ZnNBrhY/3sYLpCns9O
xVKL6PFs66o1xENCjoV+e9sZx3Q1g5omN/Suc9cjqmlG9aKfKH0oGQz4jenN2XFv
p4D05G0bI3B87XQRkvVSnEywXNHIQa9X7rWBHau4JmcmALfMEJRcokhLYHRN9E0z
k1bXsZYcPLjMtshYb1vcywH8e+bKeRgNalkP5t1dnakfPnBOzfO8PnU39YkTKJw/
QVrHy9/KcAIEJmEHjC9HC+SEWVt6ZHyny/kHJvZ9xsNF0AQlangVsVbIwyZno1IE
4Bjj7/2EcmUwAbhj0fou5iOjQ6SMtZO3e3nzsRJBusRvjS2C18Ogm9yDbuMqlFKZ
+sSOekdfiYj7ZZB2JApzria+k3lKrgPB6OH1ORzhpvoPd2p0cc8DsGu9yFtldQvf
ZvX4ALswerjDGVXbkRQUndvnZI9wVZPqQfQZN402/J3X85SJUajN5DuxnDgD9hre
CG4uHWvYIMipShTZyG+lDDYj/lijMvYTopVvRRcaej3n6CDSX2jEwv6RPD98Cjki
gEtYl5b7lXU+AGYbpWCFEIqp1Su3/tv+9G1BmnIBr0NqVt8SEC48G/dJY0soRZyJ
RTX9s0EW3GBA9fTU9u1VPEwKmFEerEgU29WfMSijHTYPRbjh+nGfxSXfKcCLGEBD
H+rs2VKIapl7AQapURqB4zIbM53WUb7bomtCsj1vp2X0ty+TJhz0JAEw6q8dRWrA
BWU3qys6xnC7hpLZnsxzwY9NnJZ0mwH51pSbLf5k0qCWhXyiEW7gqRtHicwy+odd
`pragma protect end_protected
