`timescale 1ns / 1ps

module iob_axil2iob #(
   parameter AXIL_ADDR_W = 21,           // AXI Lite address bus width in bits
   parameter AXIL_DATA_W = 21,           // AXI Lite data bus width in bits
   parameter ADDR_W      = AXIL_ADDR_W,  // IOb address bus width in bits
   parameter DATA_W      = AXIL_DATA_W   // IOb data bus width in bits
) (
   // Global signals
   `include "clk_en_rst_s_port.vs"

   // AXI4 Lite slave interface
   input  [    AXIL_ADDR_W-1:0] axil_awaddr_i,
   input  [              1-1:0] axil_awvalid_i,
   output [              1-1:0] axil_awready_o,
   input  [    AXIL_DATA_W-1:0] axil_wdata_i,
   input  [(AXIL_DATA_W/8)-1:0] axil_wstrb_i,
   input  [              1-1:0] axil_wvalid_i,
   output [              1-1:0] axil_wready_o,
   output [              2-1:0] axil_bresp_o,
   output [              1-1:0] axil_bvalid_o,
   input  [              1-1:0] axil_bready_i,
   input  [    AXIL_ADDR_W-1:0] axil_araddr_i,
   input  [              1-1:0] axil_arvalid_i,
   output [              1-1:0] axil_arready_o,
   output [    AXIL_DATA_W-1:0] axil_rdata_o,
   output [              2-1:0] axil_rresp_o,
   output [              1-1:0] axil_rvalid_o,
   input  [              1-1:0] axil_rready_i,

   // IOb master interface
   `include "iob_m_port.vs"
);

   localparam WSTRB_W = DATA_W / 8;

   wire [ADDR_W-1:0] iob_addr;
   wire              iob_addr_en;

   // COMPUTE AXIL OUTPUTS

   // write address channel
   assign axil_awready_o = iob_ready_i;

   // write channel
   assign axil_wready_o  = iob_ready_i;

   // write response
   assign axil_bresp_o   = 2'b0;
   wire axil_bvalid_nxt;

   //bvalid 
   assign axil_bvalid_nxt = (iob_valid_o & (|iob_wstrb_o)) ? iob_ready_i : (axil_bvalid_o & ~axil_bready_i);

   // read address
   assign axil_arready_o = iob_ready_i;

   // read channel
   assign axil_rresp_o = 2'b0;

   //rvalid
   assign axil_rvalid_o = iob_rvalid_i;

   //rdata
   assign axil_rdata_o = iob_rdata_i;


   // COMPUTE IOb OUTPUTS

   assign iob_valid_o = axil_awvalid_i | axil_wvalid_i | axil_arvalid_i;
   assign iob_addr_o = axil_arvalid_i ? axil_araddr_i : axil_awvalid_i ? axil_awaddr_i : iob_addr;
   assign iob_wdata_o = axil_wdata_i;
   assign iob_wstrb_o = axil_wvalid_i ? axil_wstrb_i : {WSTRB_W{1'b0}};
   assign iob_rready_o = axil_rready_i;

   assign iob_addr_en = axil_arvalid_i | axil_awvalid_i;

   iob_reg #(
      .DATA_W (1),
      .RST_VAL(0)
   ) iob_reg_bvalid (
      .clk_i (clk_i),
      .cke_i (cke_i),
      .arst_i(arst_i),
      .data_i(axil_bvalid_nxt),
      .data_o(axil_bvalid_o)
   );

   iob_reg_e #(
      .DATA_W (ADDR_W),
      .RST_VAL(0)
   ) iob_reg_addr (
      .clk_i (clk_i),
      .cke_i (cke_i),
      .arst_i(arst_i),
      .en_i  (iob_addr_en),
      .data_i(iob_addr_o),
      .data_o(iob_addr)
   );


endmodule
