
   ///*<InstanceName>*/
   input [7:0]  /*<InstanceName>*/_tdata,
   input        /*<InstanceName>*/_tvalid,
   output       /*<InstanceName>*/_tready,
   input        /*<InstanceName>*/_tlast,
