//empty file for now