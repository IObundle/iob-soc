// Data and address widths
`define GPIO_RDATA_W 32
`define GPIO_WDATA_W 32
`define GPIO_ADDR_W 2
