`timescale 1ns/1ps
`include "iob_lib.vh"
`include "UART.vh"
`include "UARTsw_reg_def.vh"

module iob_uart 
  # (//the below parameters are used in cpu if includes below
     parameter ADDR_W = `UART_ADDR_W, //NODOC Address width
     parameter DATA_W = `UART_RDATA_W, //NODOC CPU data width
     parameter WDATA_W = `UART_WDATA_W //NODOC CPU data width
     )

  (

   //CPU interface
`include "cpu_nat_s_if.vh"

   //additional inputs and outputs

   //`OUTPUT(interrupt, 1), //to be done
   `OUTPUT(txd, 1), //Serial transmit line
   `INPUT(rxd, 1), //Serial receive line
   `INPUT(cts, 1), //Clear to send; the destination is ready to receive a transmission sent by the UART
   `OUTPUT(rts, 1), //Ready to send; the UART is ready to receive a transmission from the sender.
`include "gen_if.vh"
   );

//BLOCK Register File & Holds the current configuration of the UART as well as internal parameters. Data to be sent or that has been received is stored here temporarily.
`include "UARTsw_reg.vh"
`include "UARTsw_reg_gen.vh"
   
   uart_core uart_core0 
     (
      .clk(clk),
      .rst(rst),
      .rst_soft(UART_SOFTRESET),
      .tx_en(UART_TXEN),
      .rx_en(UART_RXEN),
      .tx_ready(UART_TXREADY),
      .rx_ready(UART_RXREADY),
      .tx_data(UART_TXDATA),
      .rx_data(UART_RXDATA),
      .data_write_en(valid & |wstrb & (address == `UART_TXDATA_ADDR)),
      .data_read_en(valid & !wstrb & (address == `UART_RXDATA_ADDR)),
      .bit_duration(UART_DIV),
      .rxd(rxd),
      .txd(txd),
      .cts(cts),
      .rts(rts)
      );
   
endmodule


