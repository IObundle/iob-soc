`define UART_WAIT 0
`define UART_DIV 1
`define UART_DATAOUT 2
`define UART_RESET 3
