//add core test module in testbench

   iob_uart uart_1_tb
     (
      .clk       (clk),
      .rst       (reset),

      .valid     (),
      .address   (),
      .wdata     (),
      .wstrb     (),
      .rdata     (),
      .ready     (),

      .txd       (),
      .rxd       (),
      .rts       (),
      .cts       ()
      );
