// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dmMFKEr7wGK07V/ng6DWqmHX2gYE4ZyZt06FEpn44DXcvds+rvLI0gSLhXu5oGSk
gl5ts9L+xgDmHzMzrII66Q5UjFBRz4CH5ishU+Z5kuYQ7NqT3kyqOEpFoo7STmfC
KUMstkwHJtCmUwECO5ft3rqiL5UWkXIgQeTKT3ibup8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29216)
7HO7q4lrUN+mjP6t+PpDeIbNr2F4CqUsHfB9QdO9nZrUpqCGTt1cyv4dGzP484PE
bzcQZ/Cr8TLsYpX5ZLh7fwU8uno4UQlZqx+eDi+51eewRzPb8FzV4Ei+RxpuVTYj
yCpPNRRN0BOyDxFsPhqvVwYN0B+AFA9iDMEHiPrdiIE5gmwJhuH+0ZjnwgrKlVpM
RIyXCJCHlDcjzOhmoJtS9zpMN30KRb7CjgHFMHPT6QO1qxBNzW9R15e6eZzEubw5
/T87T7+F1Tf6h/0l6QqsNbhepL/m9qwUwZ8ScgIH7NwbAvsAqI02xEpgDwDlR0yz
f+1mHWWy+BFWaNk1S8XQm4tL5TFWA86Ta3IvCpSUbm4Ri9Ci3u0nhTohjOurN1TR
0COGgoat7fOnDyJKPrKHmiZMqygKpZClIDTlbiD8LC63brGyQmb12Cg0fSVxlcNq
CCFznGrgmgP+J4tyRVzc3bXywAEzMZqs1H7ZeaLTwJDuUndU/rBYDiufewMv/4Xj
7sxPmqSdKNJn+8F0tdgvJVq3b3jj8s74quNyHFpCiC31rioinm4NY8LaMJx7UMlp
Bxt1Vl5T0IINLhFkIyruu/9ogMQC4OCUUtVWiB2LGHe6QhOVzXx2bB9VdAHXuOiK
ufmepDh/OLF2aFNNSMMLWH/O/FHIqUnu0DaHxKhjJGFQCvOSf3qjfFmNZPAz+xL4
246PRQM37wKm60CEwX2FvxecTtQPd3o/bjvqAiRx03F1dplGI8pHr4quuxC2yb+K
zlM89bs60CcASKBgNTnSax+xnzL5tKZ5DMxF8Gc1OivZ2js9UZ13g43qKUXsqmWB
oKUGebF1doX9W3F9ZRjKqoJlYl+pU4w56iEGEbmo5Va0OSjOesi8NDaiei8mAvrp
/K9wO4cuHFT0JEV4SPdGIOqMreOwwVnP1+fBLXkkZ+Qhvp52wxB9r0uDkECo2X0S
xDlhS6KNMgfDPekiBFtX+d4/Jav2Om/hMMXoVn8vorTkgxy2Y+VW0JYzldynykg1
uL7PiAt1HfcFM3aJp19FyC7f3RlYLZYmWmxh/4Uz4dTYVSlrhzgZ/DN7ATaBSa6I
Yqlt9ktzfE5N4fVhTWgpBb5uMUIO+qX3eMPzy2rsUKk6OGbde2hnv+87I21fQvif
dgT9LBPxbV0P6iExIkDELzfzPLNu+Fr+71GxMP5hNXz2XyyxtMzHMbMT9MYayUaB
0yLBpDIfzI0l0AhTGJ3INnABLYDInXji66cBryxMVApdlOVDRV+wq/V1nBMLNoeD
9zBrO5D5QyDSjLIsCbF9f9lZCpThzka67Nfkyg7cDrkYLI5dLUsxIRQXBnvMu+Gg
GdASZ9o1nSfLiByacp6oQ9Bm/khj1vYG6KRQRYebWm05tCqohYtK0J9zE3i4yH8i
9mx18dFHUWAkD6p3nSfCcZZKuEyngZ48CsXSNmq74tmsZfSBTcH1bTbI6E/Hw65a
TiuaDjm1S6KLIN7YtRF5GWRh7DpttN9gej1uEP3p27GLCG9rux7jqKK8EgOFHhjA
jZOK4oFvxR27AEB5cvZEPTocT+b/Z2nvTMn429/R6JWosjwm1eNgxkEC6ZJwMVYB
bBXop8la6/o8b47uc2V4jtdo6KDy689UHOlQPJiyLgnaBVTiUXq/acM15R9pYPPC
ZF+4iL7jlM71EDMaa/Gk6ajDQiNs7NzZkBk263RCaISLIkHPqxGJuqtRhlXYQ0On
uXkDoljt6wOfgirFcEo4EWoKOUPFG3hgnqjQcf/tmdhxGAFG0pbGIQXgCQf0JuiJ
Tvt3ZQq+iyFdT770VanJEhXprv9xmUgd57xVi5wfxKpnwch8UyaMp1IJMJkO6RLg
MVLh1jePNGe0lEFrrie3HmAKlao1GN1jS+fS5LLDPFQi9nLTNp9EA0uNg3xK0utX
daQdLc4LPKnpvv40x4sjRouNGICpn6kUB30EKmWwMxo7Zn0oe7xG6rksjB5+RVf8
WST/2OzgCCk5ylhXVKGzJ6MrdjhVErxCgBSS7PxZ9tNgnR0xP2Z6YPwrV5t4B8Bt
DJPs2D3js1OO4L9Gsh4MH/jJ3AcTXfkirLlYWpjMPcggFZwv9oyyuydYTixT7/3V
ZkNrZLb75MQEm0zmEYHe5i0XxtLGvtlwU7SL3ymbP0SWBaqD0w+DRkpm5f5QyaB5
6/lX+UYUE1753WCW1JUTIUZ1eqXR+DaIGaf+QVDxq2yFDDvb7SpeQ79avXduQNtb
j6v3RgRsTh0eqjuvH0ZksOx6mzV0N8NDGo4OlHH9GUBsr3WZktfQt+2+VVEovGBF
uY0UyP0k3v3sAVnKY+o/iWxsUApC0BrxOL74ZIeuDJ1iRqeTg3czPU2EPw1tJi4+
w56sMeG9G9IEdSvT6+hs4aS65PJ+Fo/uBFEBg9Z+/eGdTyQJ8y1DCxh3+bvg7q2E
RJ2TWAzHPKOaGKtK01wbMVPPRRiQ4PLyLMtcz3DzMR0DTBl1GuRB/dAY2iXIQ+ba
UYdkZVDuWJ07ByAbFppntFTsfRmRDDhRJoNvtvwpr7lY/YwmwqXgsdxSYD9ncZkP
8H8IkLyo3OCTOCiHXo84cqtkA7+0Wo5n4oy7kI0/Xrpy47vIlYBd/hOBmjZDDlx7
EcRyLTJAEiD3+MR4bFr1+hUOk4CLmvMeaiqx2eXTCNTnsusuVGXUB9EsDrA4/a7J
izOSLHEs2TOnYHZf9NC0h+UTY0UGxHN7p/i5fzg3af6+vysfP0knb3CmuWBZrhlu
feZc8rPXrOBKPXCxfBXtkJsg4RF398qy6sQtp/jjK59d6j9mQ0tcU6IO1tJBrmoC
kusYuAJ7kmSE/pw9xrcpnmu+XYoj+TBInPcNineARQtqOE8QJXAhyVNrP76l1IXR
HJ9GmdDwB3EMQI5W7psIc3tuH4SnMdHXs9pSrlQDI3NzxOBQBT8UltrUVN+8ctkf
Cv4Sv/b+txwFqN6ZnF/QWgOySuVXkTZ8ffssVRYg0vZ97ZuoXCKhbP5Nq2++S4ue
U+Rz4JUPk4T70le/qVf7r7v+Z/t5CCrWPGTDxTwJP8yQnwQCF9BbNpUMLWx8WJus
Hog7BBfRtcIa4iTAsVYZtfehjw+ASnUGhqrnihtqOwK/8xzgFCXvU7aLWL5IZ6aZ
uXvsXD2FJdihRfPmBLqqX6SZPNc+xJWLLPD2bwPGEwDl5LFE4ciK3cnXGL39EZ0q
zPQegc3CFqOJsx7K68LWAWMUPRfh+TxECjK0bUlRpv4caG+fqDLZ/xYrt/GamsVI
URKFlfnp4h+tZldRG+Ibs9AUo/nbDjBNclcS81msIfL11r6pKvF1gYTq0qmxZIaV
+I1CqQptTkjS8zcuufqAla4VJQ+mq2TgACp/JJ2sL9HJQ2TCfMkw4ng7jbdda2k1
p8cd8zIV/UgmKziWPYN2xCna4r7RfszXGgjIyT2lo0aLb1KGBkjyHPNXVggPfAYS
8gt85ODkRABM6qr0IuTb+15QBiHstt284NwPJiOASiUfJbjZ4+UOI8EWtnucuAIU
Yg6fLRLSWC7lioAv5kwog6zALVnPvy8q7FOZl6/2Q2VBcsr+UiBckF7QKINRCyap
Ol4cmYf4m4Qqb0MH1Y4VR+lfJ6Kl4Gs+8wZspMVnAS3GGIAyWFpHZcZ93fZCvnGQ
qB553xKATbLsCCplxdh4qZ0L6cEK16B+VWHU0cg7FW/Vu7XNobzD9aCto25vzEN8
WyAt6GXZU996g14m319KDRP9zYUL9TC/JSSpg0urTqp58Tr3T4aQcw7t6emUbzZH
B39ra/y8Qg3lsWQPyeMDC0yzLhBSbbLxfgs37lC+ukGkQH9nz9GQ+6bYYVDVXn3L
QKGd16N1s61eIvrFE/vR1fZ3EAzNlI0Zm7juUD2MVqHHIZjYLX6OKJMNgZRi4TZm
26R3pNncyctD7mC3W7CDyxi4/ESoIOQNf10HAqGh63bRWIQ6B5XYrKc7f2qSeRMZ
mSE59C24SZ3cdK7a0yUrsS1mZAUsFXJIMFOqHmDnWbOkYrd0QUIu99spVNIdXEzE
GYJC+mvZBCVprzmIwjvSEc9wofdem46QS4Y8fzJ7uMg2sdEFbucW5IYK7CHtJyCT
m5DgDmeiq3OFqWwiGvMrTMaRQBIaitikOgsZUEuR0Ry7nbkWa0gjMRLuBENHTN/u
z6oMdWQXlz+gB1hs0OJQaREjgUpI/Uom8FxYd/w4gEzjPy1Nshzj8+iLqjtKYlZd
az2F1Yql56kXE3PgeYGl3JtNX1ADJUxz3uxGEKsNb2cKiCdTCchzX1egDnaDSaU/
ho42Rtc5EgWrZ+K2F8aqgIv6zR24Xxp5XyQpuKDsX+djyKdRENa2Z7ifLELDvhe3
ghmbcuKnAvRre5GPEV9t1fjkVtBNiPVxWoCE1EcYOjpJaIIS27uzOyEOexHbmwW0
85/79/DyT3jw9DkealMvSgFPeLKARM8yXumqkDJ96A085VaIMS1VAcHz8UgISdH7
MQM9SsxCnk/RDPOm4qHweggHn7sITExBRHzMvxn/SFoH3ZhQOL+5hv+rV1ri3m2A
Z6gS6vYvINKfoql764OrOoRdJv8bMf4m6Zxh837KQtMiXtU1hEmhfTm2fW1prXzf
61+bbt/lwxQPoAqDqPlsVWdHiCdailKIJeT04Yib7ZLkdiAU1jNyvgo/TMJcpf28
DZZ9XthzA29ZnVXnVBp7/3pd0RWbOIMtB8/CRL+Y5kvgN7B3T7x0XaIesF1N4PYn
wGIxaAex/aizUfAVxeeoLt5Bcn5IYwHLZmyAECKKNZho4fnsCueJK/QX1DXxaClX
qQWrr1fsXItOQ6CxnOVau/cPcgXHpxobclh3Ro6ojMY3mRjAiespyoiFN/4dzmU3
52nw6/MjDkkihra0XkruzXduG+QxpYmguPHVuzJMYaQbXrc1pz+Xr9t9o4UivfhJ
qTAb069P3frmE5L6glxICXzOgXqkdad52AoEdp80NMSluoFsvTGWRGxt5ZyQM9sz
f2xTCk2m9cFR79tx/bAsQrgkd4Rgx+woqNH26n1mtV2JQOI49h86W4VwFXzVLBXo
w1PJHBczXENeXbPHxIClLE+qTLU2sCJCkuepAwId/+kLZPgLjM5tJNEyc9vgh6N+
gU8v4C3xj52HjwPGp8xh1TNNwKNX2drWvZZE/q3oENsyXPAcV3Z1NjgnJ2mVxEPx
4bBRLbCxut6SJX7V1bMnlTD/MowhKeasv0qjDns19F7vVese8Uqw95K7RIdNDrmG
DI/9bTca1fg1KES/AsrgIt9cpczft7gMIjVoPqE2pdqrl2LRMx17seVwzHvg6EjL
6Z2PuZpVqFdYA/ghOo25RA1ErpdmeuS8ieTnRM7dGqYiysNciEqMyhw2jm13eYbQ
dWjPhdAXfLTVZsSGaz8Mzlun8LKKru74XUup0PXlxwybaZ6SDxHbbgPtR+yLvrMU
LBK/kH7TQ6x5kWmDrPuem5asW+nRqEoCwjj8/kS2yGzWQkUmDtWcyPZ4xCVUaygy
ZKgTeA+Pf8LSIr676v2UXiCuB4OR3EFiB0glUIFGk/gH2ZrJK43pUlnsaCzV6i5o
DgA85adM3pHfYi7YPZ6rN8bzc5QcnA0HgppEwiwTkLOmDK8Ng1HZIiOLJyFYi7EF
8B31elhMv/4iGx/tSb1GBDH/89/wveRqTQGK21nXVhtSYk0fshBT5+Y4qCwMwxtq
B9rqGDpathRBOCpbtEsUrAlylzqT5dSqWaNRXYFi1Z2qz1JWnzNFWBnqmQWUn7FB
dKQKilOpi4VxK3UwVgWh2mgmlDfKayngvLZBctES25S29gATrj8iHyyloJJXQ864
5RHS+Mx5c4c8EfFeVmTlFleAd3x7lhTM9s16okISI2vLrYufX7zc8aqf0OfhTx3t
TCDZQTA/KIQkTJu7KW29OabHEMzYx8fMiyoWfRj/IvyLRRVHF3KNu6dC1+bqbNrA
lZQ9U09bLV6ajuYj/YxlwaV+UdjYEdIww5aDGL+Ryaga2hdBo0dF6McmMb6lj5z/
g+Md0/Ot6gkCh02KIOeVv9h9hARWSnVL6SDJp52LN15zX7MiK81LkUCvtdV4cakq
fgY0bWOmOidERTdGB4OlP0BsC1RaVABqJV3M758texnughi2LwYZOmu4ylE/+xwp
mviNEqxFLVRETRspbi7QuVGJvz43bbfVFibnMQdCO97xLCXvT44AcZeEseC8b2Pj
fWmhFjElyDv9G9lUok2Ln1I+R6yFNl0pxTKqgtkx30bGeZxl72fa9uPQAc9Zlj55
DB2nmdo67KB/j0Zewjp+KCiavltBcuXPRjUrypRsrrZq6jXwMs3ti0u7cF/jgWBL
ZlC4xKcu2hZfoQ9hR0e+DSOk66iJ68ghaeWg3VP+TBzV29IKPzYVTSGZ0BeOvyy9
jciY0TgdTkJ8NBvvlpnakJXFRQtjqZOfkldD2JzCX+Snu5f+i3Pc1/dj3p3/qkFr
zJJvSXneQ8H39ULGCFODGhO/zo2IoF5GYHiOa6gAUsTErfMMDuarQiSE4uP9n/FS
Xc8PLlkW4tV+UkMusYqsibZBg1ZWsEzt7u08EJfK/5LS8/GkMjaSG7pTnAWw9yIC
y9GQ1C6LjfWYG36rlNr3BCassdJ9jZbiNws3gybwDvH78V3jd5ywpb9coQgpzTEb
yDElu+tnKR3n4qMYdE4MfA4m45FirNQEizdripCb61nzgPy4RQnHg2FfVYFPlV5m
92mbAvfcJ0nXud/ArdUDAo5cl2tTQ2n3GPGW2CkzjcW+6Pck6TRchladULH7ygNA
p+oZj2mKlh8VRMp4/2JG6p9LICbGFiaVtZO5m53er2aSfyRr2r0Dv6VjF9RqQFaS
f+h0T9oE65SdEHB+WNpc9fOsNZMC/e128n40ERZJBm1o+nI67tIwqdhKpDCgOXOi
BwO/YvxmnSQi5kAIuBi4BeHbtM0hoaQLnfPcbW+X2tbUtFEdn0PiIi5dIHUm8Cng
A7xjWANRmfPZ5ZVK77AGRda3QdPE7yRe6tucGYE7DQGKIVFC/GdGXaXfP1afXv+k
jhjnWn6p5KQXPheFiU+G5nP1U3C27t+bQfgzKCj7cfgM43fcEpc6XOxUjBMrKv8P
xiOpIAF6Gs+EQybnDRyNuHIuKMHL5JR0Cj5G7j3S0/+hzLi/+B24oK+H6Ze6ihIe
Yol2zhUzhLBaf/wj1ylCE7mQ2/+UshqEa+MQTEza/ISdY+5zPQ+UyvkzA6fQOX+t
wIQR1DNdo5IYYKJljtNX+/buftGFjOjZ+3L1kWFyT1S/Z72w6i7WYabGgZJwgv04
TdH54xwVgYvYA6bZJYYGWOi0ExvSEBSf+Jgw+peD9u+1T+HF8Lpbvzc/rJO5+fyj
i/X7SIzmtQ5tDOm6YjtPDw5Pxw1z9D7+Nx2ejrpPY/SOQYP6cO/24e/XtH5/1+tW
ajeqfrXEGAlV5yBiEOL4NNdEIEzcD0GO1Nr9LvTTBfHd/+49vU0Knm2iuDhi3Dxz
Afr5yI+h+o4TvDUEhSFHNEt88DeQY4vIdQvQsHa/qVidFYAKnPMPtwDoMYbqMhU9
6kO8LrZWvHeK4gXFkFptmHZfMoI4v5BTwoJfSkft9RMgJO6Ht4HH958my6cPzpqS
pMOKu5loJJs56xdVfCr5cRFuWNoC5Vwzb0ab70XmqQFM29RQqzn1o6vxBQxkjuxy
y2kknZF/YeODVSFoXIkahu28Lq60N7NYLmv8i1S3uxYa63BcUCT+oj2cnyE2tCJK
jeuzzdnuk9F/NPC35VPJ0yOHY8xsIYgGdKl73+D9ZA2sZ997hEhS66XwJYmqrjuI
qfqWOTCjcYolqENT9YQiTADRhGbLzvqwtqRmhT5EGKyRUbkfahfXua4UBmJl6puA
mM6hMCUhU5WJiEokhR3Sdki7JirAJU6CABA3u3KS8WyZvEfLg76GbNy/Cmb1OkH7
HY5COWba2OUDYyNVJ0lUbEbReKHi9+NSQWDLDv9pOhietjfQetoHNz7KRuVXapBe
RVn9hnAz1XqjdRAJqYR1dHLZjW5D+WQSHlpmahGAiC5bvFxbbqhw4xVDiHbbsVf3
oa4w7+XgVD3pmYFJ72M2u+9fL4FX7B/U9uxBalnWPc8BgeRhW7fRXvz1HX8EDJBi
xVMXO1O3scc5e3VySMkdOZelJnmaZwLKtXnY7yh+6vQtoqtabsosByZCQyCNfPiJ
eDMB+3teHYtVi9o5pZxF95TQMNxKBlmJX6A6TrWV25HdxRYFKK4sdhN13NlGQ0PO
x2Ma17u2exjJn7JX4me7Zffm+gMtb4hVsZMDYuU78hIpMireoL3H+EwTHF+jyS41
ZI0/B4EUsJ49yyUtzSy9fGmdyMAOO7Ii3uus92YNnEIpUxgbHn+0Ry8N1eZS4+hm
vxPS4rHJ9m2i9Td6ZTYYIKribfr2e+DpkVRDa+IFTnGtnJfxQQs6r/BtczDjq6oO
9cFZb5FxMeUrfDC6E90ygXjhiJwwVuMtSNFSrvdARIXlzCJuZJHijqyrhDye7+UU
/KbvpGTdDGxKZ782mCTU3uGgpGOYg3VJ6tKaJ3EwvHTvv6oiw8M33lUG3jEOQwDC
4H4nJagFFPSBc7BHdQXcYFU2rXZjOIBy4bF87Vjk9ekBCRcnTbbLCo7zNp4Jd7Us
YxmxsfZ0INGFVpHC1y7rw5YtvcKOmcPbZWpCASmqHAVsfAgfrcXIcvx7mrjpdYWA
1BX7+PEMXYpfsUE+pRGywpcRybOOR8NmuTP2sdb3j4V0qMupp5IWlgk3/BsOxFYT
jcFnQF2SiaBtlnt32MpsZPOxFFmnWT6FA/73I3VzJTOoT/8DXaZOmm/a5GqzFcUn
7HZTR/a+u3YcQA85rJDaaHN01j4EVKHWo44GmAgCQRqynzjVqskmgOs7Y1gxrps0
Lxj/MPuuRptAI3vPaI4Q+XVgbcxeDiHGqXcFGF5M+KNJzzVrRG37lbqF/E9MRa/F
o90yoonugRLqnYpHCePec0HbX1WYg7wyS7+pjTJtwHAdYEv+M1jvD4ij2bFR5gSk
arsPPl9gaUaUzI6XoV6BIznb2KhnDyU6a+u6irQw6AN8s2l+hJ/A+svOm1/oJNCp
lZcVVFzRPd0hKzJeBIzAs3ZiawLr9F8uCwiiZBabLo/3XlYjsc/wsjB/S2Gc3nZP
sOp2KwpoUjcXhAbNWXBBmK4ZIxdpol2KYhaXkr4B4iWLvv2nSTEGJBKJ/dpgbwPV
vRTEpoMEXdrqlrYdi/hK3McdAVFvhoKn7QMgIK57boZuFPQ8TBo75MPq7H8ITOwm
x2UXkZytlYP1QfUxjDHNClK28D2eB2yUzH+a8YLWVMgFwSl5CsLuWqp6JYjjVPah
qtIj17VrU0Fb1d69dD4j0JC7SlWimaRfUatBTTDEnZ2w90TAftqesVEvdSi+UCnR
wbzRC8p8sFPsvBQJomi6b9RuEAFnwBKAdJ135jOuH1r9oyNnVafeaM4O3wOH0Oil
Mm8lurdTyKqp57Ddp1b5E8/+LtJ2jt7FhPCUbT8wmGz1pG0j6XVIsej3PajRlTf6
HJ6niGlB638Gf0PEpPE2sk+NaAvmQ6udHBmTbDWXnDPGHx3I/RTLeNKMd+JdHWZ5
q6wyUmfzbDVvJ+OuPQtJXSzYtQb03xQO7xJx7ao0xpj5PBXWaulmimzigFHgjF8y
Fx+FCGIhQ9fnz0xJWDwLYgR6fSKPUzcqAQA31SKctg+bVnE3vlk8eEY9rh2HqcHA
gnOg0FvWHz+8fxIZbGgIaxe+xeMzPvX25/JE6iw89k9B3ajSm4P6oh6qZmCK1thJ
qh7BvZlRf2anspNWhBQ8vo6Yb34MN9mtKY/GozbA+x47ieXbNu8OqGc3J2p+CSAE
nBOQ+bqgokqYUBBauXPmjm05WJ+TnTAvfD3lUw87AXLykaCXjCivc0W0Ylz/B6UJ
Eegi6MIkM/JpQiLWXzxPov4p9TUg0lK/Rn2H5sd1K4+y2r9cFpl4LrDsjkZqaUqm
oKZm7pyynMVJJXnjj1iws757ESIbqyT7NKAFScH82maohrmi7i83Qcoy66GsIAHN
9bTG5Af+4BOdUbEpzABHl0J8UeZ4QMuXOiHnrEoIs0G8oiLgBoxz1X/5ijO/UsUN
VcfiwQuNmQgeqX1bObqPUGEm9aVTPGzeRiLiQMq2cNjTQoJyVNYYjgRgPZ7wwEd6
bENTYeOoY2Buh+FPcWttwYtKKm1VmjnLkmsI3HCoyO+fDNw1FDl1L6r1eMrFzzJx
COzA8CSJ9fZtKayQ1fgVYyVcIK/NBXw7xGCg/Y58BlNrPTMsgjJ3lesOR+kPxymu
DyB6/qFOHQFqsiA2EvFuW232NaVYxEseuv7EjEcqv2p8oigLHQeEll6h0/uaguI4
W6+kKXAL6Zke/Vqi+0YIThxfoCqleWFl+C0gRC9VQKm/deUEb/ZiH1scXBEn5jAd
VJYuVDbvjy1+a0eNSxIu7q49tewjNRAdESN3M/FDDifb747ge3H+SC6aTClzqO8f
3P0OXUfh+bd2GehJ7djd8xN1S1ZQhRT7iLiUyy3Ua+TGXXzmiDhHKpUe7qCBJyNq
eZuoy0Zf2/ErYQpGAPCYjacGYIZm5jmpw9lXP6p69Q/EM6xp21Oz8g4oOXguItka
ua4aTIA0gkm0Ez0o9oTPzwDnqFIcBa5KIVna0ctv5sF7TL2FiUlqUyIiJSFWBvCg
vcC4tmR4L45t3S+ItZmGvMRAWTf3p9CalqEQSd+BdsrbJmUVHUM8Q49gSV5rhLbV
a48qAZ4zvdRhSY0cXOCiCz9UK3Zqi+Du6ScHugfcaNRM3yT+eAGCI3hWJ1ZO7umN
BOaLPHfpyZxlk7jUtcU1KRtMi3nGhJ9WCSAbAmWtyXALQUPf5Tnf5VNLNRPXx6OQ
krIqluN9VHLo7O/ULQ+HFt2YZPaks6WA6yyKy8qxLRiTpOL7CLG8kHUVskLSsBxZ
oN187T2a+yxM313qasqvRwuMeAYgqaVi1VkJfIiJ7dxzaBjc9pgo83TtU0hIsihR
XF6hCXehiTAkQ4MouHxCB5T37egS/Tbbe/NcD2swxHP/LBYATU1VZ9XW1r4Av8Ne
tCP7gXzvcv46/2n6PtootuDgiF+aibV5N4/x9/vNcQw0FSQSJj1xUG2mitgUywj4
K+a8/+CZw76rveJXtlcxxgxrlBo1JTvUMpUgr+60zakB3XTzwqchx4cj13yen+Up
F9OI8CC6Zto3jc3Jk3+zepYj+MAkHq9oiivPPGB2V+tHkPn0f+Zfpb704f2CDNO6
zopCEQ9wHPRM/4LHfLwczBEy5Ux0/Cf48mya0LsyQ5TWJimhXdtT+nPbwPFZrwCB
8QP8A/bXZWM3JoZIbvs6qikKvga45VRoD+Utre9aE6a1IrJ2fdChtvpH4eyP2EPs
QL2AouWHOkLZYzq6RDqoEYnV3gFjq4ZKCS2r6un+Ujv5yAkYGgKNWtwaE42msEVR
6lHQzzCPXSrleXo8aVOjpLeEqPJP7IDfwiNCHC2ublmmf3RsD1dY8wYrUZekr6oW
us69uJrpAPUSNZgWp3VxLe+g6XUMO5P2FWLXYoL4zch2EMjJfZiFhKi1IoEplwZD
XvfsG0R+qjcnAMhkEZu5YbhI8mEwqSzYe1Y/G3lwPYQml9wZy3yRZXA6yLvkFIVP
fKDJI0okcLa6Mg3iFQFZcvmRWf/+YdbnyrK84TBDEXgC9FkZfLpGPNGSllYaj+/F
kn6IzWpCwilS4qaUpU5jPrcWaajpO7VreSKDnBJHqXJNOIv8F+haVwtDvSLbgOcv
2EleKPMb+6ltEkHiOBMeV+XLNBBUSx2+SNFXk2I27eFDi8gLfjgvYCi2uSdODxlV
A+A4Fy4o5hsJXjSr3EStmZZSTEzo4Aoh9pCVTbMbYT6brZGqikXjA3VFuDgq4FAt
b1y105yfb32vN4P8/K+Yi/eeGiFkwSbaT2nH8iXJT7QFAFY64sBYZzuqk3KdwlG1
+8NMtRidU5gXj/m06hIbpTth3KEfzdIZMGOBFFr0E4DFWqrY3CbpBBaUyw9IJfWK
qBj49raRo80MfkGHH4/lyfCJwgZj/xBO+SQ9UG23phL+LSiTyiLLURweo7D4FYBm
/ExTSB83a4PLu9GldmPNzU9cuigJLmHDyiLX0usanbtVTcsBHqzNB/bsmEg9//CF
Jk/t8rNdEazcbL8HAO8r/pnpbng1C/wmWJZkt3fgA5eZYB/US5KudCWe538KWvgB
H2Pt8vXPoFJGoYuaR9msK2/zGomiXRefFX62oDLHdE5O5yatlaD5g+3xNUALaHen
PXaN3Y0W/fuv+pQMywhYy7wdtax/xGmDapIuC68yZFyQOyOF9nCT0ZRjzu3FxsPU
MllfzBT9azKFH1aQabWmpTAAo4kLUaqKwh8P0CibYhRuOhsEnRk7l0Ct6Na4QkuK
qB6zaGC9XmFjhSNLN344O9APTTSKUkfEhrscyP2XoidrbL7jdLAfwupCYAEQ88wx
du4Cxno7vnxobNCeg1v50XDIIJfs9pfUcQ/8rVuOwZ5cp+MyUWuqo7deJx9zi9ES
C1cmhV+7JkTyU8CAjb6jaA/fTqTIwRan4ReufImoFdNaWbU+lh5M7l5JBRv026kt
ClPA7NsTWl1BvmxGk3nfOTdpmsGxDx3W1d2UtFAB8a2o892EVtitamd+KYhZrYbB
dEcTgJDUgYrjf5Et0ZlQLIKnxkEPrWku+NqoknVlDYv/Iej73hl3iV9GOaffSDZp
CNafaLTeTdsqS1Ofw3vase5wUeZTdBwn6v/re8qB3CS6aNhjvVSc/6rBC6WLyvos
yQCE2hxcxAw3aQU8WyAg/kWSKDQkywwb/CAjE8iboIdCg7S/NSfihYjCSwr2ZHLt
/ZugLtpvNPfxWTGQtyNnzqo3r86vbV4tRZto77Gc3iCekXnInhaD9ef9Llk1lXeH
Nze2DHhS0W9R0FAczUYGULWfUErMErGypP6eLonaKYXrW604HwUJxOdyHPk+HfZF
Sdmpy5wcAgYoEcnVUCO1soOLzmm29O/dsVYFvmECHiDG2zaCJlTAmkTcfHFPCe1X
0dOwh0+bm5qYe8nm3bBntBffRIAIfLfcl+OlEx2VAx/rTrMS2wdriJvmheiz9A6G
PZ3G8M7+9HjZhLy8TbXP3VU7c2ea6t0/dyNlcNbCX5zkZ7dqSnurkWSQezz8g4SJ
kqSVY9no97kLlBbbV8QJZm4wgn+uXn7LfJVi0nCZHI3Yonb8lfJg/NFhZlvMRoot
DOAHW3wBGQ57l21u+WrS7WH7nqOtGdt9ddyapOuytHM+F+3f9qwKfx6IuoXxll58
Gx7aSw4jQR0Y4gkv2FyLDdp8LhQk8piapHrLULnAabswZwjIq3MFMg6QabHwMs8y
X8Pu+Krk/2dNz7ISrDQkyl6v+im3SKg7pFW6YFyvl26p+ievLTHnrRJqJh6Ibi66
sXbJZbm0NncLpDtiB9R9clk6ZyoOapdsB78ztIvEwV+W5z6uzg3H3L8AGyDycOT5
r3bRTMNVtFGbrZTIhX1sF4x+ojT3MZ9+UYt4yUpguYVryZXSX2JCGcvtB+81FVuR
RbI98nyjImu0kASSgdArLGYB9FG7FOZ41MQ7QOg/yXvbYLrS7UWjJ/LaCa4g+KWT
+KDEFGm/pjOB1sXN5uqMPOrRc2BF1okGb/I3BkWlKJKjV9QfG3eWYhfZIPglRwgb
H8L+KyzyCMGm/K4Q26AYywBq3qAdjMf/85qTuI+o7QseUBmfI1ro/+MJdZZ6/xpF
G7WXrD+2vWyLYeDpdUQR3LDNGT/tMZTdkMgoG/ahpmJLRDmcomOZCxQdcp6TB0j/
BCxs5YhvGV2OhYZeRGd1fb2K8g2Q5cxuuxA6eEVzAmA/oVUmm+1fYs1hCyDft9bv
tdBAm1SCIIWny6VFwsCFWiXR5b1flVY2Ldg1fJ4RApeO4AXSP8OYY6ApOxCBJT8T
6rU8dEhiXVdWhK2JpXpGIUZA+B78FNQVUamcUz0DtS+0PvpenX7nCLJkQiRN4L8F
UMKhGLAxvNISKj7MtxE2Wjs3peuWGfKH5aszHVHTDj4I/nQhtCQ/1Sjn9Sdg4Mee
C1IHIgtnVGKOHDite/dW8Hwj058/kVrAb4kiyde1/aznX4NqbazhgW7q1Z+9QG4P
8GZBAYu/2zdbVlGqvz1SzpJhGyczi5lOVHuxNPAjLpY3hyuVjKB8H2//5yWC+OYu
COhH9aOvhmeO92ftt/p+jV/MR9gVDF8MTMSHEIb9Qw/xXuhNgreXnI7TKj5S+6PV
AuczYrP37HeKD8qNnU+Jse+cIfhjnvSZ7/s5uno+3X72z/EjMIkTEGSKHs5HtJXy
o/HZustQ+SF/DxZXM1c6vQ7tmVKp06tMFeRtvVcUshimNvbTcHSLS+5GrxJS3fzI
EGdqpCTp0TKR+gr57WZaIulOuka4NT3oddNswjs1yC8oDInky9t+yirY+ZJTlDVJ
BQqai4wxlTjgoOiLTvkZbbeht8zeWDtASbqjR/sA4k2IHKekCxflsFSMPoIaiKnt
rj8x0bbHhutf9S7VUmLfMylm3aw/bDrFBmwD6+0qitSN23jEDc44XKPBiTLvc7W/
pQgLQm5F6AQ7yz3kLUvTEqIB8VyLihAm491XqhWoOh77eA4e4dH3cEl8W9TxCZmE
V+Nmthh8rqxOJv67/Pb++uH0SQoeDW7poCEfg7OqyDHn2gAgVg01+jAH+QsRS1vA
svzdi0C9SINsO5NhSBgLuPX/Lw5JoWhVO+DMQF3OqUG/fC2OHZ0VgMkzz+dPwZWy
ODYFkyBOUXIXoJKodBs4yRagfy2N2dzaXNkkNr7bfa4wR7jZUO3kto1SWvxWnZu8
winnPxt0vzViIUkw+mFQbnBvlPW660wq6IkqYbsjATQ1VefRFBzGLeHp6oK14OYt
lgerhbhJRh406blg6qmVOuoBeOdwBI2aL3t78zQ/1zj2ZI0SBVDmuIEwk88Wfgap
FXpDxKhw4IKAuqLjt+k3yJ6PNJyeAFA20E6pCnsuPbZWPimHIO3GxDFVuldkROUj
fElRDry917w9ZlhepxaV9lLSD7LzrYHwNZKOM4IeuHMDX406gmqCu6/A2eBDXDbp
k4UJLgcMdnRPf0tL8T8WtbdGO+C+ijbqV+z73qpKYhxJHyW/lrDeSCxKStD7+bDZ
ynzi9FFOCakfaemSJ5haJ9kN7jxceGydEVF9GM1o+1jVUz2kmQDngH9R9guHKEDw
F9C4UvncdgHZlUUeMTJySG1HG5gF2XAWPnmTpN3ucTsoQDCm7qmG0PTTjzkbULV/
7EzwZTjltPltSdkDFrmo5awKJvFkXjJLGaIYNu2UcfC1QQUMNcLOLLkXSsmZ7BZr
XCzqb0rTtfnon5I5H0Esbf9DwjEaEYTIgMwB5kLCld94c8vIhM9VKQuWcp4T01Hk
jZ8HE7UmzD3anhZOgNY1NhqFfDjV7ZnHlhUWN6UsG4+4458va/vWLEevdxUI6M9S
pQZiLQppJluhbrj1JMEakBsopS4u2uuWWPXM1f97+lh7VWwc8uASD8BdV44ClZ23
7AAfdLobRzXYbjcFURnDf5yT6QhqEVY5OUlLgcTLZL19NJCZu6XkhZfi7Ja2+Ig5
hFOMb+cmpz/5ixJl0KCwwdbywhGjaYzR4NhjqHsSqIWyW22C4CNNWadFInIuORmY
BuUmj7Jyq+DxP/+vy+G4jgOqOXMZmlun90l+uwhHN5YF9LPSJgxbhq+MFf/BP78v
IjmSk/CC8S0MjU2No21OlZsVviniqrAwmX2UFImcQgmycsY2Lz9+hEnIq7yWCkkk
EP6PSpgZ6z+daJiJNniBWid49sKhYSADnKWw+dmeLMDPRc82PqJVOpG6blW6Umwm
1GwgPcUWqkqOCLz8Vur6sFFvfKgJe4d4AbM0kh1vOY8E3g5NaLB7D3A6oPlndf2I
QhScg+gsHh5zgjRrVy/TC1NCeVUMwtQWuOVN/4BgpDSoE5YrqXC+xvbvMWWUPy6c
lk8PqKhY8xR0gICVgcXu/UZ/TfOpluOUmi9ChjAyfrJ1HD6o7GXwjaIpY3zeCRcB
pDZAL4m/CDoCDH9QXgmTtm1Jm4D3bfoIG9YYdpXjABB9lcGGvcoNRdVC6eClYyX9
pm9JWkcoqFKd5SzwVxQaoRW81SGCboGja+L6CkSm6z+qDepQ2vhqp8WS7LEWxRzC
UmIfIP9HQNKlkRyYgQRo0EolXKLsZXH6i+ZVKLJPyP/2oXG5oi2xoE9B4oWF0jVO
2CPwYpKaLUnxCtslSL2qAZCJx5k62/TFZDwX2O7tGZtAetpnk10pBLuFtbdKZBWA
q70UUyah9R7+RHGRMwOmNgQZCxmEpr0vdwIerOnv2iN8GILL3WiOfQX0BT9vmG8v
kixWQuULD5lUaOrwMZNYUKlvP4g8z5xIzp17pUDIh+5SQYALRvGGKmDnuvAAWB+D
Y4LaKOKrq42VPk5gXYMzVu7yIughR3QlAuvxjm1abWvvnUQH0RsFJCqWuAIlGccA
6srRddpqehiY01R4pH02Oa+/EjhQmkekGsOjpGXw6a3DNAxX3Hgt5KL+aY7QYM9M
f0XfmtXgtv0CBDnlmqWiaBGrhDVs3Fuia7fXPDQYp4visjIYGa0kJzB4e/bv+Ht6
PW3brXLBqw9HO+WK4x7e4/vLh7P9K1d34ndk7Se0ms9PZKTuh9x2ZBPW06VR1IlR
HSP4ecDXjbVyoN6ZdgbA1eTTlX6kJKIJ3evmTQ3giVwTxL0fQuVNUhBl9464acv+
aiqqaF1AZ62OhVcPR7VzuOSv79CpSey3o8Nxx1qRwv5DSVZR8naN0qfjkYjGBt6G
SjVu6ljfwwzlpswpZrAzBUw1zwIwHfE1MXXgkTnCGR73LCpFGCCWyTnHb5QBDlKb
ia6wGWyL4N9bX/3A8dLzUVkjQSHpyOU+L7t6Smw1rzisEVFlboJ9ur+oJjX0zXOt
yBWbmN4ExWAl4RIUjMO7FI79yX1BxAZp7FLywlKZ2Aw2F1zjLydy5YbMQvLvEFxO
cIZsgoVCnF7+shKeyet8WsAPDoLoGAmrHt2IGh/svBum7U+nXdXjVUVWGFQKvU0N
3y25/Wnv41sCfeP+OBasuLzar68U48/H/blCAdiy6Dq+YJQ9BOzESqpT3o6iIftU
e65vv8/DsCdZTImgCJfhRO7vcrlK8jIub6o+OgZ89O8dGVUc7vYlqDPaqdHKRNm2
Lp17ct/VxakDOIqrxJIJCm7Ae0484gtilzTuW4erqm/YqaX2cI5Z/C3XHSwQ568f
sl9JYVPFLmr4ekbPDyo3s/okDLl9b97pxueNikpMR2ddSwUxMhtT/3LtzmWiex90
vBCUhim8JvQumB0wD4d3b/jI58H0G3g7L4mzDuTX3/2vHuQP6u2ibj91yohaoF3G
cTyAz7LQ8kXUzz1uIUNNSlcbOoyvxlxwqlafdPxl2tgOsAiokl1NPGFreX3wCa7O
O2XueAlbIAbi3BNn9AdVV4joz4sBQ0zKrI1mYWMRYba5wbjegPWgQIXVb8VZeKNP
awQDHuoQ3ZFRdiYZ+69KSSgmfBiksqfjDMc/H0sVkeLUe0pEkKIw40vsrx1XcX3I
GHRtAvRcUsPD0Xh63MwCNXRIYVA7FD9d+tjFZoXMYUNxw+mFrC4iDz/W4oezMrcv
x1sMBCHfeFRJHr3vLyzDI66yiTBMQwzjp46Y/4e8bITc/FyIaROb0wltIj6jeSl1
pP1T4cY4/MhwATJ2XZiwZ5fal+VTcqIZhykvuWS9fGiY/lDuK3uHKSxhKjeA3kGy
04Z/ZaM6Sma3BaVIc82upWIZCkcFdSSlRkGVFxlPgdlpBmCit6uXb7vP0kceD6az
alvkICnzBNT/j8Z+sV1zUg2kAZba6QKzF844lUGTUveej5fudPlj0Lv0K21s0JoH
32I32BaH4UAc2E8lqxENTecA8yVpvRYDMqHCgJWFzqUzXXC1epMyd8HYWLd0wsT/
Gbu5cjL/fCFgOzbgREAt79T6GHWFH8LgdJGeuISxHoR9915jGJXyFQwoyYK0Uswf
Lpv95bGSmT0kzd3CsXpuVfKuJsQhwjpx3nbk9/kpK/ElDBSqiniV/5L37xtURG7r
ylYMEB16IyovspdN5U8xsi36Yx7NWnABxwpdeul0/34dhdESwWl18XU6eNN5LJPB
InSnW4/KExz3mScGBT8bDnPIq5WZ2Uccv4kgvFOOT2MhGYVLIneXcnbF5EUaFVIw
URRGorFSkEikzFW3wurZWngyPcfcmgcZajFMqE94PKn6VLqUuABUAF6ellskgq5W
csWAxN+VSU6PWnzeQT7PeCCe8gpv48aqcGrCaeQt0vKH4qjgGZGTqWgIQh1occec
0d57mPql0tTzSUsghvwIseteOCx4EPDhyY8Mw9FpByp5qFDPv+4MjUAab6hOej5u
WHenWgXeqnrI6K9zUqG1Zk3wYg/OXYGO/Z/6eHd0wNfsWoNGQk/2qQzW7OZUDO3W
WaYXiNy1SPYEp/90I/WXr2HK6mlxrTWOTulE/EsWqdrxbzWyXtyfTkDvkZNb+BrF
o8AhUTZmSgfKHU5aLjRFdPuoqQeDKxLdVEXmsBOE+yXDGSdDom9eiEhBrc42YrQn
twBccbdgUyn/n6J4/YDG2DL6SHOkoKPrkzslnlEwJtKv49uJXbeRkSXFeMH6cOal
7Yfe8gczU/ADjMFupGbfw7dIyWeYSpH4rFVcvL530TZLqniEln7rSHn8b3PPylQX
LZDQMR5EZs7s/K3zab2vvPNpDHNt8g0YNrkitxr7oCmuHj87nYd18BwHB+aSmHmW
Zc35EOwB/eadYue+Po/tBFkAqbGs3X4Acuj6Oz3qWfGAP1TX/KarfVBjAybnuc91
RU4+duL1JY+SFVNYnHBRPdQ5ETXb8Uy4ITc6KIfxQKuQISZqibYUx3lCF9sOUKwQ
cavF7UKtSBA3b60h6hhRiqPfx1lbX8GGphgjlOID/AUymJjfdOH6VLe/OeAF6rQZ
4NqoSN9LXWzkH++RpBpFakStXUicdPNla+Tl1NuBmfhFZhDZ/a01sh+o86wnIs2y
kD/0+4bkqWARxNqwSxuMylQgGWeD0ePd0Hgs0blKwx/SJBYFZ6tkM4bILGk/rZgY
z7XMVEtfY7KSXXO0uZ43o9WjPKnL1Zyyeuw9CsUnBexcVjGB2PMxFGyZe8pgmnzm
mjv6CdB/L3D71FYOegnbaX/pgOmCe2ZzMOjO43eUgSJqjwZuQJPr0QAQ+FG6+3+/
4GAEQXgNcHIHptX3rkotcYcqI3kmLtvXlOjTzqud3yXmsnlz9ZDBCVOxnUdpB/mZ
koWRlQdVjKzjif4XMAdUUJEG/AEimS726k/9GyKgSuOI90wwVfjdibkNzLvvMpgr
DL2FPLveQF9Yh/dqghgT5+Qcb1pTlFgeprIMpR9rR4nTS0moYT2rcmizZ3aybLAs
qYKoh9crNkU2uAeSJq70cPLw4dRhnjcVd4dP/Gt8fsQaeSSWpFnSBuMW5qp1iDNN
8MV+FCFKhWZIL+N7dDu9W7SrlTDGokaRfgQrbp56lNulcEhbJAjStkROXj/26J7W
a0rSrKBgeibAM1EJFJPEpwK5ds6u67c/8XqLQNVCwjCvCKymry6PYS8lN5qgCkPS
YFa8OUQNClF8GQcmuQvhr08jgBbmFXOj7KfS+Dd1A07P+2cbOh0YpfQvY5uxvu+f
IAQqMDU/vH+4AqJRwwNImP6ew40wY1a3WXDVaNWF0Bh2konAH0U+sdRLPAIAl895
NvfoOuYZ6s2jDBFI/yfcbVkBQ2ZCdfwoL/pL3wlz6skosON/91sWGiZzVpXRxBKx
hE5WQ/nTImfxy6WEji7KnTTU1XDKeX1sswJZcBjnwPv0bhW4nGAZdsfwHI9C3dMT
v4b1R7/8akuk3eyBMmpAHpmLqrVQm4hwvf+U4WLsUykLLJPf85TrfNysSwIUpTWY
huK6Dmjoyvfs8P4lJfJvilSVZW04kqm9npz/Q0RBEtPBqPkLzD/42xAkl07J7lSy
ByATNyrOcNqs6w4TMMOfWd5nxoDSRnM9vOCpBVn5j1mPznUOHx1i2CjYQfhw18ZR
G5VLtqyS1UZXTJNM/1nChW/64XkbAD9fSqLWZud+Hzcf2Z0sNXKDXgWA7F2OM4b+
ihV+qSicxeSyGmsckf+Pc/JnUJpfc3YoAvZLuX+rRdUgFlfsm5/omxkUTX0l4to3
Us/Hx8rSoZ9F25InNI3z4+UH6p/sOtmw9Wrtao1fBwZLXBnxSQcv4I9A7yotrtsz
Acpn3IqQ0Cr9d+IBCEMWC+Z6OxUU+zCZAlpsuUGsJApr80E6iAG6jHYZvkkQChUz
Ht2ebPbP87OQpZTipyYT8UPVuCLDP35GeCMTs/2nLPF43RR5SiTpZt7N06QSyjFf
BNDFU2wVlvQi7epOmEx+ZuSJqox19/2vOW23xSWHGw8yrU6EEXH8PmQ5nxsgf5/+
JqXwhito6HnmWPQ1kNqX37Iw/vJ+Ekva54dH93iDfdCFr8Yyl+LoQD1HL3ptAngG
K1yAhTjNOx65MuCKdBwlt4WNUp8iBDrA+hqyXp+iFdfeqIm+PVRgQHwd5Ve+QIcq
czWZg9AznyiAC+OpeXDZIWhnFkrCxzq34dqNvJsGnOXK+UEPFqsvoZ9GV+vHGkKq
24dxG06MsGF4geyGJQc2ADw2vmG5iJDMDPa0OMfbBweWwUhIq1a/9LP/cqC5+l1v
GY9e2MUyzKu22Na1kzrR+upORkNzaF0X0ZWZlAziMqe946755XAxg3Z2RhwXjr26
9/GxMxx0dFINc3bI40/z+JvdFaHkLf/iooNjWYKOPL+T+qR4fFkznQHBRmLUsxCz
p/QOdBd3iw2ARM5UBJCEEDN74XuqKb/RtkbJ0tTIAmv84wy5CB2gx34kIV2YksFk
OVn9vjKhkkNMJ4iy4V9L1+t1B7VKMBExv3Ta9mMWw9Goyi8+WDUIxH8DVfsIjxCH
1UkyFYvecJAC4OV7gt8cB2da0AWx98nsGjsZ/lSimSnJ/WPIVAVaGyd28bPsJ38T
Jw8c+M2VsDbQN6RyC6ja2/Be4Nx7hZb3JTiYWrhJD8Ek8gAAj8kFcDcJa0w65R3z
tyoGE4doqZfRr2b6wdu1jAnZVU5YrJuvQr8ZIq3s/fJc5gty6RDc8gH/gGR6rhtJ
Q6osP68xGihoH1ualB9jmnWhBrHztMFF2P8s+6/wEF1DIaIi21X2l51/+mlHbKXT
6diuoFyuX4xhybrXHJgplRV+gLLaV8NRYi/lS95RmVIf32lWGFINcyIX97iMVpvQ
ZpIboHsyXqfHYRc39EwnpvXEUbVH/TY/59lhEelk2SqMFjGsx1ISSHwuxu0njyHP
spKjXWkEACARDrCqhLrqzDcl3EB8g+nB3D9y9GLd3zcash8crGFU6ImYpLI8mn1K
KD7V220um9k4VkGfBBEihulu4gMTW6S4e+GKXAYQIbkQdHdagVN/TOdgjQmUhENZ
xdN7X3c2KB0RD6H7jR87ucZkmMpEigNnEpETW3D99QLXQ6ZPS45MKDVB5zMC17MI
r4AQeeOnI4ityhzW/GFkE+YvkA/lur07tJg2ux2mDWrIgPhB7Ok9BOElLiE/RrnC
hxM51ksYMT7gq/r05woHkxip0Ral74jH9tCTxyxKJPSjGos7qFicmFjbUVZWmEAS
0GcLaqzFt34+7WnEJLfcCtGw9JAH/SGI4EwMM7X4tdERCWb+eN4uIKlf176LyUkE
yEwzOrUmrLmkEhgcBLG03CYdy2nBS+Ud+Ai4jXrNSiUgud8XDizLJZLplFZHGVbQ
vatENcxPD6WrrrnAalcI6/igY72wpd2wXn+k+BU0uj4tMq0JdpHROBYELSB1HJ8Y
rPcq+PQB6E2Tbao4tk6mzKQeMgSU6Gz9YB7Wxb7aZwiGareHw3ijqLVxNSdmFHHM
WzHMaVAPUFU590/gOs+7fJvqQyF7RR9SLgwQzuV9IpILZ/o8GAPTUy5KYjs4Kt2o
YSNze0SW2Q7F0ZjJHyHZ5SBk/7MPjmb3KbEPhQBVho5wX7GamB0PhU6dajymnLaW
FCPqsRSrv5JDNwEO1ykCNmFik+wkDzOR5oGjjF+qraxM94qq7LWs+8ZauzapR8MY
ZWHkvO20gudlRpAKo5/Q1gJ1ixNe9rrWvf/+EggzQXSxBbGUgRJ0rG7DIOBa1cqx
FBWxhktgg2E2iTMKK7Q8H0yoG2COOYOFYpT70xOXGj1p9I3sPAoPc3DT9tYFVyTo
DdzJEuEt74T5pAv2TCV+JpaEG6ELSpMH1iFiyIcUxRDxcufHqrbWXd8+1NDMWozo
/R3pVXmVbxp/qMBEIzR420AfdQ+KgtAMhLAxHIq0uy/6tnq2BIEvIKJQc82uwdwI
xlaqRMr2T3hbjlhq1yttkqKo6YNbny/xQoUhWXMuX+Q/sR9wufSrb9GQIBNU9+Mq
Ua0z6g3URzUFNXIv2ZKuZMx+c/pd4wUvw958mFXgaakWG9hd2SLLe/scXnLPMdM8
O9E/7zccEOlKXGPesY4MKAYlhd7r4e1zKTW0CTyP9j00NQzzFQO1QWbLO+Lka5kJ
ogh9Cvbxxz4OHmEjCY8lQB0hrjjD2LcJluLMZ8tleAOe7kyeOGywpQ5w/7PPKz2r
D4roplBpuMXdU7Ps6jQzBZi6yd9QgME8cLDFajNZ7Zziy8K18O8lTmPz1on3Uezx
b2+9B2YnuQiv1Qggz1fnf3yMySE5SG9QMinFpOw28KvTpZt9kvuiCq1eHV/bVLiu
YNr0ADYnziaYWDKybEobaj+fL2aWtxKk523nRyb4Q1yFCTAxC7LHZaj7wzdvMaq2
f41zK7C+veJY392TkrpfS2IEPav3LM6lPpriKI+eTmECfmfonYepcBQ0O77f7CdF
DHXr7uuMb2im4TNC7kOt9IhGwC2liu6n8Yh5bb6V/vu1ji2usjOoZ3A6poq+6qDw
RhHqxZ4vxPwbbKHZZ8ww8yXbbNscKaakagMDxUEgn/RxM+PQ1XbO3u88ZI5M8h07
fHQfoTnjhCftwMVizCnJnqXLTe2J5xevHXPJLxYHfm5K+lZgCwpiS40JS3IfZBqi
G1u4CGhzAIUGpQJ0Z0YixMCO0/Pjg04Svgfjb/oA9O7kJ6rC6bftr38pqSqdtrhC
aF5pDLc+U9u5nP/L1LDtowY+x4ks1bM3dEKZ5yle6CLepCqBxYtft0M+3N7KeZiR
8M71b7e1hOZ/O5fkg5mbEv2pZ1rUbA1N8MKCTFlzVSz85vdWBnhiTMkZ7A+Ksies
9Cr3dW3L8PASlEIDCOHnwr3/hjGJ7Y+ICDCM2MP1uwoT6nYP6kIzveDvGV4r43Fz
PzVaYziXyQyMUBwF/skhngwZVAfd2aQd/hJGbcI4ppxzsGPNTgODvF9Cwx8kBScS
IUtUobTIG8LidEZSfRqOmrhTOS45+k/gl3++pbfVtcDR+ongdDpchbJ97gnpOonS
0syh2ZuS+MPtjcvU7WADJ+7jbxwd0anMeN4lSMafiTaSVVJncCNzvKoCU/GN3STd
FEjs+PLzrwKbQ/MtcDk1hVzV9HIuz69RL5LeSMIK/RGf4mK9KgBIlcH7xjXAa/Ei
fMeuK7HmWUz+ETDelR2Du31Z5SfumhzYs/DajHnc0UOLF9kjCOmvfa8wX4OBz1Oy
yZo4mbsM4nmOw1c1aD4yoWB6CcEqBHxNvCRPytzHIJHaci1MWWpaYlveE4ss5fzT
5rkV2KUD18BBLK4ImaG/86Le5qB5IgdjOB5fE+WfO5SYrqQmSY6oFHv7oEUGQHAq
Fpz6jkOApCgP67izLzvyJmYTQfEXGrCrC30gxpWUucEVVngWTPtj7L9wka5oziS7
kAroT14Mm5qbeOMd2ZdTiCZad5j8f9TZx4Cb6Xz6ppH8KObMNk3GMcF1dlX2xZcn
BIdl+CGHFzqAV4GPMuzHqH1xMR12LIvw6nSSFRB9WJkN//AOVeaT1lAicxsx5SJK
kJu9TiBzAFBmxR6GRt8XakhMbJigG+D8nufxbl6EsjxLzGzfjOU84D04US7xGpQb
6m7QsNkuKMPt7pbRSTzKFkc7YK3LQ4uM1QqhNC2WjM6X5SmF6FY3ru/GcdYXMQvI
OmjQTpvXuHqromktD2Ahzbv8vTwhWeQMEDlX9SbOggFLEDg1vud7d7lz4Antf5IE
53QOWoo9G4ubbeCDXsstByBA0TQMXww+P3G07HO19T71L0MJbEH2/8OH/3Pwrvb3
1stJrAy2Qz9G52WmMC42qJQmHcTEbnpanQmyB1EjU3K764gdZHO1yV0Q2tqmlK0Q
xRBfmW4bDs7dlmevvGBDbJCv915My0ueIoxOpjTw35x+PtOU2xu8cVNtxKaC51vQ
l+Jnk68NI82EMb+8WZkMoliG9d3HvEuTdJrpgM14++Re1k3y8r5lOnws60M/WFQz
3bwWY0BvaMhJTiDUFH7QYkDJ0L0IWD50i8xOIA3WdPnjJd5kV7IX1rhMak7Nc62N
kHlUD74BjUN47SQqKy9FHK65DKrThBwXPqjtoYKXF5or167J/et9GF+1Ty2krAV4
f15qR+fjILfMNfJJvhDNnBK7oU3K33CRv0rce4sVw/rAKRVXAcrx8hjSMwSjSJNp
Q2iLKdQPms00Q03TbSnXxCYhbpaAOEzQVa3dTA6xbOsmSWiI+WtIRilc95DxtTh0
YcEryaqx1qnBEqbwHdjMiMnhkxY4CN2p4EQCwPXXRYRvnJ7wvuylH3sEAUjXNzZs
rkAQ2Ziwo8jmXAia0YJ/LelqLL/ee5eMvFkw33p7Y+uQ9X9WqpcVxYV6/FyDSnpS
euxAI+IbEc9DzmF3sN/7+Ri6BNQu4qsOHlguEnACZalihw0eOWMWIsuRzO5VaoFA
dI38T9BPOUqVLXTZzsg2t8ctatlLWkRCcYqUSTdcH++qe2s1gfDqViZEf64KODSN
AOIGWT3TXT09pq/hcDoEUqviOPvRkc8hXskar8TxPCYiek0N1IgYrvZrSR5th5P0
nY/MC9l0wIa6p2Dr/pzRtGJTb04iVB6BhbvtRanp60b/GATNpF8KDTlGinMW8e57
ECh6XjiFh7Tjx/NHF1ZIVP08ShSJKQe+qWt/HF9GUJ3TsAMiqN21N2LrBz9bch0K
AyIgXSokt8pp7WWFiPsEp7WThK0CcLvCzK8BnQradLzCmyydSHiT3tB7wqiFz/3K
6v5m92JoT3VBv9HSb8jMelEIDFLsdUO6VIF6B+aSfpDNzHpqoRCi4rsRbflo61Ax
TpGh4WQ2gPwWNomt/U8sTx1ti5O6YD9NiLeYZkQThb7JbAuunNZxqjZbpTmgNpi7
zeF7+k9ukGZ3mPS0WtrH2f9HjYLk7sRX3DFjDVHrJM3FI0Q2vMPuqQ/pV61Zdz3S
VnBtpcE9tEzsYw9jIBb/f49Ct+v4iJRP4YzzGaLjK8wujJf+qMjJAykWIzbDDIH9
HRfM6kdAYhycPs7lf1l78XGqo7dL2vz3RZkk5DuFf9rES22Fg6mToP8FIRBwDkdn
htob/2JmfpaURbzsjrqzCTakir3k0Z57Hf4FpOF4hsNIEwZCYMWIG6+Lc9mhWwYr
IrdzYkHAgXylm81ZLtpkCcmQVRc4edbsZiuUWz2kLz/X/wt4ZaYdLzLe3T5DBLSK
LpFWsIyFBSEGfMPKbAJP2BIc/KLyHda/bbiw/lrR+TDRBF+pf2dLu9RJ5tdabxLp
6ysNi75U7RsQjWp7GZbUG2ytkQJJKwbzE2DmQQuH4SwYDz9morSuI31DjSZmrnP8
e9b2y2ViPudHIZ0sN739K2iC1Tr9FUBdN5ek7qUOZZ2zNlchIQTPyl8Dc3p40FWy
GI7HejNPLwR54qEhjNJfbQ0cfMd6nazaYQLjzC5vKcZwC5vmbsUyJpfEmP6s7MXg
LlyuY6i6SBthfhJJRTfnRHNV4Q3Ca5HHfoD566mM7sDDu7vlUEyPMjhO1LdHWZai
AcfY2lzbC9pqy5aNUnGFVL7+QNzDjiDoyCcWXyCmSsupYYiQTsmLynxzk3ghdwjO
3JO+e1qs6j7NoHasZKH9OzLsbJjfC23C1pdpAtyRmXEmRRUkEXljKI99AUqgP5M+
pHDxp3qDwyCXML2flMyIPsopM2IDmRjOhrhyCnUoKH+kK2LzW7NJ4L1+pcrBen25
kosm12Thad6mMJHxBFPcqzy3HHz3HqdzHE5xRzkfT5MOWgmnVYyk/jcucZLFxuv3
/saYmT7EG5aBbFy3SNvbPafW3N+aKl7wvrnLvQQPsUpdEyW/jciAyXudIe98muFj
Txny53aG+K8Uy77KjV1ewTpsx/PVeLFwZZo7qPNzmCCqeah6JTWmc0FXjegBbaQk
6VdAL4lFkPi7D4jWlVNu98zoSGhXbOwazjNuPo8w8YSIWiC9JkRYgpvlCEXI4sw+
uDN4h0rgaptVX3t/gh+3tsFLpegRfI8uoONUA7lLxI1XrwCMbH2hOcWE0tuGXAAt
Oc7/I+AaV+JfsVXgrblRDjWPzJ0BlhTyR/6HEuDQ2E4GjkrfBQEOYKE+6b+daZAx
eXQei2KALCzcAEoUC39gy6zPBaOliwXPm+rJgkzl3DczKYZ/Win9e0msBGFPrK2/
wE/uzgZbKTJ7fFL8T8dpbIEdaUU5/Iwp4xNqcSaSc3MedH870evinRtguM9yojpa
KNnkx+DD/U1Df0hVetiHv/kWug+SP7VcumbvKHdnMHfwKsvItTyJpENXQvn6k26b
GXYeA4Vm1PL+5a2a8Ok96kWCAJLRbme/CX874wuWYBGdm1OqUQgEvbaHt/xy96/D
b7dVGYVMK5KJoOpqJccXFJ9ie9V4Y/vyHHypIna3NLcgCQ7LS3PTC7J6kWQABto5
fi6Gw/TvwYAIbDNsj8+fHGuf4Ph/nFNV5wbFHa5ncIT9On4O1Rzhn1w5EaCLyQyB
sksZc9XVioFXiimEnTmBk2tcqfgTLbNRVSYLEM+3uJmE7qM/zQ0k2WFxYVv+18gG
X/sTVHywELNZ38IPkIiqGxa5tPSMhAr8NvIPusq5Or6tjokpLfrtrhcWOA/kubMQ
8FKxlCSCUc1hejQ16Q15EthdhxwMXGHJrlYnLk55RccWtKSEIJDdRBrQ0wG14/Ht
I4rb6Z4mepLpAz8cLnuTJpuVl8JcBSEMLv1bP/Zfn1kKaqYzNNEbo0fS96ssTCk7
EmksjO9ryd4+GBD1YhIrKY44w1mUK5AjVUupXo3wiMBrEKSQlM0jgPZedeNJ7HWz
QVRgHusSaSMcXWod4Fg9HetcPxYQflksfeDSKr4hpSqGV24knFiYz2ZKTJ+yf2M8
zZiunyymf1J1fMLWlaBXGoiA54E6Gb08dADoW8c1za8XyNKsmnIgWtEnf3A78Hoh
3Q6tbof13vdh0aE2FEDDTjcKFIanCWRWYeYTEMixo/OLSaMJ8+VE2/Z3D6SdgrkS
8f5mAwgbXLiGC4s6cSeBIl4+frVDMDBt1+Os1XQZ2GprR2D9C4QIKDJgzem1vkKQ
KCV2ZZOSQJtFsezkmyRSLcJQx3XdjkO6Cir0ujjrvsu8x+8d8+1ijkdJuWRHRR4C
Dc8ptkqV5pnGID355hfy+MpQT00scG9+r3loPeH5Bfcg49qn0DYFJTywwYmwiELU
viXlR7j9f3XVm4gJW+dRc4d5Dt0b4DCWMwNCGMlBa4lKEaFk6orudENMMPu/oFHK
mW3W/zT172UBJpt8buNtndVD2OBsL8Dq9NHMDa9M3TO508abt81o2Wdzy9Ji7cve
OzZ0Mc7LA/DoosG4p8bu7KeLVWDr8R8XTlyuCh/X2ZB8mEa1wmlAYJ68TJJFkDCo
Awrz3c55HZHE0CX6DAURh2WVg/4p10xBDR+0l2BBTCJ+c8LSY3GYObbNyDjNauOt
neC6Fdtg+1NvNrvPlIBedGwHrkFOwctw6VLn4ZX1rvooyCQvhbVm6XRd5+qy9f7u
VjB6Cu/pD71QAbLEWVeGfcwaztygRGTjQ3RUDPCmCcq0bbk1+860lQ+gM+/34KfT
mSv38icsj7gYkG/obVFdnMV5Q5CSzAe9EUo/1ajdq42hfe6s5/vAYGebBPjWDFPB
Da0yW7c5PPSvVT2+e4LG8RlcAG8HQpiwwrcYUglWxqXOk1AICK0cleN2OnePgHci
20yapvu3qC0reVLywQSOG+ls2t5zjfjbWQAIIzQFFez0YK9Uzw4Noa/FACflQxDJ
87BpQm0C20EfKdD01IrlIep+PefCPeyrkpCEJv/sby02sHBp4a+Gu3aDhrWqMH73
vhmSHtmBIkQdPqr2qQRWUyCPYhKDf5Q2QuUUyhPVJaq0LreJchbkzxHjVUcXtnbD
bpht0Bo9PrsEnl+r5pnq5Bc5T3ECpu+f+hFnmrCUglCzhl8KFQQjxdBGdqFH92Ro
M2Tza0xZTsy2VMqn/4ZISKYBNCa67rf7a2KdRtRjPNtKoGTgo6ohb4XhsGndR3WG
rZXP5Eam6ncp2Pp2IL0we0sUxSiNRotXU6qj78rbLYCtQJVQtl90pmifC57nvwkO
mxKB9+xveZ4Tn+iFROjEM/LopeqdKWx/cINncBX4le37ji35Pgpok1dFq/1WAcCm
QenXjDr/c/PajbF5HnwPUhaannOO9Fzi3IfNuT6IB3iRGKBUmfVmrx9OACykbc6/
YIVml797mNqb4b5MnAdojuNux1BF+Tj/P2LoTmv1eOzTaOEcuXmoZmudwRoQHOOW
JqevJ0JmrlLmuJZBE+HkhDAgbyIGpOAA2cUZ62vxRjZJSFA2GvSi+xtkvhbTLTMO
meg4BeYQHQBlsxakAeb4XVfs5a5nhPEme/9HmLqYoeOKWBrCWi3LxniHQBRpucl7
q28p4LpPefb5IvnIYMjdV39Onq0jGDFUP3x3R1LlrdRFHj8HAYFfsv6ipgzb8Lol
zG3zuCaYFILCyl02pw6zjaQtgclplkNvra29JDpbWLvcIG+YKG0tV6aD9wx4FBVi
LpgrIyIRlh4TEyM3GAe2kdpwSEMo3PNWES8sAtRkhKt2hd0ZwfOrPcVIXvAUBKUz
Jz2lmgUE6fKT3m2GvllpmooIuGj5/Qj++LZAJTONpoP/jN6hBo3QCTufTVpNBOW6
J6OjLyYBGaiSmQzUoEeuqtT8IYi0zFBog5PzkKwwjIriSsIPdzWSPxz4W3LljBGF
lJjnR7dwW+7K2L7w0eFG8zAAT85WQZCB8AI+hO1dxJgKOnadwLfBukEAZoolHXw8
2ee9znD4selZINrlr6z63nHgilRBE6c/THiGPsLrJ5s36WbqhN2O6lUofZCDCef1
QJB3BY9DkWNqxESgurGvfoN1Rd+r1ryvIVdX/8bHN5QmGPZe2cknXxCQWo2k0hw+
Q2BR/3e0rykcFVHxYqKKbiTXo2bXH0gwlkcyyFPeDFrl/WE3VfEHhVQb6wibidoB
kuCAr1UdILAbbnq8wxwM2spTR0TNxymNUMitxJIS4FTkd7oc91pTRuM9zWO/+4GI
wbKFcrMZWGkPLlhm++z919wnfyQELFs8zh3aPkePLcYvfV7gxME+5k0y0WEOuubN
PBDUUmDqMoXE/m1TpAZDVBWT72clMqc31qgVDG/ERiYxbgb4tp5pn992X0nNZceJ
/ZIwGx4P9GUkKyzM41xkK/ied3ZVOchjNUlEfleRvoVCx676Sx1dG/hrhfwqg3k7
w1qeSOQ3Xf6TUt7mvuZgIlYgdNpy24rS/2z7B1BH1K41eKriZnYScXZRfQRvCNpE
8RI5H0726Zr1qm3ged8k7lgolp55ZzqS/lOW9k7z+HK+Gtn2NO3xQ+mT8ay62U+y
9VNMs+3pBj+LBN4gGJ/V1Q3TGLINNRuMsgXUsY0z/kqJQxwXmGx53k6c3LKWMUAm
LTv5KAMdECajXfkRn8hrPQZRP3sMnDN6/L5b4npYbWoBsnHVMNcOwQ6mnoccWCw6
MzDpeh5HkZj0/Nt28zuM95EZhn+XUQ6M7kzaFwWVP23+WwUmmhAMfs05xwDUHmgz
izem7vwzU5bP8Xh9VU4vmJNBc1p3av4SAdeq/F1PDkYkRuvFGxUedj8IBftVRKuu
BbcegSibKHP0nOXEXPBYeCyq/PgS6QOBOvrcZs0xuJZe1m7coVypp76B/bMJnbvr
03bMFJ4pG2FVkgpaLAVtO9+Em9AaKeNNgj5PxsYb7SyX9gjXYM/k8T7ZRqdqoCVm
ucAJo85y/b8K+ndv7e/eyeAAEZE6FfhbkHdJAkCNmyMK69Mk0MmcFiGMB0img1G9
phb9zIZTKZELcSnUjSgy37UzN8rgLkR/yaJWGMsHKn3wCCV6fgYSdJpsfrVRmGKZ
ZBn135qNj5uQqzVbwsUTbCkJNFOkx8FOX8ft/W3X/spt40XRRzHd0iDVyIa5ubou
QhZ02rMCKFY+GgoxZM1QxiR4aYtSjFKlzFTSud9OqsVfXPQt2fi+IbHvNc8z27Fr
jYCUC5hcUQibQUmAjAv9IJC1VvYVGCxVhgt7iVRAyEBymiB7n6ozMTbhQO57AXBR
DTjlNSFJcwfHDa4OklraQfELuvV42nPR0qy5VK3heS2zD4O9J7KEYnDoEZsFzyI5
beMndAGjz3NgtIYrvIJHMFOvLa5/FrLc6XQoXz0pwYjxGe9APB/6nfG1Ss+RjNze
wakx788sD7UUe1f/JLL072StxsnZLxecLTmwI+y9TSvv/hPnM1db24eIHOW/HXpj
BbKvwVjM02BUKij0calc1BXRD5lZvH8rH9UMA1uRG2yFs0V5VZ4+Bu24xdQeUGt7
/Rd54Mb57rbpoxn4KNvVLwCfn/mrRtqCZRq7SNZpVbR5XxJ1Qi0STkGm4Y+rELgF
Z2Ocgt4bX3LmYSahsmzk6YlVL7tVyYtN3NSASEcu8QY96Ui92m4TFlj7nyEsRJHq
ncX4/UPDEhxf1MgDB3O03701Zk6OiSqJSE9jJkRZkiPtHek/mqnI6RIjEqk6VOuT
ENx7ViP1twLZzuAje4AY7Yc+JOIMlJwHXMv2hICJ86/3ArGG5RP9Z8yPEJca9hfk
zoFjcGdbDFMVqAp9UtjPZpfDOBlpPpDVkFt4YeHNyLZyGH7zoxpY432Yg3HBJ1jc
c7wPq+z1Q3R7RlSCd+BrVld5DLn6oQe+C4MNfTSR6suJBLjpAegyP2KF0MSzVX1b
MtYK9WbK3KPBbpipqI77PVx26Smebkec4dDJCm4RpsqTkmjDgXnSBe8U0qmYjXKg
Gd7R35UHletlWCSr2D05W7v1oP1+Zf10zSrbKDXoPwEDase3ZCrrQQwKEVSPwpPw
fYNEGf1aa85mxAJISmhlFTjA81EoD0iAkWdqwocTRv904nR+HyXbm91vo7ff5XGl
SBJ3Z7I+lJ2hislrHw9QbZ5dLJFu4jc5F1ZMay0C90A/vZV8GEOSoqXtekA5dTW9
veLjh1XKYqlZ7m0Nj2QqwzIpVoK+5MAXe2CEAUmqJpDUahuO7Ra7cBrJdBArMIA2
a1LoVMVIzAwtqvhLA7gBRahmR5lw3H+cz1kyAl5YxVMKbxzZ/SlUOmyt6f81MzOE
WX+f7zysYliSaidnKUVC0GIG3HT1HP3Xk0cRvo8OKBx6Q3OJ+2VUE8RCMSExOxIK
Kt1LDFEZlj001oORFCzQiQ1LjMyHRY0r1hkmkZVGMOUZ7lEP4cOuxFcahPiHfNWk
A2SdBoFUuvHE9recs7Wy2cqo8I85BMEOeRQXwSG5ijufv3g0KvH0S6/tRva9kCXK
ey4pAu04JwB6sSlr4Kj4V87DOcIjYNRRNNQON2bTIw5ZqKpkSeFtH7STjP1ij9jI
s+hHYY0/3CSK+QlwBDiBjqTsbPRTYA7/EYBT+BpOoFsucM6H2FEdCyyZXjfn3fDr
Qrq5fY36nbDxo3iE+4EjViE3TV4oLLbiiVfzjZ8sd04Zf3AvtznsMQXLM9JXo3RH
o5LBvrS+bVLgRMcHdV2Zcvb5brDGh2WeF3+7uOzeUQ8v26gOCF4Orf+DJxULjIJT
Dz+xqs5nSqkkcS4mxXEuGisCxoy8z9xS+yTpJvmFCb643ZMeDL28C6czk/5aKjzT
+9Kt5ZLPQpp87o7xsbHTgAE4pyOZ/Hq4II4psVspjGqA7fpEh9QWTyQDzPyjLyt3
hOBkxc7yMunI1S1eKHYp5Pz2qeLFxyZXzfJKqQclpDEoa8EvJ2Qro9fY3ueTTGu6
Gt9/DwiD2No+qE5kbwACmmcLa80QskWBiH3Iq20W6z8JnRNB/kvcgJoDpQ0kKGzu
ipWjkCrr55CzXiMzPIy+E7m5J7uHE+VfCZOlBdryq+Gm+k6XZbgNUZ8DY7i8T8Qx
bycRhWEkO2VmNMPaB+Ro1yCvcvix9Cfus4y74VzBdnESw7JfzTHDf6solGpaqsV/
oTooVCjoHHodnPh7UdfsyrOVKgEt9BBBc/DIO+/sCLJkuXJPHgKnOdToxINTueVE
E99lsgUvTLdxRyEzdYWVIFl84d7Jy+XyHuEfZRk0LvIvkhk5bbGCFwUjovMhJgOi
qzgND3tpO3hEAvMu/xS0errl5NzyrxshlbN86i1cMf549HbHiSsbpgPj9zmr2+3F
10R3UraiW1aKqNmn8R1Ln/+PZ8YCty7My5/H+BlKbd5POM8VIlxU2L9PIif521QB
GXibGkd7E2HzgGGi7C5XU2gqO5mQ0ZNh4E8kazpN6caQ/EST3/I+QYorUlxvMqCq
7BfLnYSxwSi565cyVh8Q77HDYA3oV94IFgtQ0KR0iSvhhmuE8hqZ+kl1zRL+1yTX
vIZBNZBmZoDhAc9ImXRM79YiEmeQeTTGKRapFJ6XDJJdu2/LRUmSB97g8Ho1fyCk
w7NO8l71TTkDDcjiolDCX9bbnPlu+L+fFSc7/lpMGlNCfr9XgeJI8njnC6IEnCSi
Ws1xTeZlh/hVPMabuuxts20alu5Q8+DTgW0mMdJpLjb1JgC0k3MVKexHq+nVmlHG
d4OZI8GxWYWuy5aew76FmaPXuImt2e87jqEz22twC0gxU+kq/g+n/tmRfg6fum3W
22y1K+SoxCIv9yYyjxIWoMQM2Abh08jQxw/MfCrCP5mwEpLBv/g4d/oL7mjfk5an
qvPNR6FjG7W5a1iL9Wfu3DZy3X0DZ61nlF02y+JPnGLPudDVrOZnu5eeldHHWBQK
cUNIWXcUCdpo+iEaBAw8lREfO08dL8BtGFUGP4kkIicjQkwlUidZ8YSEjKJcpspF
1LyDJj+ZnZdofowJZ/ebhjwkotC1McyxDXlxxtVCysb6UeYKB3Sctf0jXNxGVUAh
g+6Nh6Lf7KJqxl90L8h8VFOliyU1urDf4He/TKL0Y0/OJCpnscqcsOuS4xd0thmg
P209bympY0glDtFj7s1wM2oImt8DOnPOtjrtfHe83aZ8z9HLa9OYIKENssxYcQjj
mjVmD+Ojth/6hlzGSVvaA/FygFSgj2T4CDu1DswjMYzHiKLiUCP5fXmeA4MlG7QO
aEzRG6DgVU2Tx3X66hQfCG855J2hQir3AjYtdvVN0i1aEgGhEf/+yNbR/dOjdJdm
jpipKgZXHp1htH5jjesSWhVZNNlM/gE590RFPdrg2rclge9CvfJuaYmXWlxQ0XFK
bkfFjDlRZuKBCnlZiJNaTpoxpbRilFszBVTzw1poFtfhRQQv+FIVZWmeRg3QNHYb
gM9SjEw1EdTy+TCjj4vEAW5QOibS3PuZQPSFgl/cv7xaB3f9k/8QQFuNVbMN3FBp
7HV8eNfN+EMcHztIkiKmtjntr+BQTc4UHaAlMEGQeuwGts5N+EyIBqZqTYW084en
GhpbMOWLFkpcoFd6ysmqKGeD+PbcHKHEqZFkcf5nAwAHMC0vezPWJ0l37m+xTJHE
F/McxDkwVMhCjqg8j2bl/4J94PZTd679EgJNPBDaA71xQMs0BR5LKCq+zeTO6MJH
mSff0w4AzOjpNqX8/BO5m53deO4OOeo4H1PdH5cnqESS/O67X1X4a6PdzxS10smN
piFHTxYjBX0TqO01Cs5X1BllaLmS5CFkl7QZZfTCf9ZqmS0G1DkLucujvpVvP87Q
Vhb0XPTC5/TfZ9mNxkrzOlyvxZ3EOnnkDKwXy09s6k5VUCO+fUS6/8e+3JWKoNth
Kqws/9QIo+Q0u7k5uVLohtScbJxMp5dp6WlfrKGu4xvbIN7vyRIrs9NjXTRBFF2s
vFuyz3l7wCnZohOaFSwtLKoGcCnRpToC4XHoI6Vc2+nBsVSXGP13YcGTSESgDvH4
UYRQCTiriPcvy3EIRo+TzEBwuYZ+aTQZiITds2fl3AxTjfegzAKOkn5cKo03gN+k
wx7Q8XEmvq4tdjS5c0Cv+1k6vP9Jh+H1j/2KhKYNB4nssCgOTZFL5WaRw1a7xwkT
B8OmpTgRMLY198ynJ1ErJdjemG7z7b0VcyYcb1JRzRtwnjxi366HlN9+PCM+CIsA
Dqs8GEyjx+HBwGvBH59QJSPfBQD0beHROTtBw7LoSZOoSCQYwJgEHOKs7CsoHoHM
DUUHv9dk2WZ3cSJt5lO36GjRO7j1Qa5/xFcOEmuB+16xIiR5LhCtpDtgV3KZ4+WE
DmTe1Ez2ubFXyZIVko1Xpf4naeBwrXfZSiSoOPaEtXV6vfnV+46SNxlhZkloYUwk
QOXkQ55feZgpPXsbGMOE3SS7zWIHAyDmpySJ2rkGGC1fIaHBhzbeYQVClXN9e2Qt
SQ75mIqgAs9YZtBWIIwRUT+hPeatiVgVkUIrZx4s7hMfaoQHip2THUAU3iocSkf9
u9E6IIgIyStUa9Ddu33JuEqNHymI+yp/d2ty7/ITTL6Ll1/3t5bvvipQDaG6t6Wp
ofuXu6Btc1oSlnImnID7+4K/K6rF0H573IpGmLDRGI0SaLEOcOyFTDS1a1eQJF1X
bSDCs2gXncEcAosEnAOApQ4pJ3xnbonC+BOfjSIU/bGTFSmUUt61ZfXpr60Y5pFl
/56BCSQQnTnmCCTpZyF0SIY0+CLMTcB0NthXcwWA3ocEShOUmdMhTtI+M1fXAboa
va7s1H5pvAY9fyiFYhRTQsiCsr3RvWiSb3Uh9qGK0JigusZKDGVV1znCMS3JFCpQ
ddSCBl6X7qex+F7aa8BskzU63hvLLyeoGBgr53u7SdnrX5v/0WhzzP9rRKc7d7Nx
adXRvBY2BfnYSbeYQNxXHXFND4k7Jeaxa1gOBl88PP0AHVXf8P90foVEVHplXQsL
tviXyxYsv1BNsQon85/PWhBtzInSRAfrNBWkl7RgKnsckJy8SrsIhb6PAIRq0TZJ
NSpEMhwar9C0T2vUotbd9eLRdySamT4tWjhm9hREI0dRobMBrGc0PXvvUfg3SRaR
UEqj2Xz/02RUkbczEJ3739tLQLUwYZfRNxYCPv23E35VEI3hB3VzM470Ccqlp17s
SkfQSkTv1+FARrw7uWiK3S1x/ml6YAKvNkkLm+UnjhdzQTvAFTyQtw2aOqN38Clq
Stxrwn+MQmMntvNyUkZgX0nc9C6PiEHyz577MF8qIiW91vQv3nd6Wf9eRcWYEjmd
dUHx4KVnCNk9Rxk9NVqBSixhw3RPacZTKlE8SAz3oXcNR1vB58/RGMWuB6YnF6fK
kQjh8x65IrwxtkKRHVSth1FzP7W1Uf6iqAsEILF0r+Z5pd5UvFQJy8XYVYHszXnL
5mbI333y/hUqa4nm7ldYttvw5jNdpa3y2xliF2ZcEfnBJRqAicfZJ44J3itbLqOw
hTtfqsXD6HyMFNSbDzO/7urYBl4ko7cPgVsTk/YVZIuDbOutos7q6k9hdK5n+pYK
25VKPRgNVknbcYooxvEWcs6+lJvGyFZG9k0H2GGBMaakE0L/EpRCUM2ryfElWkv7
DDEnINOccit6Lv5CfiL8YipRuV4nt5pOeZBd83o70UC8BQkAPDxZ0KF9YNvmj+aA
Jfvro7yIAWv2/8iYyDCdiXAknbIpNqrB/wpBn8FMu/ThP6ef4uD+s6mZE6h2Xoyj
RhujZTELrFOr5nwNNuwLjicxcfACvyN8+kKkNJNvkKYAKHOUrj3R76cyqXmMwFnV
nAI7JjC6UiWPiTtEkiYD0mzW2CuHDgxzLjkoPbn8AVASLNXE+0nMjCT1LPcEUNSO
aNQnbNyzyD/FfuQJz4jCL9evSEa1G+ykw4y2a9OByeTKS5gXuvpCpvmbFCq2ltPz
dcjnl4TEZbIOKPztqqqHWxwwvObVrhB5U6CBduwm1QCNibzfsJfXdxBF6GqXh5WB
/Wlq4CCQvLHN1gd6BhE2INRbrHklSdyB7RpAFtogCPBY56yvb03o5W3y1/AP8P5F
06TWoiOFBgJSw4Sza+1sH/yinYGvfq+CtuQPi7TrVOy8tdnZ3k39wBlzl+6Ak/SM
S1M+T0BZIcf+rdoWX4LDjHe9X0CRTSvWxfDrZ5rO8QaxLORNCiHQH7l4iHtp1elu
QRr2/mbk4iZj0d6u9/VK8AFo4MdrWqHziuyoDipdQ3GGAR0Wmsw+B3P3BMoma8O2
qJULtnu1A78WE4e4Jm3o80+4xvbt47FruKlTZMqjfjPHYkEqZOc9wtHz50DDnFXK
5NdWMax3WLnKW1IXG7At7HwQldCMLLt9RdlMRfcoRJkXNAgXkxiImMMGeHrm/INe
Lk6lKS12PEVqfuHU8NjxBhAnSZUHo6HDxc6FFCbQmdRqGZVq/SO8osHeuX1k6cSM
qkmsOcoaRlEdC+T8g2LYvEJveUpnSgH8KnFZrw78shNAcvpkuyxZ0uDscRi0TFnw
e/4ms0mXP9B9Uz6zvL4YGCxivUmvcUsrfKKFX9Nh5zFilKDco6tTLW9nWVVZU6ja
xVJ8ZzNPqFlGO/1vZdhGPYmRUIfQQUi7xeg8yadBoAVu/v9sFKBm2SJy/u5h4mr9
PUoEPHt9X/74jdofdZsZrDqgmuXAv71Jic3PzYYmMgVSNyfXpbTHPp2PIY/fADhQ
hwHV91C5sGr5C0pWUGBZjUz+H89DPF4VoUgXlHMJK5mKfa/5N93aUavN+qI8jLhg
kjj7X10VMs8ATWxlSCx2ntJtGBE+dE+n9goMD5D6p3Iy4uOt2nvPtKUzm+piUa8o
41tgXCVC2f+rUMmGRAwZIZJL/WmMJBNiPUKdCIiPIzXB/mFyZkHl/TbnIV+UXBgC
edqlwagvISN9AmdsUQGcr54nHo/xISNDhIatojWOg8vhNQ7dfG4HzzZQYWxCSiYE
Is8c9lWaH5pgMUDXGeGNUXyW1CX0hO4xw5x5bgnlQKnGvcpDyoxGp32l1zbDTINM
RmnZAT2uCujhLYeLBpUOFYiIrQ0sqYPoiRvn2I3PFnUb/xHzfZYSYOqgn6sT3l3P
1S3h/yC2BLbgWfq+SQCfzUF64HnJFyN9KAAjDDWTiapXFtJOsI4ndA5sv5i0aSW7
frpkC68GnKTEuuXponM0Yy8or3c/WoevCa74FzSyBnMdeN2lyySn6KwbBjUlM9h9
4NfW1iOOF9hawqXRHei4zqwWYxXfRilpqMgny3zVs0dtfnVR4zkIuxTtwMBOx68G
M1wkpfClbfj1w+orJyan+qfh0N+vemmjF0BipptcwhxpdM3rr5w/SVvgwkaeqYlO
aEJYTrD3Hi5T9VySms956jC+lVLDc2DyfN3fER6rtsZ8qoahJQgQZaXvFGwTxdVK
KnJqkvyZ7at97iEK0UseYiIl1NDlIbH1v8ZX8xnOkqZoDuVJzO/zyTTcTSS2lE1d
x5R3l+fD8gyZxjrUz0I38PSC/TjmUv5FY+H1yzl4Y7WCRcJWuTaGOopdRRam9+XD
6WBFRUSdp8EA0AT3jvUNqN0xmeirNlurR1YBogyn+kwsoq3hWYHt1wTzVit8Purs
eNA03C86tA0OgraEzF7QlISbrdtmSfZ/PjEESAFUzIBRwIjIzzSiqQWb4dnSsyte
B1lTtQGQsuvQYBA5Q0jnTFHaXR/hE+5TmxGxkRnC0tto1ussfMQUTtlx8IpVWEsn
1MZsrBpz/xZ9DNn2yTFk/bvMcnnw7GhTrsUNh8gNKFFShTe31g4uPafcxijARhjA
Ln+ldcxd6wfFi71M5hPR7XYtYAuumhVCFDvEQO+Ky1O1xs2us5ei/c/YjfrNiTo+
bnhaaMKqm3ByCTf7jKuvph5sGe+ppIsgB9t7YC2h1WQL1QCau2k3TXNmLNvpQOlF
1hu2B49XjJBOs68s24QgwgyigBJkvB5etFRm4DvnSqQwfuMXRqswp3a2409y5pvX
ow5hRgcoTX20VjuGfE8G5KC+hB46/5qvh8spBNp0RqFEi1QA+itQiHQzVFbbJnnJ
K/kN6A5wXMm3HqFpQPaGHnSaO/wkI9rWSnfWZ18BrB2SX/IANVUxqOIxfqiuXKXo
g1uZWjcoMn7//vCGmscM4acr9iklCzcJ1458/AU6qZgZ5/FAhfdIDL4sjWGmNZU2
OzrsV1oiRINV3daSX6Gs13nA7Qb8RrhMg//BFc1Q9uVZRhjM9ZB/EFrxmIdA2397
2Jm5QpB50MXPskCJvj+ReYnQYVteBlt9phNdsCH1Uig6WXZbboJLGjhPqaRkNPJb
+tQ0B4yyxPIOzd7MGbaBQZ424jeNE5B83u57a6SJf7eaQzMUsG76KMtvDzH/DA3/
4aRmNQIn/fr6UdY0mD+tLMRRBqzcUcjhGGjNrte0Vy54fv3RHArqRPlsT5ln+3pF
h//Ny0VENOqXN8dbY3CVeGXkd6AgrJXEd/XGeU5mPxYImvKpLpQFWNy6ua3BpBDq
7X2bxVRq6lMjHH8xH5PEykvET1kzV1HqGYJwOjKOXFneUfBs46+rLXVdUXEsTu1l
tNnb5Xp7D3p1igPW3vZtGjHawW0LgmiyD+zuh+OuA68aLbc1aFkuVDqvsUWGVpjN
RGgwKajGRBGLpEdIuSSvUz0lGpTJ+rT3uP8DGzoihcka+CB3WTsyU/ftne55hX6d
RAp8y8oq/kmUc/H5UsrrZe9gutxGltTrgz0y9tk8xJI=
`pragma protect end_protected
