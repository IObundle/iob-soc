// QDRII_D.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module QDRII_D (
		input  wire        pll_ref_clk,                //      pll_ref_clk.clk
		input  wire        global_reset_n,             //     global_reset.reset_n
		input  wire        soft_reset_n,               //       soft_reset.reset_n
		output wire        afi_clk,                    //          afi_clk.clk
		output wire        afi_half_clk,               //     afi_half_clk.clk
		output wire        afi_reset_n,                //        afi_reset.reset_n
		output wire        afi_reset_export_n,         // afi_reset_export.reset_n
		output wire [17:0] mem_d,                      //           memory.mem_d
		output wire [0:0]  mem_wps_n,                  //                 .mem_wps_n
		output wire [1:0]  mem_bws_n,                  //                 .mem_bws_n
		output wire [19:0] mem_a,                      //                 .mem_a
		input  wire [17:0] mem_q,                      //                 .mem_q
		output wire [0:0]  mem_rps_n,                  //                 .mem_rps_n
		output wire [0:0]  mem_k,                      //                 .mem_k
		output wire [0:0]  mem_k_n,                    //                 .mem_k_n
		input  wire [0:0]  mem_cq,                     //                 .mem_cq
		input  wire [0:0]  mem_cq_n,                   //                 .mem_cq_n
		output wire [0:0]  mem_doff_n,                 //                 .mem_doff_n
		input  wire        avl_w_write_req,            //            avl_w.write
		output wire        avl_w_ready,                //                 .waitrequest_n
		input  wire [19:0] avl_w_addr,                 //                 .address
		input  wire        avl_w_size,                 //                 .burstcount
		input  wire [71:0] avl_w_wdata,                //                 .writedata
		input  wire        avl_r_read_req,             //            avl_r.read
		output wire        avl_r_ready,                //                 .waitrequest_n
		input  wire [19:0] avl_r_addr,                 //                 .address
		input  wire        avl_r_size,                 //                 .burstcount
		output wire        avl_r_rdata_valid,          //                 .readdatavalid
		output wire [71:0] avl_r_rdata,                //                 .readdata
		output wire        local_init_done,            //           status.local_init_done
		output wire        local_cal_success,          //                 .local_cal_success
		output wire        local_cal_fail,             //                 .local_cal_fail
		input  wire [15:0] seriesterminationcontrol,   //      oct_sharing.seriesterminationcontrol
		input  wire [15:0] parallelterminationcontrol, //                 .parallelterminationcontrol
		output wire        pll_mem_clk,                //      pll_sharing.pll_mem_clk
		output wire        pll_write_clk,              //                 .pll_write_clk
		output wire        pll_locked,                 //                 .pll_locked
		output wire        pll_write_clk_pre_phy_clk,  //                 .pll_write_clk_pre_phy_clk
		output wire        pll_addr_cmd_clk,           //                 .pll_addr_cmd_clk
		output wire        pll_avl_clk,                //                 .pll_avl_clk
		output wire        pll_config_clk,             //                 .pll_config_clk
		output wire        pll_p2c_read_clk,           //                 .pll_p2c_read_clk
		output wire        pll_c2p_write_clk           //                 .pll_c2p_write_clk
	);

	QDRII_D_0002 qdrii_d_inst (
		.pll_ref_clk                (pll_ref_clk),                //      pll_ref_clk.clk
		.global_reset_n             (global_reset_n),             //     global_reset.reset_n
		.soft_reset_n               (soft_reset_n),               //       soft_reset.reset_n
		.afi_clk                    (afi_clk),                    //          afi_clk.clk
		.afi_half_clk               (afi_half_clk),               //     afi_half_clk.clk
		.afi_reset_n                (afi_reset_n),                //        afi_reset.reset_n
		.afi_reset_export_n         (afi_reset_export_n),         // afi_reset_export.reset_n
		.mem_d                      (mem_d),                      //           memory.mem_d
		.mem_wps_n                  (mem_wps_n),                  //                 .mem_wps_n
		.mem_bws_n                  (mem_bws_n),                  //                 .mem_bws_n
		.mem_a                      (mem_a),                      //                 .mem_a
		.mem_q                      (mem_q),                      //                 .mem_q
		.mem_rps_n                  (mem_rps_n),                  //                 .mem_rps_n
		.mem_k                      (mem_k),                      //                 .mem_k
		.mem_k_n                    (mem_k_n),                    //                 .mem_k_n
		.mem_cq                     (mem_cq),                     //                 .mem_cq
		.mem_cq_n                   (mem_cq_n),                   //                 .mem_cq_n
		.mem_doff_n                 (mem_doff_n),                 //                 .mem_doff_n
		.avl_w_write_req            (avl_w_write_req),            //            avl_w.write
		.avl_w_ready                (avl_w_ready),                //                 .waitrequest_n
		.avl_w_addr                 (avl_w_addr),                 //                 .address
		.avl_w_size                 (avl_w_size),                 //                 .burstcount
		.avl_w_wdata                (avl_w_wdata),                //                 .writedata
		.avl_r_read_req             (avl_r_read_req),             //            avl_r.read
		.avl_r_ready                (avl_r_ready),                //                 .waitrequest_n
		.avl_r_addr                 (avl_r_addr),                 //                 .address
		.avl_r_size                 (avl_r_size),                 //                 .burstcount
		.avl_r_rdata_valid          (avl_r_rdata_valid),          //                 .readdatavalid
		.avl_r_rdata                (avl_r_rdata),                //                 .readdata
		.local_init_done            (local_init_done),            //           status.local_init_done
		.local_cal_success          (local_cal_success),          //                 .local_cal_success
		.local_cal_fail             (local_cal_fail),             //                 .local_cal_fail
		.seriesterminationcontrol   (seriesterminationcontrol),   //      oct_sharing.seriesterminationcontrol
		.parallelterminationcontrol (parallelterminationcontrol), //                 .parallelterminationcontrol
		.pll_mem_clk                (pll_mem_clk),                //      pll_sharing.pll_mem_clk
		.pll_write_clk              (pll_write_clk),              //                 .pll_write_clk
		.pll_locked                 (pll_locked),                 //                 .pll_locked
		.pll_write_clk_pre_phy_clk  (pll_write_clk_pre_phy_clk),  //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (pll_addr_cmd_clk),           //                 .pll_addr_cmd_clk
		.pll_avl_clk                (pll_avl_clk),                //                 .pll_avl_clk
		.pll_config_clk             (pll_config_clk),             //                 .pll_config_clk
		.pll_p2c_read_clk           (pll_p2c_read_clk),           //                 .pll_p2c_read_clk
		.pll_c2p_write_clk          (pll_c2p_write_clk)           //                 .pll_c2p_write_clk
	);

endmodule
