`define BAUD 3000000
`define FREQ 100000000
`define DDR_DATA_W 32
`define DDR_ADDR_W 24
`define SIMULATION 1
