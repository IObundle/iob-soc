// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:09 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V+YaqwWXXg+sIKJ24WCvK9wS44B7rqHzB0Apa93snS+zELXiWZZStLh1aTYiBBWP
ZR8dABN5WkJZLSKHSkD9D8TF/3jdgQ8ti0j9rWBJhkNmFGJpkQKnn272+gdNqYQ3
bh2otb3WhIT0U+UE6TemP2zur3F4a4mbdPyGvzcGjQU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18352)
qHOb09Prh/9Zmi+HqISrKnIHiTuh511xlutyIO5WZqj2axaapPgZwRBGnYZMToEN
lKLadbRlFXY4nNdQwsaZ7WQctyluLv/PPY495mZys6YCi8OfMVB7LmjVJ4R7qcE5
aIWKukiAECTQvWPXqHrNoXpjuc6Sxi01f6fjqW9ROm3tzc0EKhWllsTdVXuqeiZK
HItjJhrBLKl7rnOiPODBk1JUwaltbbohcDiBK/bCQbUk8cExacK80SpZVEtH0gDs
D16NXrBWoM/TwsvS0V8wG0IzyCRvaaChcptZx6dABK7ZFl8cj6IWNrHp4QKgQd0L
OKbJ1Bhdsdn/RjTcMMDlnZ4Sods1Rmqa2tJ0r9xh2zZ/4D8FVlPdANILt3BkM5aH
GymLOu+NQ47D4dU/dEGYVHGNkQePThAHHovwH43mo5r5ymblUWwa7tBqCJFPHk4m
mjYybBzw+KoctQhMoAfceXf+VJdkig3SswhDhVIVzUfV1N/tcmnfd9npbvNJFW6j
hy4wKd2Ic2gX76MYGfx8yYGS1oZqwBZi0vcAPSKX9jcBe/E3LVAoDhFIJbfsi3/W
fZE36SZboxuN0s7JQwMUjduEucmJ0rxMgiWIqvO+mBx6EmRp0O5LlxEdCadUxMVy
REcrpVhqfmuG7aXknjP6XTJFr31LWHlZimZG2fjZk+KcnbsWud11gjJUC4XbU//Y
YCE09zGYey/ZXGrWI62bTTEmaT5KNUivZQ44ZG1F9Q+lgc64waVj/P/63bv1kFeq
TkabDFpaB55vlmvF8NZ05blt7MFZA8votXC1ekyaowLvQ5vL5SQ05K5Oe/gZZ74y
qSyJTjbq+8LVMsFYJ6uZ/qZ25icPKENLcQSF8JrrY0Y+YB3H0koi11Ls21043IGq
wjxdb9TN6JW8fH0wPHwMzbmTYr04Ob+dKYSumygy0PimyyDy6GnNUcGKDoB2Cm8u
HrreKKwoptJfimBTEWgN5YNBY0Iuoc/aBLUgDLEpMw5f/44Lf1LVCoFsFGDpoJTw
o8QoJtWcbnQD84TBLWreu4d6h8ReAHkq56e6aBVGWAV8cXy06a2NLEhcBjapKwoY
1XoLLxqKIafl1eGtNl8d2jE+rf51+C+tD10XarFIp8nWo52RDWi/0pc0A3W5bsZC
suu8yX+QinaBwgzpWYsH/0XXrk1upIGz2CTCeU9lM6cDEVBCfhsmNRs5NsNkG7ZX
EjczccadOfJftk0Qv80jUzUJ/kV2hUJ+ShZOWj+QtMWCWR6O+XzkfHeOeDWwd0QK
3HRT+DZUjYDAeXO+SGY4DUxwCC1IuyMnoKfEBVvf8XDkEU/U6I26aRC1i5vRRVKd
pxLm8FbNt1RNV50nhuObz0d7Wj6vJj63md6qd5R7VDVWFbFn2qveNUJ66FTa3YrY
RuAmc9djoN9NN9gNDzNHnXkIa5qms89iS8l/lH0/OOXr6K2ZrVRMorc4xaHu3vV4
A38l2smdGZuS/srfedJuvoGFGUf8YStM+achbQFa+bYO8MhU0Fa3avMI3qbn6NEi
1FaUmxHzgdz/VN6Ehi/LrDBjDKkgBl33MQ7mhEIjQY6y75XEODN0Y+1Pm4WTT937
tQvaXRdDsCua6Z7QA2YhKQDuftwVB4SdNG3DM2/Smb1u2TExRJsTrM0eX2Ude6cP
9VErzFuor2PUiOQV3PIV9z7hksP+12xqK1CMMqYShLidmWA8NT01J/MK/B/rPUPg
v8BFwdEunXV5yuQV3h4q80n+EdoGBqRZ29WQ1ADwrRtV1KvYl7n1RQ2kG+Y9kVhq
CVGXhrbmdCWM0jDKiMvYmalSBv/lH6R21bb15k+0LdrqXjGsd7joZ98243O6BATt
eK/vxd8g1MHfgX+KxASaEDSgEyt7sNcWFMhrPrScuZksH0Nl5Sgj58dSrybpBttx
crHlbDtQW6/B5FlLJ72WzCpaNnnhoXd2C9sLl+gWPZI3x4wlv3w6XJrcKnE5NT5h
WWbrgWYZdwHyzS8bRm9qIFbrh7TH0M6ZZ3dJQjhgUzHyi7vU1SX4vwGnncO1lIcf
Z6RzTDT5zjvoJFj+W0WuRxXiCsfC7B0ynlNBw/L1EBc77nq7xXkVIXzUgZxfKFWz
HKcA1qPjK0SaiFqxr6ZQIXJRi+UKftx++cQKyBK9Inkw17LPqCv4ouYiFU6SIP6A
A8j3bY/2LbnlEVqCo+ChqmPOmd1Zjbxt1oKxpQS2LcoxLiY1Hz5CY2RJcaOL1FlP
I/E68HUBZDG7po+sDcWJpE600949gWMcbpom9jQwKLvMcF/EjnkckEMYtONtzZDl
sVvppU8WsepWeC10NYtQt0p0aer7hW/3+ryXDL9dp8q191x5XZ3j+bXlPGTFJGDR
MU6UsN5aphH78ZFvVlQ0e6uq+kZRVmPO9y85KGBdIa4v9LrHAMlvgAj5XBXq+jD6
TESNmUr+Klg+sXlrcmBwwOe+DS/fQSouoZ2E57RyUUjjxHkKTcJ2f3TWlXWPXAlP
89k+dMz0syBDOeu7bBDFV9CFkAUKfKz4KPT5FXmigNao5zdXfYK2qa1f1NRoWZgo
TVDKu2oQto31hqefYQ9PxN84sdM09QLzWRAiihJ+eRCL2UiLZwP10vIio717MYxU
pq1tbDxMByYrJz9F/p/uNvMd2kJMSpSGMfvzDIsMbN+P8fcHB8lT1xANxdbiDiKu
qyR6BqBu4zorM05CZQsrBUfb+TLwMv4zhv99kFncn1j6r2TrClIoyYlKDfD1At38
0/KnLdX6LAfpbfkwM7g3/vxJwJ5F0ofNLZCMNyeYgZRdk9KeNzLOw9xPeAWRHnQh
rrk4Fwo7aI8xx+X9ViUF6gTuXYfikLOXJKeYKBRNhOXMSWO/sW8F+sisDDQ2mbPS
/jndZdF+xWc/Ra3vFMgoNv/419Yh7OPOQk+tXgKnu7/u35k2sXlsPnBsNS/6JvTd
Aqb9RqbZzkDMkaYBeSCk5LzAv/2c0Ay9CFeVI5O1ZcRej1c6R5YEooMYN0B56pl/
zCr5HcuwGjBh6QP/GvtRL7LNxHg4WDDqu76HbBp0//Ut3K79BJXBH12O7hi4kLbX
qV+xFc3BiCxJQHdjkE2Pav7Y6fNNGnnEg3qVldnk9RvFsTWR5gMwQ66x9IJC0ghd
1t6vDZxoyHHSmGC3/aLUEFIU9/fmuPlNbdhtXLdgh0TBOYIq4DhbQJ0ztEDld3LD
lt74SoqjheLLdZd7y0Q+QjxMXtqfYJPpvGpDjC/ulNcf08h5HmLdJ8HxStzOJQNn
ERcE+aVf2D4X556+XddqyYfpaZvGMSUM+A2vFZfWm/sHCVJASxuenmCSSIEVeWNH
AR0QCwJp3kJmH1BK2aed/vV23HsOoVHTWB0ODBWu8mDUnC74Dun/B22LfLtLbb16
USL3UsUYtEV7uqUSVHIHug3TUIBYKnT3Gz5eiPVSriQe2vovQ6fPCfca/s7Yp8do
wsbSND24du6J0cd/uInJSMXT6dDNbokWsV02iaqx9SN0fVeCZjH6GpXsVmwrYm7A
a2wjjsVIUnYNKCaFji5ylqGHQFOkYfbBFU720RgpmMrocRjKEz6XVe+jMA1DX+rk
Y0BYOlGudYQiFTc4FNK4qdBA1SMD71OL9xBJm7oZLgq9Ns7SQd3NIGO/W1UhIbvV
qXxQwYPw1ZYa0W3Y8ycP3ufHdeQJXP/lvLfKW/h9alqz9nlwbFTciFQsPs96TODi
OOG3bHmB/KzEJE/7UgPNMS3b9V6mI5APMdIx0MwAFyw0BIio7wp7O0C6Z71/ycM5
tZefSfouqrZlmUjipE2cNdRHfYQzt7M1phESNsw2dA3WK/T8M4E15TAeozXWumqV
wB/YOsGfGlpl+SYDqg4A8ILBKy3YwZIHH0BiqJAF2qAlr1tGCUMqr66xf8p+FBIt
MmetEWacOVba5I0AmAJ0VJFGi4dVfFayNfMyJOnGPhCSsar5DjTsmrhF9Xr4qQmy
UgyskjILsqzx4RvgfIkKgto5bjkK2F9+/6qI/5AXLtKXcc+qlLy5X5uCkDtMHAPS
2IzyPkuZoPuxzFmc91hP6WizoynQRo0No/xe15MWwcYRos+SqsY7q47fBwFbqi1M
zvsrobmoaX949ntVaCIjrFwrxRa7CLEnQZohM1BuxP50C5adOtd2v3JWXFF5wSKV
9XuO5TZEv+7gGhWWxWMKaxY1jSS3Gp9DnCJBI2q0z/PRCiPR5A81M83B/PE4Mzpo
mWUzbE1KdudcvRjzIsahKK2je987v4nThJKQtrXv3HiXjidBRqEMtU387RQ23zot
g1A4zV/4Hm5IevKn0pBSpEwVb8/6X0W/XVYZLwYbxN42ifduNmZFZyfVwcqrYqXB
7AhkOQhWdPOIyqCgWoElN1yrR+3Py+EfcCDHmYifkuFLKhP5qKMGMv59m3f4SpKp
yuYmCyu/mIGESYkl/E2fFJIbZy1bRyrqkV9CsyN144ZpFuAP0PbVHG4V/MZsQmLR
X3YWjas74eCSVcEkVXgEfsTyKys+uXkJsRkqsPxkbULInqbR7zv5mTjlk81KdDEI
XMJKNG0lC59VokRZoD7sYMHhyO0g2nPmw4ICfULQ38MsoQ5SAPWijlo4opDFjk6W
cP5TTUOwKLNfArjaE9WEPh4YzcPTQEXY0goaj1WkKAZ2cM5gjvcXJVcBvg4YuAKt
Z50bE+0JKQrg+bUhso4GP62VwZmJDw3BgbhCe+CpsyI823ceBrTviQAH5NLKwKqt
9p0u4Xi478i86sTzHOqgVRAiOKpjmiju2V55305pAiC4DvlanMfotzo3RQ/lGrho
wiF2n5HLx60oQEp7UKRdRMV0z1gnFDELd7nwG8ZnMYOEwMKctCrFcsdiYVoTIdat
BYLB02ABe3NczZOMGpgz5crTKwYwA1YfMisP7CtJVK/fzHnTbEDcoUzq87KyBvW8
0x+g8I82uiIQSfd6xc9tgYn12G7TEwk3qfqTJZZYbc5DyxQP0tDwPHAAU9x7rV9P
+ZXusrj5GDF4mqCW7qLb8BaqhzsRRJ8i8VycEcaUjQq8+8ytPRcEQjmwjKOk4lhy
AxIHIo15pIYTB4dDpfOMSSS3s5BXNXW1J8YPnhKrqMzYx2eRMG9mL9DjjotTpj21
FQ0SskHA4qNE9ZbUe601DdKr52ZQKZbmgJIbVwKloPxYMoTL8P60xtFpWl59+VrL
KKKjxjuorRq/1yNDJquJ8f9exlRnKmTDuRjootPN4Nc0DHpW0QXZmIKxPbEweZov
31pfztUusRlP/lOgVcp+o2XLl0omTRddF5Ak6q3sZosqpxZ6TatoXdPVXC4w59kt
zXnQtJp0fAGG+4BYmknAvldzkzuobnJpffXGiRNsU4gmAJ/FixSnt7KxuCvv/7QN
WA5UpzFwa266+NgFr+Q0OthrSwBfovfqDx/hBvpVNgy8XImFNTSsBB/gq7yw69Ry
2CTP4kTsrlmB8DduvhGdI2Fde4oAYVIAUKb5wZglZOZPPXpSVtIm/jBzlZZ6t0NI
SsW4iNleQBPdVGFVi+OyhPL9WBYJWnJsSU7xxbxLqbkDczEVB5SCFcgHA/ahRPn7
V8YJiPOLLe3ZzJQgGt1g9YpAnZMYMFW6OMYBKePHNpSgtATRPTxzeBHBB8t7rmK8
CGhOKmEs2zMqyB9nruAKdUCuw/qvttOd10Xx8XQlzrLtsnFvbauXyprA3NEploOc
8LyCRlajrYJyjo+cczrlOoVIW1jMbiSrRuvBd1V3Qg5PKA9kjuf7fGVxyHoP1Tt8
bmg7EAAkC7YS98ltQ7hlwSMKMekYrCJLM11VwT3RHEXIIbiFUYMNPSXqDWiDQpmR
t6CPes/2NyGXNIXvu1fmvKGdihrq36Qo0Q7LIBQ2v6RwUXWaFOoJ81upPMSA+DBx
vZ0cORNWLg+UQuEpL4Zr28QM4nzfh0Xm906VqLIsm9hKSWMuE1e4yp6Amna+ODTW
1UGWr/m8g79oCSmjXSR5SAR3Ubhlrh3AI/kaBGNSw+FXaQnGhEtgrfeTZt4OOBZ0
PPs4yPrVQ9lmH9pDzX/O/FUWo5/tz9kvDYST5+2NeiOPqnJ0SLMo6RZPmcqmhyhk
1V98f7Rnr/P3VT3SYoyo5Ya4tJAhObai4aluj5riqUaqzSyUW3HkIhFiKhJdt28C
faG13ZmXJ+L8I4xvexobOsCC/NhIOngGUFtwGHw+2KmF/SV/kbsq6H8DlQ4Abvo1
hjUkHqDlB5AG0oIfSQPUt0lChxAH/FbLiv+mP+ICPJ9KxJWrGG8HySSHurpV/62p
3NdZ1lExxboapPF9KyVIEXGC0DgdAGHtH2xbkF5iHVfRoma18hpTkNak2AWvM0fh
HQ8q6u2ZubAzqdT1+RSIQb2cmavRQnH7+FyBMSjpY5tSNelse0Fp68PyLaqNLH4X
088iXs8E5RO4mRide14g82J2EaPedGX2oBA3te1o2gaEWTxoc6TkcRXgrfK0fqgy
99LlWIInaRmysJTbWMtcfH2i35zSCTExKdqmykCXEc2zNCqamcN3fasZ++aOao1O
Hm6YbhWTLA/mU+nD7CR5D+OeRXXNYru3dT5a0nqQQlp2yvWMU8z4JFDU7yXmXxP9
6ZG/IHOVozBLwinUdxuFP7uUPGFxeb6UzQ77a4X/dfkmdRnvr2LMmDWgH2umrdHG
roup23yIu7laDBYUnp69kFAbwm2gPS4AoMUCaTd9FQOxr+Snl5qcm0MXSQXKS++d
93TsI9NwoA0MmNNhJ2UVPBHpz87w/8QXED+6SFJRnEWLhfgCEL3n+PiK/jooVxtk
NUzXaZMOV1djJ5QWJKJ0cKLx+vbPVdKgEoIX+kMQ+FYrscA38UhwUGnEw9sGgh1G
ER2Z8QmvMevvd6aRNlA5VfASf2cD62otdad8MMlaTtfw9Y2lg4tvB6ZyhNbw4cON
ciEGE61n7www29oKp7GVSK3JmMQ10Ihr7z8FYEP6xzgw6QQDp3TqBRJas7Dy3Kmq
EvIePcGeOUpU7xm//2YAkvjqtAk5IsRC/xOTwIZL6cDGwERnH0RV6LRb0Fd1gCJm
oFTOJVNDH5vb0ILiyDPUgyP6jfOlaCBkU/sEmATBXzj//9s9EJ1nVxAZKLLye5kb
AqmYhTE40o0SbNfZYS9YSIWYvd4bo6qwp/DEGWPocGwnqIKuweCpvN+oqoYaxDvV
ft16PQMIYhOFVSSsIV86HRXTixsucmus7GFr13PfukQrHBaGnVjsZkHv6GEefmsi
3KFDWW7j/Lwco/aj3EqmJ/Zh2Xxi//wQ+Y0utenPOARzhmsgYoJT8xdQXR7Tkw0r
nb2/ZEH6F5d5uNPWlM7npvpGpwz68zRZmu1afEKWKTSeSqgUmjHmQ0Pn0mOBOJoo
vv1eqwRuTadgUodTa3QgjHELprn5ZBjsGcvk26AN8uBIzfbqjg97UmVKGzrBG+Te
L0g4IKXojsHj7vjjyFEOgBK4yIK/PP/W0xZM3hYIJAJVPwMm6XSpedsAa1x4Ukul
3pDkGzGrXKKzDP19Syi3Oj+HNpetzQCFPE+A6BRBtXVytMqCPyQrpC3YiOYzuS0U
vUOKA3i2RMRovrOW44MebVjG11rFPlKegq2zLY3HuWO1ytZyhaRRB0/1Jx09SP3r
3Tq49Atpt/XZOZgoIw8os5wKXzBC1EPV2wLV+0ONhMfNupbtZbKlgU3zlbZE+0ws
o3wKIM6DEtSabmvl78NHwGT/GEaTNH4/Gum7U9/VmWoVPIpviWqYSrM6Buz+0/wc
NMjWjDCaQHl4dP8pg8w/b2KVRciMsem2LiFra7kHz5EEU1e8bmP3kdSg63ZSM67J
fFHErqW7Abxw8qc236RjljeudgZdpTPBzuaZpxJE4GKXhLE9AvpHMuTSvxyiFAD+
S87Kof1xlEQ04cm7AoTCSDTieaX+Cok2yxXT8vud6nInjbbEXtzUwmpuB5SA3pi3
Z0qWXg30HF5MATMsopNMADlMU5abSt/Wke3gNY16wJ4+2TenH2GLWSlwL+vlOcB4
dw+i3meYx1Mdo75zBpbvPf9ZfW0f/h9jlqJLa7vreZNZrn0xkpJww6EE03r/xA+Q
+lFRLtCLJFtvNpB+ZsyT/J56w7Nz0sd9/ZFcs59XvboKYmKCn/XIC7Y0WpLkmnVC
xbdRsRPxKOUjWFnu3IzM1MLhz3c/Ki/XZ/d2SLPP1NYnETYppltsHKwKEJ7DX9cf
8qAMMZrcfnUSSDX/BHb3HCGav6PWYS5YdW9XH7gQ3C8mqeLAEcDVTZJ3o4hHlXdq
bem9j7+RAHGB/AuZZCPq5UxtgSU8quv6T1m9fu70+SU9EiOlsmitQA1RxBlestx9
RvGQKk00pUjeUSAtl1+UbNLohFm0OzBr30mzG/HEIZThWOMoL9voSD/HO3MCJavK
1XYp/6C1c4K/DhURjgIje4UhMCMO4CEDJ9dO79v3EbKW5BzGnc5wXMuLJE082Bqp
lE1faPrbRM3//r81mYF6x0nL4u8rAtbtEgAduJHDl64z0i/ySjnKlnlonv0AcIHP
LSLsQlcvzbtgKAPtyoIwLa9BSFgMtPqLc/kQshcw3Ju/dp598orY95X2+JRZin6N
Bqo+qqd1t0SOmYAuMmzEqNJ0cwQzsIn0UADg5WZ/dIWkWIWqVyvprHUAaLG6b3RI
LHujist8UIOh14V7ImQDOuxwPiw+TXYK996IN/EIVv/8lSQsqlIzu3mFMo5e+m/1
9ogOhGBpD0HLh49rcA5cxYIzrgpvvQOpt6bNchO6YM299FwPa4mAlSiA7ywlfoh2
kA6+iPD+nvBqfHvV4dJguJ7lS52HoM9dzzjSiWDEDzl948yj3rXWV0awtXxDsDdv
uWpgqKXWLCqAQZboW5DbZhHXvo4VdV7ErDRCHH2j0V1auv/R0PRcAEzI267OZiA8
BBQ4R3PFTSiLYc3wHgvSbmVlCFoRkiv2X4+x45y1HxmyoBol7hYLZhzoHIzB0H4i
isMWhnjHS1rrieL2plokmwZBNnyUi4L/EjQa29E80P02RMftwXGJjTELAys3UQQR
D4rTG8wyJqD1qbGKg/8Rsa/bRXmQWckBMW0znXZgzfAx9EgcN22EPTqhqDAhT7PQ
E9r7p9KA5HhTMsaWbDufA1W/S/H0+TuisYyGBe9nyWxkXVHtksI5COEPC/+B2Md8
78ERbI37OEQxYf+n7NsfCDbZtJvGWPwj3SJpZ16IROyMtLeIW1MKJBYMKi0a3uZ/
IK1GahvMYTjkGj+sgzsJxqQVZZS4GNsUNxgkFVMhZJlFMFW1Byl+1q4F6GTvV00Z
NepVz0TbXTL+6jtAXIck93poKNDdpi/bhXdW/3FW68/k2cGi1ym7muwSL4HjMWfe
Bit3N4VPLh3b7fFC2XaqEOy3dqT2/o9onZSudKJTGwCPAQnZQuHRcc2xln3SZkcO
Hzamzjxp7hGgazStC8Z9y1sv4A8n0/+gzSrbXp7iRyqoXSvXXelAD83Fs7bAxabZ
i/zjCQ1OPXUNT5+x7vgcvyc7uQyvCdAAWWJY44oWLu1KLkQ1taM+hczM1DRd5Fcm
dS3cUgmmNpZDmFgmP93rYdW9xK3s0iZLMgy2wjd6o4igBRBTAL3UwE/ElENVuc3i
qHxPgl9LeyHu21d5/1c4el2TcFfjiMQYZkWZQeWtZ4hAx3u4Aspl7izMLTmHGVtV
k3zBptmUbeqbizgOFOMMGXvqkEflJhlB+k2uc382PlqvfIERbEfVTBffJrmEfkdc
9KI8ed59UCn34iNK5NB8wAgcuoWAxZjhallBIEOV/SgUhU6clUrsh4MPqLohLxAJ
U5C5JQveg51q46QAgLUCBxu/hAoeiy0msTFOfw0jVTfLsKA/krNzU/ylGM53ljcN
dRdQuBIjPmKfGhri11EgHWPC4tZU8iM502Kx9n42PqyT5KelWkjHrnYggo9lvs35
yAb9IQvWWj1b8bf1elc9jsLdzvCxG1RXNYhSHIM0KjQ5PhOFAqMAU8Y/G3Wu317Y
Xz3zHOGrFtRT7VIebSrz7r5QS49dmwov1lbNTeUWnvwjFRw2H77qR2FsSBHqGSze
z0aIEwWggpR9n4pXr7cFk9xdKXSTOCqTP6PE453YQIVOU48iTLWuL0UJgmqN8CMw
9vBzcUueeKy/ukTGdkJUia8QI6YsJkPLxqwlNeL/difONJtPzAOU+00SRWexwEeB
eeW+JGQKCu+Oz1Fw+w3LgohPMUTF0Ukv5JM5TR74ymTrHOiLny7SjMfQRehV7mtU
YdLuGrzXyqu2PDvfj0S0z6ZC6m6Nztr3PRYEfIdn7LNmHtxHinsUi4miuspidq5p
y5Z1EeS9f99miqrnfPKcH7C40ESSGqn9c7KPIS9hDly/UVQJkDsg++7/KcA4DDHd
f/76LZEY8mRvkybLJJkUh62tXyFFuFdxrM/eEJT8hePTdvXhfR3HHp3b5iZADHeC
KWb6i/0oDwEyBjSfT+4VIu5H9c5oyDTlHsTMhRmNL1KUaAzE9PFDawRokptYhkIy
FUgC8C32aTaUtxwbJ88fBI6nvQWChlBPLOsADy0/wuqjld4vaL0Ce9xP8++7LPzQ
webAgpsnJ5LKQzCQDehKYm8CNtPwmn1tc6Hd+uOGm14BifBEEdJM4khDJzxSDqny
PXAii43C/yD8lLWJN6X4kFS7WuSjL8mF1MrL+R3Il3m1DYBu15DqqHlN/9LJEznY
aBkpRBWIqgGWOxOLqcEcPagUNiaNfRxaQFp++TbHteC1/XOJ3hWSr1MUGBbdqpJv
SlS9FLn17Pg0QD7Llx8lB45rGb+07fkC6sxVfPc/KtiTPgEE6RG9VAYDK6Hlg1s/
68KxNevoRJ4OBv7NyAo4gieUXqAzvxXmehihlVmxUAbYIDEv3gH3vzG6HV4kirYQ
+CYtAS4b20nDDO26UgNrX5JJLtELGS2M0zKDz4cLI+6ILOdFI1kHYoYPpOJrDOYe
fLe/RMlojvewzB25NlWCPvnBUlk1W59cnZs8oQWtfmUbFihm5JxyezAq3gziqwU4
yIeeDdLgPiYzGsXyJ1N5gCxCKrpvr+TZGG4w4a30i/GBCWp/BEi3zSpg6gZ3KT3E
V60O7zuUHJhxXJF72/yTjSKFGEMhc+td7XfSESoNhYdWD+DgoqJxZyBl4qC0fhnb
Fdi2ahwL1F6XoTUCDC33G1GcuWUvFlUUa0nP0pElxBCLlVjC+UpjhiC18uxzQqNm
2NDg5F5WL0S565KIdK2/0hcEA3WI4S2oAT3nssmMDyZRwsguxnEge3Gt4/b+B4cj
CrUsJ1GHNgkQzKIobBiJM9KoVVbqEKFg4BCr9OteAbEJvr0SWQgAHywt+XLL/aPH
IBJCngLJg+MFUBRFXCivtJ4lZ0mJxEphXQJOENhl2g/F2PDML5V9NwHowTqXLwKg
1VfPYEmco81bSyHRrcvZMJz0uBHyQh+/k35BvSv6hNpjSLgWWe7bhTA5ZImgB7n8
Ln/V9aID3uJxZW7PeDqR/AP3f4pVeEG2/t+GYwmmn1UIUP5Io49iGFASagSuniLB
iCCKgjU8RFXupN6hLOCAWJmXWFklm+ZuExFj+32L/8ws/yTKnaid8zCreZcJ6pL6
RwFl72v9ruuKDA6oup8JcuuO4Tvq0IxnFaB8CGGr9X1XFCSSUhfYD+kzmjrvsOMU
yq6okOZAnwbQXu+xd6FwrDQjqSql7PoiK9NBO6laBqFw2QwePV1X1f/jEGY7DJtu
wG25y+beTIQV7PFHLm5300u/CTYTjXVX4Ab5nI/LGfZ2URAgqaBGhKXEDxcY3djz
+hpUtyVQhPV+lAmJDeMOYt6e1IgIeybSU13cMkecSUkVPg0vYSAQrQhsUxBjQkY7
73JvcfgdO5AQaW4y8zm+/U6rzQbStyAJR1ajrx9koVYAsy6OjSB9KI6tWLC9Shq1
9/4X4A6bqA83f24ed2QwV+Xl3Wa79MmMpNA5PPGPA78hFX1uOPzCI9g34VYrFrXl
mXypqVbE73AL9DkDtScABnuurmchSmOxur45QSx3V6u7/EGPclu9WBEj09AyE0jm
xOnuyhK8pYB43uYsOufrpF8JX0nmslbrikzcmlpMtC6nU1KTQCAdwX5kdRXuFncy
JvwB+HB4vmPmnP2DG5ulTvRLO7HNodSpFVJRTDNo175xxbR6bzkwWkKTIboL4oVl
lvmbf4gdZtYhkKEISVdkZDVog+vZR+yY/HyCfZy92soeLjlnJm+5a1v83TuCqw1u
WZ9XjVjFMtFrQWDiWC9o4T1mZiK1ZLrKefhC0jPCxJEuAT3/C0c8Kf9fdFAm0t8W
I+Qij6Qw7l0PVA+iVgDy7AS8Lqw0ZBlPLvtcFdecwEl6sFnS9qK4R/t0eQTH9jhh
w4aoXW0v12DboVejpato9O2g+tanUhwgZb19jTipXpsi5UHJbAqNG9QKkup8xJyb
4NXfmJSpKxuYyqPVO8FjO9ke+/oZyckFkDjhUqQqOAVO4yA4iIuntHjalbx/lsAH
2gilQPtpbyx/XZn/eCMQ0fo7w9UMQV4scElw2YNkA4BQp948yjgmI9EuKTDWYQed
CjQ8pjMJzqaBobjbPrCT0vgZosrv7rgwdb8V8R7ssxyHQ3QkV1mLjXxQ4X4Tnml0
D0Ap18zmRIQ6FzifmPznUH7FIvLBLN5G7ID5CUuAjiXJzjruOTDELaRf4CbhJVm5
ztmqMPoc8tuxKVPZvW5GqAG3cSXuXbklq2XqDuZxRzsJzhXmgdqV1ebrmOewyKCg
E/VLXaf9IcDKkPR5rc0GPFvYOtbrXTaXephR8ePhKQjdh/mixUjjtW9sxgG/SuE1
SURQoMpJHiloGP/bE6Q9KxShgy3gA8PlCMaZOEQjh9HvuoiZA+fNaCFOSsHJvhWP
E2q+MrbVnAOjiL6DDPImW6aHt8J6rQPxQRI52TWeK3PnPkQ0KbIqqdKZAPLhgPT4
p2L0Jw4kA+lPPmWSp4piKi7HrkGttcr4n5DEcl7Myy5qVdePLYZMZXeEwP81XCH0
z21YHsZYAA6GSUwuGlxxLcvwKjRbrPZo/xIryq0vKJllzw78VaU2vnf8oh1Jd8J8
FCbhnVGUuyMeHRw6pM4WfknQmsTJD506V9fAs1QDwxw4xdTKJcaXy7O0RBq3CQwX
p2RX8TvpAHBBV76W/9LgwIAoiqwzVqbe0MDaAxIW7FpahAiw0WUx7lK+SWoms2Sj
S4g3xD17n5mzImnnAm5jzKzMc+kMISRkIi4dQaUbKTjsQybyVgl4ZQWALumOxoV5
vMk4KKCBpRLfgSXj6k0sxxbzXmHwXQ98UUfZ1heJqaoXN0B8DNB2uLhNxRe+DrK0
mURa9gToQfqU3/eZlsCku1I/I5V948Wim3LWKRi/oSm8f4qk0aLocdh94+jOzcVR
8I7ALWf7sdiAnvw7yyL3B3zAAWxUkQEo/olaRcF4rRInDjp/E1MpGwFxlL56xTWY
2vCqUJMGRMzts6DIObvRLWElfLlNoojp2na0d9AkkOkJe3F2wSEk/4sSSztANZ3q
wvVY4aR9kzWlQQRNLmQsTkZsI8230Xxo46fJ50JHkvEbRZTZcEm5WgCU54QL8NbS
2EFM5hZ1om1bwBvitSYmTZBHW7sZwtrVqh3bcU+aCszVn8wgQZP4rYp02b6SwH/4
8rYbjglbwGE8YGGS4E6Y8/iq0CrQjKhp5bcC18DRff1nbgZy5HblCeClhMz+XW6s
1G7+VT23n7aNxCNyGdwJ9qpJ/VuXliQJi6w7sQdWKOYR2S05x7djpZN+4WyklBJX
rFZ48miy8WV/BtlJAt5OcXxLJ/W+zDiNWGX8d83IIaQJL2UIXLaVtw18GRLLfBVU
JaQUY08zHmw2Ou4JhDc6Xi6sSKpM5woozGePFoUH+R8YdTIW4w//1ukRulMfo2Dr
OEZibd4C3HsyMfcXTcwPdy5HkTqA3xrsSSDSV0nQXG6y6zoi+/Zu/z5Fsp4wQYpW
IPILPCnLGNjGBBDV+UdttQ0pdwsvBXdf2BKNXLKy4v7g7w8y6or919IUWCxtlA60
3W3kkjoHxPDuB4u4jgJNWR3mAto6r8DWeR7Uos9W7o4h8o+zmCS5xbO+4gvpeazJ
4mZORrFoeSn02iRNRNNeV+YG0fZCTRwWy3W2M0+uEuhxxcq38vgx/xEyrcLWW44H
g9LAUmRQ5icJ6EMAWFLxRgPTqmtQ2B8RjVA8TBvtkajes7JLl8lvpGvOJO+ZcWbk
x/wZ2e4StI+6dM4ChlAgy/XnsECMtzAqdR1ffuyhnbmCyi5352JhKemV06l2hPTw
E4YaP5hAYJSLpfm7cD22BgqKjEUoRF3gaqymS79K+ZBryjCpJ/A64mNR/FT+/iF5
Lx2BwuRclU6YyMR1+QnPbg45LxeVG3lJMgJFLtvha1eMER9czlHaB0riybxB38Cl
pp5eCO8lcZRSp+nujQxFN25l/94MP4HetlISVT7Tb4fDt7VQWy3OOGkBSvSo0oug
i3jobQwM8PYJPBThPja64Mtmq0kl42jLUK+TUQUaR6tvxOxrT+KFifIPbwI1xD25
En4+1xGWFyqSOcBAk/Qcw313vud8Cqd5xINxdf6yyQGig1GJV9KFKd4Xqum5JIMu
zyaXOS0wf/cQ1JCLePfuOmTcM6ci5635bJSuwhKruM5PtbLopzXF2bdh06WUZJlV
cDepAq9L5/L8gGO0UIIsi/hSyLCVvbiY4XLw+0lZgpJ+ujiX4I22vQTs1E3LR+vZ
uQd+2hX24pzuj0asYmoFHQJ416RD4XwF0h8krNhi8trIjBR1QuIm9T/qr1vc2g/c
QUBdR+lRpcep0qwWthrDCtGCqoEDzqspuXmWNbvZts/H+ML2sJ3IBufkDZskx4zw
+jAnz5fsqudfCO8n+n4rWo3GoCkn+FGgyVBiiUT71tU44xzlZidC+e7Ulp135cVZ
zn75wWxjW+zbURIqPlubW+HjcsiMIas0GVctRzx4cI1l3THY0TR5Ez0g2N6Eadul
g67lclLuYu/98lPt36pj2ob6Ie3oicIPDVC/ofyRqzXuOA5MGYHXBIKv9XWVFM9x
gTSp4ZNABA/FKaMpHpvC6+LDndtEuJP8QwSlX7TyI6lFXk1ikuMbdBqw+uG96ekt
1q8j38+nrEpcqYbeoT+Imh2dL/6H9sbVrOBferkbi6tf3vMkBD/nAQOGSBhuLwV5
AgIiN7EIAz4+oIMLRGxiZuZb6IWXmo4tlAn72nIb23UesQBtpF51w7YLBnTr1s1V
Gb4ROSN01e8ib/PbZWXHLc0dmAqyRTMFJX7jwsu7uRAJdSlkxoK/xzcS4Ao85mPE
Sp3ouBpLoUqaU91mmip0XPNNRdo7OX7Zf7I9i4F90zSpf0N5hFMp+tIGae+PMqr1
UYFz2sGyO6xQ/jStK5vkZxJCzP35tY80XI9e31+YJ2WmRZkXQzsuhra9s5NEjYCQ
1lwj3M7+48uTHuIkVu4c2iBz9XxpJJlHEcDL76Axaj980e0GNkkgoXQaZKMTE0cy
DlSLR2z2PxRw7ZHcoxbZkIlRkiu7pRrSe8nb3bmLrK8QR5HMp/LLo1hUxw2JIQWf
5a5sImy/JF8uG2Vb3fhzbwRu8+qEjse8Mo4SJzy3ztaoPRExkmAYS2jl1QERsBSp
upFMHo//RoIfI3pvrsNQeOGwVRIXju+0NjdDioSoOa6j5+7mBPAMAgvO3BpuxvX+
AwCj96CRBBvk2R8/oIDzrPKM7MpCMmN9MCsLC6aE+pthHH3yoBLWqGXLKwBFAo1c
KE96zfZlj9FSghg/jOo+o+xHyubj4J+tOUl/rNxwJtpAWW0MCEw2XJ0q7tcialfe
xVognTVAV66dhMJDQDA3+6AaiZCXcv+g2ceyUP4QIbUPX9rJlx4nsTTXUtsshR0p
iIjMqxV24pSePV7GcWWsPNRBF4NgQ4MBlCN90Fp473bxi2/6I+5gowKJgRfEeW4U
Es2azeidii0qR8XBL8F6R5WTzMu65YO63k7uoJ34yU15SixVPqPlLF9To7PLajH7
mScrROsklz0uoVlZnAMLBn7OspA/djFllQCzQzm51LIGuFBmrfWap4YZFrl8AyB8
HMIKdYjlBEIzo2picaOtGZdaaYdQ7yx+F4do8NkoMa2zxQvyq0C16p8q1Su/5mBD
ycmaQFfz9/bNITpa7pcf276R6IwiAMMc9h4zXDI2PoSzQ24yVYiSPRWMG4YupI9E
cIbe9eHfWXtBbWi5ytHDNnnhZy75L+/rhscnt0rseVWjyKZ5bsfAXB8xJXmA7EHs
52mfrf4v1pE3Ve7OTYAVEFt8iD3/eSMzUg1BsmybGw2xR4gEPU+gXTLaNz54zAam
7VFjQ5v8fWfgJKDh9ryesgjbkYYnpwPr2r+RoLX9xYptH9fJaHnirPHc8cS8+s5l
HsK3ZEE0khc6wR7Y1rW+FlA6OIZrwm9vlIeG6dqyKYR5+ax/G7pBsgKvJg6RDB5P
2iBekqYlOYxvrbldX5K/sBkS5bkUWhJG4bsx5vcogq4yg0wTF/lfSyjnpdCWttku
2MvcBiITgxVCV4/7AQL4zJvHPkUua69rO3wsrNzC59hO653JxYIm8FFxna5clyeQ
Dg65MFxY+tWJBZ0xjIAvZkzyge8oXmOfAGRpJDpwpgQVdEHBxh9MxECrs2Woa65g
HAdRsxn7qESoBkft/SLdqKe4kOAV4RUjE3jPgZkvq70vvGL0SDIyzbm2lUh2KV7W
g3+7mtRNZR/DulOqntsT8VG7GvtlgORT1cErg0p+ruZtY9jzLBKDcdosWhXjFKYd
M7DJwhiS1H8C58Giss2FIZa1fdvQyOB9EwNSO6vS2HfEUKUwrl0EAhjItzy4I5Cg
DDXmn34wh6Iht9J+wbyCytIO0JlL6GufaT6mb/RbI9+6EN9L5oPEcjKJu3X0x6s9
4DFUkijFaok3Mj1jPXwJ/uV7ZBZCwzvJop/Q22eWegs7hYzqT6J60z8OrRNK5Oc6
u9B4BfTrTgsOoT3U1QnhA+jkVoG4ImFuckMP4X0E2v47HLqJa8FVDZaffj9YYFac
JECTczlzPbwlweokZK+/OFtxGy70Bx1T1K6Jsp+10Nxw4MDAsyUUIZ7SNW0xaI/c
vGvTzJfFVx+pMRCyhWMwTyL8eCPGyKs6y6ZptwGEfZB6+eIRGgc5svMUXICxqHNA
x2zwpFzC0RkDRv7UICvCldJygRk7CD/CYA6fnHOI6eAqSLRJ0GczqYy9PiZX6Wid
GC9v0lzodIcWevn3W9CT8BjyHFV5MhSk92UKa7wu2/IwDd/0gDVsL/MV2EFJvDjr
7CDEsyjs8wj+4UAAtB60syqZHomVcdBRFkmvre1IqycvGevTHaRKg4KSGlMqcTzj
6klBbkjUB5Y3LEOVais8Rif1eEiAurTIUKkW0nt+zsSlgzzIcw1crE0hSSrKdZoo
2PbMfZ4umO08+byEziqq4uqJIyX4APv5TxoIEEMEPwYYMgLWbe9t0KhuLR4/jrOH
9R7wV/CNpxdZ7q2N7+JwEAved8xST7ZIzLe44Asx1gBeXH4YTnLone3Kve2vgCx+
PfuRrWICyAsHWLnWai5NyZW9pKrtFsAx38yy+UW4U5D/KCRMuihUU5y9ih0aGkfn
6OUP97Lapc4r5Zryn05cvEV/ZLMmojl39v2BiCBvGjcDkDurrdcVnAT9RbW/XnjL
4dwVaZ6dfygtv8kk4ueUSLfWLd7fa2HWjFinA61XKGVRjauSy85BBupZ3z5pArG7
OZtL8YQtLV6MUqLXiNjko+WEnP1WMJLNydImq+XjB3O7hngIqogQG3p5viJjOOw8
boIDucWrcsyqkYhTfu5IOjU/MRPF6OMVTLHkVbmN0khhfNxxD87p6gQCS/aebYM9
tdeB0E9O29YkdtB/eLt3gCDwIbuy0QfD8nmUxUaMHmdmJ294n3EPY6q6tqzELy66
UMxWuIRDsMwqvdXfsRDqw4/YzXbxrhU/wnlEp8tXu/PLFQvvIPzxARPqYjbCWH01
oG3YxfVXfUdPsQVJc/fvKYfHZ4MJ8SdltMUnadwEWMFFHdgqehA0j/SHqPJ0Whpg
XVSbjLRLLDaJUOgbz+f7pNWwX1FVIXuLx0EQvBS5z5aADdDFkvgDgFr7ynn0xpLC
/Pzu1A8ncxFyGg8LPOFzjWvTP+W6wtTFU1QDh0IpbL9ehWtqvwnCavU+A9r6h094
/qS9P3h/NQPjnAi06LO/8+Vg7UXmd0FVkozy3iMvIUqUkqLCXrhuUoPTRuOt6e60
+/b10W8O6VfhIJxFFEROeE1kMxAkKwp3d1p01B7ZJ6Otyl0VGR9BIqT4wIFjXFUC
VQETx1Og+qQvYELSMhL1CfitFZL+H9kV3Ar/MVMImVjNsQHV6f70+3lZaPcvCVYN
ToiYcwDmC46A+vOmvJi/kXfsVTGo2/BAUAIR/+j3Si2tlvFe06NgCVKFr1uvamev
ivo6651EVKPX+YkSaOIwLRlGjoE48Q/kEtqJyNbUPa4bfqqeYONsqLKH/FyQQUrC
UQ+dUqHcAI9s/9JNjPrLTUuwB4CRo5mvhu7DuAQ/vLl2DKLla53UjGndcyGWjhbd
YiWNAAM1mI/7c7kThYOqVcsl3aSdGnLqHD6ncIXb0aMWWdiIg3fKIv4Vi6X6lRZo
8oreWUiRUhy9CmvfHTatdYT9GRE2jrCNj6TImLUSqcRa4atskf/tIYoUfTbrL9g4
ytB5Y0XEL8sEQaXx84WKk3w6DND66lb/RpNwEsxXLqKfyiaHIIPwvckNWjPp89ap
MpJrIKfUYwIqj+b1uSmuVr9Q58qGt40sEZ0b862+edSjPwbhk94oFg8vVrfphygz
3ftzXlatphhKOCjRHfsDOClYCWHgWG/SJTwd3ohyRRPhcN0hbrt6xSPmYsY1nOQH
E2lJjntIc4gEpaocb/uEZwVcvBORnPQkiPsy7uN6cskuH6RFRVy1Fj0tECLp2bhS
DL32Ea4fWRiQVGvr9GAThmDe2fWSKZ2uf4Ie8U0eRZHWB6I4XQ1/qlui6ElqBLWa
k2jpq7Quarg8WyAkX2yCtPeZ0wxCINkFvVLltRoqeCtIZ2IF0wRaC1YGLtEny02u
baSa7RyFTUpZQ5ce3WC9BA6MwbDivegNXv7u1ybwBYqmJFglzWcX4qg51DETgU7h
ZvIWzcSjhVXsqHrHZoQ0IkoI5JWceXkHfhUsPf984BouHjQ2BJFcq7cbjcZCqaBS
E3MxnbUQgf8cmO8cdLqxJ4LmpyoPCEZ/5kqJs1qlcC9UWbeuWrpjnqPOYiQAJzD0
gBaU+fqa+ff2K7+ivH4QqI98lwmFlWydXAKP/P9KtSxwcs8Rr78r6B5ovAd9yite
t3cWT3viSMB5fta38XH4AMdaImTeNXldYIyslfdLRmcaINI6qhn74zmuxr4XhM2M
0T+u2I6Tu4dGsom4wDGJUY29FXKk0OTqDZOXxw/PMrO7PsVBlLmKvLt/kXcaQRmv
kdhKF2nutnM4i8N47c2966/cckBhy/rgwUcMmJbzi1L7xCE4S/1w7NI+7WwtpJ64
Y56FbWDe99RBdI4lH8DL90Rb16j5YyEeEYRQIk6LE0/+iIgfsq646az/Um03x53I
YKTDQrayJ4/EWbjnApqtwOghmWIgg3QfG9Vpd6OLKJQ3ZQtYf1pSLQEsDV59VY+b
ZcVrn/DVhIr6N3m/LS+oonKa6CA2PH9wvxGJCocLkZNQstbb1sLj2Ciz5c7usdfR
jVZRsM8kQlqGZh+Zi06EWAA/JEcLLlwaRHLOzP/DTvtmZ4VunrZ83VSv3KwSf+BU
j4/ZYL3Buk5o9RPNxLKLZ8vigp6FCjiiBDpwbmKkmhri633sbIDLB8k4yn2pg8cM
3hQD23GaNKZ5lsxqC4hGyJNe2S30CE9wOQ1T6g1P1EBC9cvWyQlHIgOm5p9IYmn0
zIHZPI83lfzp9+pe2ttcRVdosdAx+iT7A+BKi2/bbCYAL0bF1B+hyHW54cRU/bSd
4M78/05pnNDB2roTxMI9N14xLiflM7Gvp/v6tc92Mxdhd/kthXMZSLjqac4kD35B
hHAYwdoB7UCnWAba9q1aN8UYtj0YTi0m1LlBWavahohVNdtR9qR3cslfIPeADlWD
FXpDNZgr8GUYllJVFa+kpPfhTCrk1oqN9eS5ik+MiQlOl6ySYNnrpFS6CEmaUqn7
hOulUOwn1S2OER9X7kzmm7VtNSyMRVCji3k6rujkRjlJ31WAPfFmRLcou4SmBy1Y
/OUpkDK0UVtY0H6L/+rxAff4rASZGBS7vWqVRpG1+UIvtHdy8VQUxB+HWWhuvd2L
7gL2SFeHoPxi1x21N+NKsZScuLINdXN0mZSY7XmY3eP3LlSbyDtzX2yxbx3BjRrA
FUMD1pynSLttmX5BrTGGrCGYS00QSVBCdm3VWayEnE7mlG5ludrFJX6xmXFXiTkk
3bVdVYzZdzOK+pqVhavO5V26nnL1obYsPbZnFA30RwXguOcUeedtj+UZTTBzoV8/
bxqSyzpldjIotPzn0PMHypI3SGdg38cfZQriW7DkyYkbcjRuJtz5+8FS/BiPwaEE
WbidNOMaBWDzU/H1HDCfJ2muqH8ZxpPs6SNHIAXgln22TlXurvPBuiZnjTO7k511
/sWtFKLuvBmpl9Iomm9SWJn/fHg3a+mfk+g4A0BfVVRggTSrq9d4s5GjT4KgSToe
LN0fS7giUwjsK3w7fsmuI6iCXwU+uNH1VaqmcBi78GfGDvL+1aQp8QbTzmkeRLhw
gMQE7XdWJuoHufuOVKWpf31XyNNafyTCm08Hzwo1Ybd3Y4OyWew7slhg9AdNn8Oq
oe23v6VXvAIq3Jn1q2rsOD/L6YgLA0v0fxQfxRGChLuxRGi70F9RZKq4J0+3p4PU
d1Zj6NtGwas6hn6JPst0LX2HJE4nGH7himdTCLeUC8xt7PeeYpFEtyQ5qF5L9EdU
q26h0wvaZbal60b/N8Pt4Gg/z2iFXHKHyRqo++mntdxpIPv4pMhjXBH1BwLFr2Xc
csXYX4BwBTmO2jARmhWWa4iVnOeMelDgimh8xOu/Yc5mlFbEPGzrX8jV9Vd2J6JK
G0FDuRm0gHU1bH399YfHIbOI9rKN5WSmhriAtLWoTVhDlnfC7XrbFK59oTvBcvIY
jcHnZCWUeEKS7P0I3YXsPcDtB/9K0U4ar4BM0Ckj34PneNw/EU/J3g0B5QUhtdKq
bPDIUni8IUcUGr3waVNthuBGuFZXWVlpU1FOJMvS+QW2DJBAurD0josTJxCbzDb8
wtnlklN6+uoJU57otwOkmTWDayRfSuuAHhLvVB6LWP4FiDr49rx5OfLO/Fdh5tk/
Kq9rcLwFgcsnEJ59DMW+mT7UeQLVqaNgRYt9lY/i/8kzmnLfl8Ml008RQgaUsB1r
7l27moUiBpS14AhLGkKdqUuowdjBd+neAmSma+nrLr3Hc3el9OB2F046xxs8hC7E
fPf7necclUKy7uz+2WAcg5f6crkgIUVcoY85T36s3GAfEMFj2DHH4yBcm94DeqCB
BCAsPSQ6C1Ni+4IfKW7DwrydORWzA1xSjd1DA0Kgp+D6OeZ+GKWFr+dA/6Xbdyn6
w/GC58JRyk2HjWJkvu6rkP1JU/YaIyxgh5PFH8bFdCYqPe2AEau4idnRV1i7OnT0
NPjG/pLTa4NL4l254ntqAV2blsu/fkkbcoAIn4wgoswiZF0B1dKqAwPNrPEQJJyz
2teR6gpmP71HqzzFESv0zr3BwSZQCrPzD4fb99or4ELFzv6IzjwzP15vMn3Dpen0
di3revNviSgqF4TIyzrJmmGuz+pdAg11jCljBA95OuxTBRQeT+4RUyAg58d1SKdS
fJDcxWJGC8VcYaTpzDxnCMtcvKXFAObsIldpvgwgcxY3yYFYSr7JZOSg5KZ9GP6y
UWcIGTalockPeNTK9fGXMsW2sCCSVKgggWEJKg1gga35h4tw72AIYR3JuFlMHDzT
2cpQvYHEDt+PMApSS0G+WMRz8fUKjCaSLSRUzV1aydubizmWUHYe5pXUYp2wDGWZ
beCCqGIjJEhIDJhD20Dk+f9YGK/cdymIZHcZQhgtwK7c8ve6uPtXEJXGphGjqGwM
FDNtGSMRDiN2Sx3ydOfGUIJCG8rG1ftGcHWOQ2ThnOLYg7zOPBHjJ7N/hL0bIwjd
6PWhYg+nDLuBghQBc5jQmdpRDwoNJpoVh3hmM8+zKi+gsSYOw/ECzPH14T/wU4B9
rFHF8/hV04VLc3cpuV9wrBd/JKsMbGnKDvbJQgAYK8nXREjdSINiZ9wBiLZxKlfU
2+lGJQekmVa/be/OCrMz0V96qJvxRUZGyc3XKzP9l+yCtDIdCQsBWEvTRQ0MlH+G
keklHxrTg+Alhhfu26vA3nNR63iKtkYjQlwZZcSJhEyxEWsq2MGQ6v95DNH/q7zu
c0d1eYJ2leGNx6Y6cy0vspK3fXkGD/Z/nALYK3b5tiQJS4JzKVxVFYbT5FoUhYpx
Lyr8F/2nllNKNS/LBqiuYKCu+Sc/URx76jZEBKd1uUFjw5k7trooEAZf6vGlp468
wRMHXj5Lf3qfTGoQeMxm/U1V7MvHOSrlRQdXpo8pOn1f6ecOVw5OA3zLJv6Ebyof
/cT2cBj3UxOqGavjeBQ/R2Sadn0C/MhmDgzHDgamhanB7bvA8kor5+qZmSaClbfc
aqphoWrcjJBxchExnbzQzZp3PBlkvwf/ydbXu18EhadOkKcysiH53AmbHEfEa52P
AuiZIBoTKQXVCTMemAmgowJI1UyZ2k+SqCKPbaoAOxAb7SbOOkmVJfrGhzzUqRGA
tD78lZJntBrKHKiVjjWjfu1wFMzelBwTEKOGWAyJCiObadCTT/nLtzpZf1lbBg8p
PHgktS7kiakHCeTnPC4MiAdEhz70I9K6W21vcXKH+H5OTNMc3wlhMsa2jT4k908h
cY9LkdhDmE1GcjaaJYboa4mQNMgnq3wYd8zrZuZxCKRMDNm7B+/f2vqClXpPUcvJ
Dgi6t5bNVuDGYIWzx2VSGRMrfTKMsOkMJNm96ITVmWtyJWsqiCbxS17/Gbx+ehoz
Bvm6Lw0byrUsumMqlNFsfmBCeFmfDc2+AVEOOxiYRNwWi4I3dlBw+D1m6diezNBK
E6m2shzkkwGAwXuWSAr58iKJ7SdyFYd8j0c8TGn6BmB8MLiK+drVaG8Oox/F9rzN
R5Rdx4LxQx4Hfpu/c9Vc69VeVTlYWwQDS+45KGQI0Y7fKY6kQpokRcUOGi4pfeMi
SZYcU09+xWFFyU2AAC3xt4j35zi5/scrCLcitGv9pgu5Y2j2U9saTJZAnFtQk9pZ
SrcmhNAS5aufN/33hWnfohxOvSfu2L7LZLhz8HW3dA0d6VWQ/4xKQohF9rsu3sPV
WdGnXd5Gocya426UECz0kViUzcZijQNbne1ON8t8XQX4uGvDBhUYOzclLZd9DNgO
b2u2mJ2giEQUcgSSkd66tlIzBvCzxXh2lDVUjN7g5JdEpLhbjiUElmWPaEKOy53j
LKvQEOUi3Rk3kiLRdgo/3R8UbqE73aWmRXcr4c6Jkz5BqzCry0QpJ6GeHEsVLbcH
v85vvZjVBtiXVF95lH6TznDorRH5692uo0A3oqdEwPl8YdarrvGv0ipR9kRvGIZ/
qG+X0StSkTIyC4BbJuKbjQNYYfcJE0BwLvZA71SR+dyqcTscoyyQQjxF0626l1Hv
kfyCANJYsk9k/S1cQSlJTqLNKVZud3/akycglmJmAUewDDVbTRJjae4L2cCYMaJl
sU4fkRm/zv93q0341bLmtRP8FA15xyiD4tedxbzpp2kQVH4W5coLTJAqbDPgo/fX
3L3890GocfZMoj37WM6d2tjoE25KZWg42Ozg6vKcBCYvBDj2JL9wxHtoHufnXAnV
3glarJsmvMtymHP8TvjCynbmJ5EG35qqG7rVJEBT/YAmKKSidjQ6K3ydXIYJx3NK
MvPIAU0VCZaEFHIhfU5B9c4EB9+98dNSaBTtdpxl8XnOkV5dkOkrdPJ7nPIHUAyw
+jUL0wzva+pm2pVI2X4l4/iygSZfgpBaZ8HX3f/QyeVep/kSZLKtXYW2VxCMjNPk
uR2G1/vOBBBrJBUNMe4pVoCTbnQeLgK3mIxCcri7kS0ih/XmstZjjgSmQwFGdGE5
1PiOO247NazusKFp1mG/iIUz6PAbOp9UkQ953gf/Y7nbgp/1d9lzF3n26e+WAMEM
LpwMvKCrPF7uXaH1A4izltxHS1NxHTS5Q5O5Bv3A1dDy1Wa+4SoYG03HuWDntPGZ
bf5XSEtIWVRWwCcTGKLJBqSH6Z1f2EvQl0vSRUA9ZYNCHrFhh84T+nmgciojYTLQ
Wk9zme5IQxffV+NVwtGwanRlMAOVJL/hAOumnPBuN7gbHhOeDkEH7FiKeywr5Bu1
VZdlBoQxmHH5Q6XN0Dw0i+yiElT2Uv2Mi7nyge5XkmPM2SWwZZr0Pp5olRqpoCKT
COsbBVVopkRD6Z6bFFtnow==
`pragma protect end_protected
