`define BAUD 115200
`define FREQ 50000000
`define INTEL 1
