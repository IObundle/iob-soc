`ifndef VH_IOB_SOC_CONF_BASE_VH
`define VH_IOB_SOC_CONF_BASE_VH

`define DATA_W (32)
`define ADDR_W (32)
`define FIRM_ADDR_W (15)
`define SRAM_ADDR_W (15)
`define BOOTROM_ADDR_W (12)
`define USE_MUL_DIV (1)
`define USE_COMPRESSED (1)
`define E (31)
`define P (30)
`define B (29)
`define INIT_MEM (1)
`define RUN_EXTMEM (0)
`define DCACHE_ADDR_W (24)
`define DDR_DATA_W (32)
`define DDR_ADDR_W (30)
`define N_SLAVES (0)
`define N_SLAVES_W (0)

`endif // VH_IOB_SOC_CONF_BASE_VH
