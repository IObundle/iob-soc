// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z4VNR5D9wxlBtQr6/JPtYDg9T+6j1DoVEOccwo7URnysbFuvaG2zRzWNqLERlnlM
PQk1jTXt+UWqOlqkyPmiitOT1SfjJq4eUkR9l47FB/EoB2qnjoTcExtGV5ls02w1
nhYxVrqFENL5tWLcY5vOKtENq5eAu6XlUXvB5mBEeqc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
znVst79d9fcOjc17Z35j1i7O5sAMxx6dTrIXeGMC8lquJKlmXpeLTm/vqVbDaToc
26GV5fslzxcwBz47UAA4wsgbdSUtQHDCx3Fz0Mbr/LXg2e3Ch0Ad6UkkYN1LvuTr
JXHNGMdJhSddyn8jd1lkct37YOlnRhyVwKVsx5h08F3BUrsGygSEqFTkAlqnLTKc
8W+BIuE4IDg6EwIePOYg2u+aHHNLMY8/YTlrDHRvxAOhjSxStrLmBG7FWPCmPVuD
afB79wwVEfSrA9vqhdZUcGQfbRxeVdy36ZQ9lKnKXkyqULurbDQOjzc+rXkKvVH1
rDcc42mX3h9DUDcA/PEbvObYD/ivlcSj0ZnL7qlVlwJ1IBnTj5UIIJEmbd6g3GIg
mIEbKYyWlHaxoIOjg3ek5MoOuBCv/4veVAKwaKhGzcCFqnH9RhkG5ZZFFal66h0a
08WKStngmc3HRFCqMP0z78WaU+dtERTm5ycqKIyCaSLi3fv4M8OA8u37veXiV9bP
Frke6RwI35a8h2IwP0Vc3MRLz32Nf3wiHlyILtKi1b3idcH0Ozh3jYSDlIwvHA0G
eo4Ww2G1/g0yXGj+DCrM2R0/2YYb0BKNwtXybz7C/ZayBi06jR1AM6EM7HU2mbNm
hqOXKDlSX+5noV8bcd7mRFWTjM8E+mge0pzBBM8Rs3ZI0waBsjZaxKXyHeYWbuId
D12U5mAmb4pkRglZUpQldT+BSc4B+k7ggNrs8dJwS+rGwFbPjdZpvgCQWZYh/ibs
dZkD4Q2dNnXkiH2tdo5+HJrxKdSV2griGB+28EYTC4Xsp28fpGIAjiXI4ogCIHTV
2dmBxNzImCy8FXd0/l5QNaICIR9VO2fI4MCvp0zqiUh8IfH6MFrR/4VAYfYJmDLL
0a9LzRWXd3zsT9GODEoTB0ILh9u87ngMICEv14LQuRliNtaYt61FhRhzb/Vc5TAT
veR0lgHngDXGI51CFCcVJ+2R/TEj9v6CO1oqtnANyKDk73xzSWaQ05zEUP7rm4Cz
WAYvHDVpWOvDMIqqpyF4PPgT3atkqZAsELHs5yR/Gpcmwr5+FK7DBfqmCMmb2ugK
lJNC6WJeBlHigJKLlslf2VrrYxM+U0FhMB2UB85A9E5ZnZMqExSyUb4T2wmBJTKS
HZ29UfBGanhIqRUe4gYVOfDDYqof4HiwQPo6XsNha0QOieRUF3qnqCJC2tqazv4b
dYeRVPpCoTbAQf8z4nfGF82GsHCOmzUJ1FV3ISm4yLXH+ivWMJexFqN3diXnDp2g
5pEobKCZhb+3E1gLk70m5dy7WemUQ43eqIZIYiIeSaD2AUUTtQyufnL/En39OPWb
pG9xtGt+snokvfvNxmjjqAqAhdczgJjs9+jSGEySwhHruiJYoyBI+n4Ij0tIRYw4
msGMdegrhTOtBkN9c7jh60Y+mFVlYJe3fP/is2Xt8k/5b80Xdi9PvGz5+/Hzi8ks
jTHoPAyATw22Q6FGRRNuWeoT9q9Hqf9nesRnoYmgxT5dDwGJm5VzcJ7/rDBODEm3
CjVmgG3FMYfPR+jWXrTTWm0zekBLbs08Cf9uD8+fikS60UWt6/8TE6lz4TkLCqTk
+AKdFMcHSBxD2UxhVbPwH6vWWUsDdoqgmmWxMA9ZR8lgzQDdZRKdbxzPlp0Ze+BA
IQtHpYI4/N6sZslGW+yArwpXWuPHlTp8SF4cpHKLmXYCQjYa0qx6LzFDJdanEguF
AHGU8jeXDYzollPJZfhn6ZXjFVUcXfGQeSboEIo3vz+HkMMtC+6GI0c8nIDKyJZE
6uOxIBgY9DSvs3Dlgru7CCkPmIPtWki8uKpLAl52wjGOIJKWNPgTiiYcvTKesa1Z
osjB6+D6fwuZ5o3PnZR9S7CEoB2mFr026IcIlYk8JUZWjPxol4LuoS3DHb/xFyZp
3NFjWDT+PyiXqP2XRqb3DhFdArVe2aF+JZ+aVHjTfKFcamNMkJSOiISGnMYkpHkD
5+uRhBfI6JqnopIWpa4RuH5IDUpym/aft9yCR9sIxTT67KuAKuxV4Cq+bscKEx87
MJbhtJ5bkypsBBgPyF6Rjdsd1i5O8LF+Jhv/KfHmklOkWsUNVLAdFc3ok66a9jZJ
RfqkNextZGjrmGLtzr3BLKOQw9OT5qyMsjV77GBU8cPzCFE10RAQYAtw45NSn6a3
QEt7KPINFbniiybdg3clWAm4ufr6GwUl1aKd1YmOpSkoEnt5aOItOod0Bxp2Aosg
lz4sw2K7gr6bqrDLgNcecdkG2ktgPyIUam9Jfi5k6iLNO5PZzELxLBuzrn+MD10A
nEmZJrN3nnNKmlyUa1BEwV9ltIkqngj4EQH5jitfFftBeF0IIE2f7tr2OuRyaOiD
2PtYRO4ZAw5JsLli14nwoD1sc1FYpcnTDJr0JKLJjrQ6qo2yBvPNvTayTcOur6nQ
vqiC/x+HqrYGjlOe1RCU24DlUJa6L6+ebfSiS3FxvSm4n8C4GmP8N2rlDkO7VJa3
an3bxFmq11FLC+vG31ZXfrHQuomPS8Ip1y7FxPFTMlxrQu+RALXVAz4ro72M9Yai
1hfEMsCB2fU4GxXJWbzm77mk4M0MDnhMjW1EwxxctC+3sItEvyEE6OsHzhDAQvNQ
grR3KldRr8wuzAIKeII+Rlt6qVOR78+W+tMgr7Sk816s3L8kF7VN0MVADit37TgM
MqTeD3SSL6c6iH0sT5BRrcw3WYiJi6cx7FKsRcSrR3fvG5Oli1kYk6lyVTHvYfCP
3Ay6Km4YBzGlYh2urnGayylPURnpyt9sGpGzYCeNpscCJnjVDQ9cIIB+5RdSD07X
in0OokPahxDPOS+EMU3Floz0ebsHOKWpFpOLcsaUE9pP/jNjihcswLhhjmC2I5TT
+3NJtuLProEoFzi/Y2g5TRwQMnMBz59pJ/XwfXrNhZfkPFtzY1DYv8nBMBMp2rPV
dgGuBEW/G78ZbxhvzNZ9HdkQeNUMLPGVO9a4i3TVd8US2L5PNR1dsyAdcTfl4ktn
zg95V++13FItTu5jcoiCKzH1vO6Wovts/L63aGsvHywUOcPpol6ksHNCfYcbwOxj
bVZTpratcrGd5gTSejE3ZI4doECMpy9B3UJUEowHKKH6WgxXMXsdhBezjKLhQQ35
HI81zsHla/+Bj+V7tX6RJ9BFzCPiOBVKy9+G3uUFAapll9JLfNhZy8S5n4EBu04q
iLIWDk9tJ08F3+OVt+Qzu9lzqS8cSq5Mt/Sovh87IH1PUnhRniKl/V764l7i4nY1
0UoGpwZBfIyU/3gFWkv42PRIQpGDKisRsE4/eWaY6HgwkLCOfhWdQs1bi6wP3XBZ
aM3ml72PgVgqWfahwQOCZh/Qxwuigas20z5pUwymayYh8PmQzHlm+ZTY32YXBybK
ELWOcYvtV/O9GUnNNKOr7REuTnjCZLUwVpvmQpAD/OZnXZcaeUcsYYvwrX2U50B8
zHlwKBHpvG/GBVEWkJFDApgqDJpJT6r5IEn05yHNwz6KrUaTk0ogzlFs6cAa0uqH
qU4ONPdlP1o0Mot8t0bp2toLesXYTtNGbu42J6Zr3Hf5fyolHaVdW2SrDKHGtBLU
JraZ/ZpOkEJXhOMEQ0ki01WaqQwKo9oc/thQApqsblvELhEMbODxf8D3j4DbwpJS
89QcZ2ZH9c7Db1oJG8FpizBqjFrk4hAmFn52jF5IKTjYpdbLL2rH+kYYb3jVgZj/
dmSVXl0b+oTknFUWohPxfmkZjkQCeTC1+gF8FU+tAttMM07ShkfLZqgYqbxBGanw
bQMt3Uzd3WQ3C1VPO3mcK5vCuFUMJnROxCUYIVsfmBxydxLX4UVKj0fQ8kgsKUMr
amrcm3o9hCNjSCkg9dUwWPIz9MaUZcI6wVcn4ttuynhZikxFOBRkVLBCs+tKsPd0
YcIKLztJPG9QUB1I0DD5JOBnLwGXfhQoMVzWofJN4v6EI//wO4Li0ZHB7WTwPFf4
s9y70v7yDt82AgfE4W1NWSoMN2jmxT4Zz/SnzeTwxnr8Kx8b1fO/R9MZaw4eH2j3
kPCegkLwTHIGVO5ngs00f0SGybMVyzDaUTj6veM+QxpFewI6EvV3US0sr86lZHdN
H4HSYfyoUQ5RIB3bbFTVrMBiFI3XwXIeOZhZ7eDj2qkWQ/6U8QwbQRmyGST2clxO
rUgdKKZEYNZ+JnbAAUNlv7ByeciWNrWkxn00WXu4nCLMRJ6g81p+ub4OAFXqsO91
atxPwrJe+oWYFxG1MWaetACCDU11SBgObDrjwE/Jxt9SnmIWilQf/vDTSxz6sxWH
XgujhJ0boldIffYQAqhhnbBXgi+llK1zOSP3FkEkSsneGF3JcaFtknEZxHp54jnO
cZwetnJyyRn7wLbyr0VBLYcfzxwqAsZ0kbgEFcgCvwojEsccOZSWEQrTM/X4Vhqy
csWSyOhXTHuWbID38w2XpkdxJeKjahN6Bxpf8TMHexHlLgFrStKf9R5zpaMiOXtG
zHmE71wdtSeU9BcgM+wHu/HgJbXTYGZQkP8lkMynfKMG93qDwyZRusIYJ9wsCX+L
OJ+myjHsx/661wEw+/XXlmxxjmTy/yv39DZlcE6fhWf5D8nzcpfmWFg5Zo6nsPP8
CStzmDfKTKWj5jcqVGzb+IqzNswLDCJ4JbIc9fwqf9baQ019dt9FWw0SrnlJooaa
5Ct65jZ093JNXCDvZV7UG41Kho3aEO5BxLbdP1w7JDE38p42XPIGJAbrOc6J6itM
rhhPKxKrlPtjsgybiF8MODBLtbVyMzpohOVw1LoLjLBHNd9rW6G6tKRHqUxATQtx
y7jH23kdGZsgw9SNcD8uyYvvNSWMcR0kbGZEmA16tA68jhm+XqrS/5rvmvnMRnSB
Tq2F7c11xpcJN53LrfdbqNSF5P+o4iVEBx9dfz9LSxIvUSyeEkC9JmTB9v7qAYJv
tWuAg8W/q9HDRCHmTDRTUiSZsrS+cFaX4hvEX1C2vMdOIs79x0HeEJUvrIkj6KLW
j1aXDp3QH7IfQ1eB7kDqydNddC0Vcs5xZkwKE5nfi4OlxIF0SV9OVzCZJW+Vduvc
wNqUvYY4j4AOv89KJcy3pfvA1AprMgJrdc1bmtSdB6n7jbZr9PTW3EN8JXLoZpiu
5WJY1pH4MYh0z/ISRuTtqMzdRST5FnV2fD0xkKvYpqFabAr1XVLkBaBYxnbxwq7Q
3YOAuzpxbzvxyH48MXTBxo6coU8oWVhaeNFPCQGWn2rQO8V5XVwcwukQfFZ3x+zy
KB5yX2dvL80wX0i6mJVlXMT6lgpmHQWUFkRFSezEi3uSEt5UKE0KxTjqZRlb2s+r
88TA1Wg7CBaRflPK7OzVIBL5SvosjG9ShJCZhfPtmYu7+PeYNYuUL6hUXykevAG+
xJmtp6HE2dfsYhYbAihXdSQPCZdlXUP6NixiJK0bgmo2cTD8SRgmdC5sAknwFaJ7
CEi7Bn/uwZ9+obHDjL6cIWSEz7gbGAM5kby7BqS3HrFupAfU4BuYt/jqfwjzE9k7
TaqOSyW7smbg6vO+PvaRGjFB+rndYgvJn4A2pFbQ2oZ5WtzfPhUAKlxJOVEMe1N+
dkZCBkNXg1eFfF17lhkk5HiZSeihg0Ts/jxbJmSv2mlHQBA77HLDkebSpX9JFMLJ
CpWfejfRVrFfJ8xri8/4uqKvp7J+9TBjm2AxbB85Txaoicv/WOi1EvrZgXFtv13z
tCSvLpZDQ07ZE2khFKc3kbk9C+bmBmXfF/+8T5pnrC9gdDDGn8HqXVEEC4CQdLOk
KCXdyupVZvteZPGQHmNjlARzWJRtkyA5ZcSP5cIYurrd+XhNWzfIPHU0xRb+N4q0
/Aqb6iChhbamh7E/v6hnzsr1ZAJUsgjjMVgYakk5oJPofbcE9pEXcA79WRMPFnI+
m6GTKAaELJFt+8LLEnt+5y3d8Rbzc93/tFXo3zQRdlsdUqHg3ni3csu8Jfhr+Bki
vFnpsio/Numn7xSCZPw66C0UikrjqdrgYkFipUce9EqEZZe6/I20LLSxxP9OCe5E
7qmGMHsZ34o0sZDO7ktE5VYiKWSfkKTKgYMGuWBbo9SEMFJOWGvhVLYvNqpuF2/x
LT/K3Jmq/koEvGqD/a4QvVVkkmn8AV6b1TMvQkWsjgLB7Qlu5e6R0R2R/x2rKDq/
Xp2MZRR6H7AuKNrp/t1MSmMmyXTOXGH2Q4YOdAfl3cSSWH6D3w9wH+Wh4O4A4eYS
nDNJV+k1vZpX7QHQv2S4tPCJ3qJ9sxywG5XUAI/zZCh8frZ972jIOjISRgg6iOYA
Jc4Zw4+OfgiBE2irPqD9SZrKsy1KQG5QcdptBfRiXN4wLqrvOZUyhkuusm4eRg6P
Npp1aGBTI9n52tAS127WFFZkZ4sr4YaCY85N+75Je3m1Zv27VkJU18QRWOHjQ5zJ
a7QN+3BVwj2DJF4bARxoputiQDNh+p0Xmt+A/GaGBK/K5ErJhONTHL0atMVtJA+4
k0dOsIby+/VYv5WT6O1RkHlADtgMKZOdGHSDI6f8H7wq7NWJPAQHZgPql167QOvo
HK1u9g6tUMVXo1PmJkT3fbq224q3AnZaHjPHl3q1O6nKT/rpflCNbFLT8Jn1fUXt
1fHqSoQLdQ433m8v5qmbfxMaVh1/3JYVFcHw8MgfvEqE8uLi7UXt4LSyYILYX9lX
BM+dMvfyV7PTbrbmWmod77RQnE9DoRhAIDr8H0xWkc7tM5mieuAlw2yTXhUKuXg0
Re3dsYw8ivNc5PFASKZ1NMYXrkIk85GWuIazsGK85sETENPcyppQm/79ZuEqXEiY
Fo/d4cS6jWP+61js4nAjiv9i1nVaLQi4YHwyev8IiVhtXe3z584o8twkNxA06ZuH
0RNz+Ufy/TOMyQRC5/Oit6rSFtfPG/GN8HWPVHAnIFbcHy4XLKaTEl310qNL7Aol
ivMuRNsCBc2TCf9Nm1KSHKT7c3tS39Y9/zgPD8+DTM/CoSJw7+7XaSr7KlcMOo8U
SOB+lV1okoGVDxHyI6wINqTmwXD7rG/WM/CLlg4XAp0QahRTnyXBEikNfG7RKG9Y
uCvmjeyJgrBSXOCiJ3UxL2RC7Nyl+Ai2UJA/UCcBL1Ly5jld+JXiw1b/v9Mtdiyo
E6C5HXIu4FVDIWd9Dhjel31AUjua+FDVOIrmYHwjKqTuGa/icBoRjEZsxdzbbwWH
w6gJJ+NW6RuxlL16yPTVuak1QSg2udk6YYfU3HOcWEWqK5MVB4EQ7Dvi/IJm8zHr
i5WIGbjhsThKfoPTtBcN6rKUZ/TDXqntfgMtWVM/b4X7ta4Hk1KN1SLiXJZOtAK/
k4kKko89aFKTwOw0T7fQg3vKJ7++kvjjqjDoV6XBQtP5wgdF/dvldXbVG6Fyr0e1
Vtwt81mu2lQCSSnvvC+RAVwl5zsSimbgQ0C0BgF4S8HnuSKcw84cg5vODmKPK9+6
rmQz9s/WgdnWVgyydOcurI7vkaMLkhQOGMTiG5uMVtS+WR689N9m7E0+wkBbBTgI
hqbPskOZeesG0vjKa+I7wtq3pCJhiiJOoHzEpj3bBOTLF0X87qbfvDnMVOj4xnhd
x62IlsFwp1u6Wp4UGi2ZOmGiaRCGlS0lcXVEDUVax02tPgSZ5p6ehvL53idWfCD8
UHUMP6ssElRjJkulUZWct2VO4zNIvVLjQ5qfTbyQkCXXcZ1lb7ZWpKGDqfjA9kih
oEMVQxtIqRMB4Qak3l95qbh53NO+I65oz3yHtyR/DcOlMi1IMBpVmp0454e31HK4
KGboULWffxLwbAbwVrVk/Dvtwd4zYa/LRzqAwWmy0tM=
`pragma protect end_protected
