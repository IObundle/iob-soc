// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
porlQvwgpktSLgzMcf+SYKeRQVDb+Zl6RqahJY7TNEbTnMCAigtSznHcM/Klp6pH
dZEhpNbk1v6VL2J9MNTh8+NXaVULhgsN9vrdPT824jb79EhKQkJ+xU54nvPLq2vW
fuGW1ejKSigW+/u8ZpkX9NyE2NYEYwPMGJQiqvp3MnM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12784)
OJb0KrCBiwCeq2lM5dX5cv6AP6Y3gHT0v4Ve+2QDd2ogWPqFG3+GKeO5p7bD+EE1
+XyiKRVFgHHDAdvPiqyrXuMcnhDOd4CiRXwTEuBhkpCZs4O0HnlmzD3dsRAr5bZB
HkcSqRUstOu5yZQIifKd13S+lVauWVNkTmGfVbjQ299oxP92jHhirdnGs4GqcPuR
n//PvtzYeCFnpwY6I2orzXHi4r/QAPqrV+GdFR6o1QWUgRH24m8HmZrLUEPc4rWs
mR+9HDzeTNL3tvgF4xhwQSQjAIDkRerCSc6q4RTXo2Ovpp6qAXjpwZH0sM/WEva2
7yMtPaDrj5j/9FJZxOtcpBduIU3TyhSDwwikSSU0P0Su84sGf3+viIWgMPRPZuxs
mU33lMLcGJITRTgvTP0YiaX3b98ErVGnPmzNIy6FcGN79WZ+QnpalkDuMUIdNVOX
E8kDwrtH1kX+d11fUOLqlZU0grTn2FX+xwH4G6OokY5Oxel+0LpwzEQCgv5KTCIF
cciOlgLQ0/KEJ4P0heJP7rlX6I2EZ1IFHVq1ez78ATwJe80zN+iXtkKXw8Y/+Fps
IDjsq+FBJSeIa4q6s45v8B6FbsOHHUL78fdKlurP0ksrCaip3qFRXySeI4o3UJ5Y
FLmAf0wJmn8qoqunNxN3VEQbSfBLCegZ0+oSA9KZ+SmUzSfTHhxUDy6jt8lM5uZ3
yuR+TfHjamsLGhGnNxzIpj4vpotg3A5ENE+ax6iwO2ZNM4940CEyxpY6VTgMoySZ
ESlAqgQ4eKmE6rjXdHhUuh39ERAZDN8x8RQJfgoYPTd6KVdmyPfl7VyXI5lECyBv
WuNfmAV0SItYDRhRV1iACJSTijzZEMacEfWomacnY2y7NZyC/cwRrkAExCkZ6qDV
tyyi2fZi5jNWTHQSKRa2txAuM9FnB4bS2vYSo/CAKO3YA00EWwrU+LXGsprGclRK
NFOWjowvzLPmoW7ej+bc+p/vZv4qlEfgsAmvhOTw/rPGMmM05ZjANZHpB1J0EzId
pi/9cw0OJLzrC5XXPrtZMnWmggw9kCQYh7nvfwLayimVTI+2keYhFgD9Px+RJAu2
3ssYWOOgPwJDZl516aiosgpQuWCkwgklf91CHArmGYaPA12RjD7JHEFSUm4QSLLt
fn59PFy+9U3Mpa8qN2hV4F399bqfdSdV5gw3Ir9tVFAte21Ys6hkTYogotg45rsJ
l2sfVAPz/Pys70gIuN6jQdhMPGKMGnzGmLweM2t0Gq7I3dzIsQK0H5sW1CE2cgcl
a+EmDAceobMJrUAkp1MODVqnCl01ezYbH5l/tEPLXcWUoxhOjCNJcO7tjR1g0yt8
YKBuE5YiB0nhjkI1hFie3NXxbk4adKexmLmbZ0x2SdZD5oYuwM8MKCJMdbFmlOvZ
f6SB/CQs4/7Os/U9NpL/K4FwEJQdp547WDoVg0acXl4jQ6hCPSdWuRWhAqkYNMGY
cTRJABYTb6Wro3G67LQqdPr79CgxRDVlO3gth+rdaNYedxM7txN+Cm2iBtKWFmoU
IV2WVmq5ckXICjf0tkafYoDciWXkIR5e3CTe2HgS51gzYcWh2AQfRq/O6SmTZUAR
J/EgZPLqGtCYCGBqOagLdY24clsXutmO9X8bbFgJeJfoBoC4K18Dby9mt/Dh/5cO
b9iAVRzZ46VzpXYc3RkJqEUWE4oPtvwSdBQ0zeAlNN6Mgqt30HH9rGu5EdAovJNQ
BxMr40es34M2cT71By2M0vPP/9ItAMfvJpDhj+TSpI4inxD+b1vbriXu4HUafunp
l6AFD55xhtLJ/kVYnLobO9CwZinZs0Wk4ARJEPv1mT4T8eMDCyCXsil/ZlB8w+bN
ajynEZY1t7bhmpgF6QXLRBM8QooJe+xkumDGpPemoLfAzcwPZHeyADbwi8aU41qT
N2gEOIpdbjSPdbkpcwW963WhJkEl5Ho5KDqEgvG+pyruzgYomE5NeAhY+sDyJJmn
cPQ2Zmd8mFcZNJHnQ4SeUSpp6QR40Hjh2yB/KlSH9mIHhx9CYf11nNK4EdWqxESN
oReLNDbXDjqkv3I4RU8rGEGNeg4VVqKIYbUxKb3C7rQmFABNlJX/ZpEfYQBiqSut
qSOXcpucXLd2Si9KBpR3kOeDns6AvWWH6PwhccjI799I9azTbhrngxc0OOX/MEDh
JYlzciISX15NBa1fidmYJ3ymysLHYA/sGVGEFr5N4VGhj4J4P8ktvrnyh9wwoq/B
mg0Ub8IsIz9k8+Rwd1AmGCenr8bBOqtLk0Huh4qDqfTWGD8qQii57FKewDZM3/jZ
UL8+8Fs7YfZ9RZMCYKpRuKhGl0i8Tb81K6qsPmUkqNyl6JB7l5KGIPw0lqrsr564
V4vkatRagXRuzFdsl0/gEs4DP4b/Z0UU+IZaqWxjwbrIy9mhUcJQSDgHZJKhaA8S
X4y9uY+lefVkKJQ/iLS4ev8mrokUUMo2AMfgBX8R4W81BHMacwOYVxDrWAu39LbC
4IpOyUIhrJZjSkGqa+MHBKLelx6e6/lusOW9VM5mdBrJT6tDXBaLfzudcJDlwIOf
Ur4zLBCqOILsAvO21/r11/giaVH5dJVe1GMTs/Wfy8uta/PJLF/3YMY6f+4wx46I
EJANGasrIbKF3mbRGZj3b9iyEQCQSG/AUnIcgfhjEFfc4IFZr8ac9uXzjzljRnIo
cUBIZC7TIcCZFe9zJrRy5HhONMlr/uQ3UZGFIWrEJU9pl0288rXi3mkxYrP2nF0d
5PUluzZoIFIlMtecU65BMnEFABuFPnDnQQcR8Z7MN1VYUWtdYn7+3Kx3uXlvwfCa
IIooz83RixMhFAszfFrIQBVRnkF4q69S4oAv4tRwfqXiVXdMh3hvTLbz3LXyiKDA
aHN354Cvka+tNkI+biTYY2DaXU4kyjdVM6uYyfdHum3QOq+SMSm0TIIOwLz62qEv
8X38VWBxUq3O/bfXu/3qUJJJU1gMW8VD+TT30yfGWkxhDxKPlKhthOYrs2w/fA5Q
LEnWDVV/Ik/pEoEcyQP+OngpPO0r9YhHSa96Yuk+XhMBh7FJnO602ovx+/9yDzEi
VPmJIhXZEe4kPdiVP92vzXExsiy1WFhv67aYsUXZEnQhOZRb74QhapBvNM2b1Lq4
xpTXl20gqac1PTxyM9c69lT3PYc7suzZajavQoWuYtu7SWrH63z2tFB/NjcBJa+R
QlfCu6X03Xektp/ockjHFhMEntuELkRx0MAGYvZTGMvtWyb89YbArKKpEECNitpe
2DeoUD0SDPZkBUpWpIDLylurz+4IvoOK8aUf0nR+aU0x1IwV+a+EImAjF0iYM3Qy
m81duXk/kFedXpC7RWDmLaXhM39jLBzEWYYCx+mCsOB6ZR16jFg00GfpQjbsKLE3
ErS36wWBXlolPmlio8WNsH+U9yPntL5QR9i47nn7J41EYsfQPNXhJcfdZu2n444O
fzy98rP2dvuTOx/9aWLUnL8B1vpJFzUUR7O6CjtWkJGYW+NwdrinzkshDU5hYmRn
6flsT1+ytOCuqMyp2lfpqDvBd4+fztbrUwQstAjtMAxA3OmEgT7YvrD3f3HPIQ0I
gOiVLCnUdMNvFY4N1HNE4g5FiBYMe4zsOc6MN0SoJ1qr0cEd50e2u+IKpNguO/B4
Q8YZpAe6YPdOrzee3ls/U/Hdghr24G3HwSvv4iMADMv7Ynv12lT74O0n1FTQMKjr
sN8jJ4CZKWMi3o1X1xQP0uHVP2SwC3fdA10aMbSchzuqWEnTqqFt0hQ9RK2JIiWW
AydrflT4zrSaxd997rMooV9CPIRidcA33SoOSB1uuSv2be9VwazCGX7iIKnyX2rL
IJkTAquKpneZ52rQXgptK0puwb5NdXHq6YpJS4oQ0FnugOPEJI7UW+V2pDrzUHwb
CG4+VITVI/yKU32HFYhciN334ZYuWNkpaFzQZ2nwCUwSKIlPx21hakGBAxsC+Fsv
msKeRT/kIsltHoNeCq+Jt+EnZPmkzANrVLrOEjANLSuaS3mop2FxxBD+eeTVIdWE
99DCqLBdeICrRXIX17LLl7POY2KSKJ3OXwfeATphuhfdvkCpM15gskv+W6r/t3qb
7GZ+llp5EhukT/NKiTZZ2CSNiTUFOSY0nRDH3b3qS7jKjM8Dzh/b8BxCfjShi6w2
z1aVikq5JRzqYpmjs0AlHLO3jX8jSljVhTe6KxW5ToZkZsMftJGMK2jGMmimnDNW
wYUVMhy9X1/L4QHNXmoapOBhyet7uKmp15uKY15VZ80IqoCf/ya2PLE6bi2C/mOW
6c4VhJhaxpkq3uRgLvpm4aNOaJ5xPImpZ5c9XeVytxnH7///0Uql/hbd9nVjDdUh
Le2bufcMHifQALPa1puO4WXaO4nnVMnjtUc7tQg7H0aoTT4TZqQU6HttHpK+eTRp
uklDO9PbCpcp0N6CMX/HFFyiFyAHAzkvVVWAHqtg5CvGZeSQVd0iMa+J6GLcQqQU
XajFfEb/pkPV2EtPlqprjZMV3ZWLj2OuBkszTbGNHXVYxwb1TJKI0r1FoBZTc4Q2
fY1iq3loqfvFO+rQBST8fFPeVpxETgXvnVkynrpeHY2paAz6xZ9dmPRjkjKW45AZ
g5dq3MzVRQ2Lt6LVyJJbvqV28V/t0ywhAoq0KLTVkVNaUtI/zd0+bPyFkunrQQge
CfiBCRc4HMToGiGTUPlUPhfCxOWXjNq2K75QbS9Dbuq0nHuNyG8RRY0ZaOblWbCH
q/ayI0zV6MkRb851DTIr9tlcg8pV+r5i3u9SwizIMihDkcit/YnrUEh4LwRh2nQ+
eGbkD8oT9TO1zOkk+4Og+B4RAR4WzXTzyPl4D9FALW2CFUUCgpwO+sbtY99aHSZJ
3WjqgcJZYcRdojJct5jUjgIPcXDAjrVKZxlvm4DDqxPAWG+smEfJSbfu8qJAWjUT
2pJ89w9A+edPIX4tMS6yN/9GBQ/EBwC+Jac6JTh6gl1Xx8y29FC77oUCqiYG8Bji
UX3/boWYRBCZRKzPZSwxL+G3/5Bm4+Y6BiD8iqEtcXXr3aCRvej/FHpKIYAk3Ww+
vmYGJw3BbxtdKnCmTnecMuti4cQewSYpl+NzXOku5q+bKL5hsxNOBuWA/+zsWO5E
kggOcxCbY07G47fl6aMwbUh4YrYbbW9K8J2i+pMPPzNl3zCQpTiQV2Bm1USDeEtq
eEko8mQIuT4wWAZ19I9MII3WXfGns1X/RgLgok2/RWiqv/dcLHlYJVp0kP+zicMw
PlV/gtjDdTGb16dRU/AgJsrV5TD6HJlNn2gTlk8gW1zJnCXYUZM0dIyzKd0kZgy0
L/uRUaXZ4iEyvMW6Txz9i3AfMbEN+wSlWpMBn9ExaWYCHgVy6QWz3g696XVQEtaZ
eSQv5NYWMOOxz33hOWrJctFHlgGdLCVipBz5qi/JPB6pCaVbszUDS9lorJoBJgvL
Jsunn35FMSw64D9g8z3aX7+WZqW9BIB5fA0OeIobRwvtinTe6FNGw3giLZL7+EBQ
KTwi+6j+Eb75PCzFDZibiL0oL3Fo5Zu1DVm06YkyFiEHLshi46CR1TOzkdvMrlYC
e8Z23iQp1kXx97G5WA3FmjQnMr/4qIhoyDiObKNGMyVIs/6tli9Za9fjRlN63Yh0
zz9eBOEQGbWxOdz5immZe6vSPLnzOw1SMP7gboi7i1Ap/Fwz2Ne3hafTMH2NG3Gh
jprcf6Ol5AZmXpv/oe+xaEmvToFyGYQmwt0aThQnfNcBT0F5/M6y0nKEXptoQgiz
wDAWajOBXp1sdVf1Uh7bjm/D+BORgzB91Io4ei2Ne8mnzC/SlxXabkpTwuIUtsyg
ZGWewJSEWt3l2v8hOVQ8srtIZDqdqCGdkTjU0bBiQlGMdwAGhTADHo8QQpTTUBMU
plIxCmWbt4HekC4z/45o0vkmWHUhH/3CkQXiNUqJHMt3mLZukXHhnynuFj1zN386
Ca9qkOE9LNVSMA9wI8migY6az/peYmxbhcphVgd1gdjSZtI32wBfJ5NofhRXcR1P
otUVDqi++/5NtOoM/PYEg2OI2ZoJLml2S9tqXjpl91duFH0TWNrg45Uh8vIG/hNT
qgd2woYelpqRi1ZMBYh7mNlPwhAIFboLGp/NjOipCrscT2oxuJsvYQYZIM1AO7QZ
QjNkAFfjAoBpnYTKlbI2TYlQJhgWeRwAWnyHu7w9DTFhCXWnGgdZtlHOfrW28C2g
lUNJZ8zqWai9PBoS1v91Rpr1woRGgLRc1TvEYjzMYoABzOrm0ZC6Od84MNWRncwr
/blgxF/Kea6dl78t/tGEZly5sSVuRTc08rmpk60Nknjd6WXE/R4gt1SzfP7Qi/H7
Kvs2AV71jBR/NHdzPcbj6AaQ9qnWG3H9rkD7RjBxOekaDVxOAtVM1AiD3D2kkmD9
vRIJuhJUFgmvLeGicDoN1Vr+Nh31CVtPkKYGaYmTwpyfdlgoJJn8KtoXNCErq2G8
omezGEnEQxsXGn1p+cqjS4c/Ft3xD1FXQ+7kpfqSOYBnNJCdUR+cluDOm99RA7ok
hcsSxFjjfas7D7B/zpA5FS6i4inalVjGQYgfZstVWV9dl7rm0Qc/nV+/6MHt5A3U
R5O9sWtjLVXgzG46c9d1+1LtSLSeITQUZ/9mdLtVgwa6NM0uGrIFtNkUBzH5AAWU
RR2fg+UqQe67fzq2qC0baAzEQJ0SQv7W+yoY9qayzwdpK1vpUPVqPUwqUq1vkeSA
Prv4kTkGErgLHchmBO1qFUZUS+NSQ8aRV7VUxWlPrD+dL5U29XzMQGGr6EZEL3uK
HXm2xhjAhyVXOC29c5ZdlRqnaGrUU3fhiVCzg2j7/exhcLqzDRQ8g3kcR/hMFtyk
p3V5ZM+QLA8vQry/Jd0JWgNYupf32W9u4tTQMJb/LPUXjIlD3PmDAZngmV3687Op
zHc0YK1wftVgr1/DCtcRQA20eWvsuntDdFv80//RJypResjxnCGjtak0j50BxIia
2RW46gUH+YHhkiY5XnvfrVyZnrQU4lCehl5wz569Ono/b89yzEt+eMM6eAE+YVjr
lX/N3x5XZohN1wTc6ol2buW+j3eaD506hKr3WExanmzCmNaTyTvwmCe8UtGhUVUU
8qtnaxazqrucY8HUrR36M4fDf0pl9ZCYVM8CsRQAintAJCrXgUolEqKio4jvv1xZ
o5qScpYXoN/zbOVPd3Uifa0lnVDIGSvNh/EVPZolHuvtA/LVByR4ZXrL0hblF3zV
VvcjdYBSwiAzwoihq+9RNa4wUMQB0gUgl83B6ftc9Bi4copmJUHt7g5qRiHc1OkR
F509Og/D2BekkYIoM2ElWOd7PodB/RlumvmAeblV7bGYsDAg7oQ489FJqIvhPvDp
v64w/WYUUCkwZ0QDNKmAapE1eXgpn89j6PCxItBqJ5ihWV9mhBxKynN6ZYFl8yr1
kpWJgokffMNij9Ox+XbS4lN/K2rHjjkjtlUbT8CnZy4YMT0LNUmdhdS+uhSPfe2d
KluaRG2dMk80wPlV5P5NDO5iHSmbNyxP0W3IKXZ8lJaMwXmShdJ3ofpzTnXloRje
dwu4cGmhXY/xfw0ZUgKT9OuVH/a2YsWwp1cTaa0KbRVYS+C8HeHTXm8nABFGoBIw
jIICO5s4BqdyhGA/NNspqFpFfcjiQPY9EPP+btUq0R4O7WubvEo+XfyiaSHaDJ/v
tAjZKqaIhaLPDXjknxrQTNmcn2oihBPpUmV+pGK4u2NjF9iIW1YgzaEdo7WgL+PA
1Dx2awNvc9POSkJni2TQaT7D+9KmhiTLzPtDUY9wQTtj3agDSChg1kKPY8/9vi+Z
G0XtMQSGFoTRvtElzXtx0eOiVY665it8qX3BMMobpXLj1eSHR7r/4AbTOqCFk78P
LTcOFTTU8OxL8Zx7gspxT7fntNgknrwNQ1DxBDIpXiG5zaNuHnoy9GosuBzyqoze
sXHYC++lDMfugN26HkXjoHqSxRSr5+6cmtImzH+dTv72IO1n6Zc+Mhig62tJJVCy
0W/hH3rieM+diGYTJBITeAFK3UphZct2mZqadKNSO5l+uyAgCWHwJlPOrTTusMhC
pcFXp+p8Ohd6r9xT+r/pWm/5bzuFf6KEU2zPLyCF8R96hcrs4EqqHZrCc1StCelI
c1JpnlU6RIDP/DL1sjsxFk9C3YlXBLsZeUDmKPOrpCyZ6q+/dcPPSxVenU67zfRY
G5hN9EaQIVy/H2T0X1G5utKVtWPNnpTNqV/6IaAdQgRDOpRmd6AKJIhMak/X4Z4Y
lYxE2sFjNYq4U4L5A8fOgRoF3CulIEQr6XfnTQIHTOtVibhz/k0J3DGFKI8fPGzQ
oGej/8ZTZPLqL29byHE4HqYpBgXZRt84iLcjmowchacekJe1SDoEocNVgCI9u/tz
ulyYVgpP/5+bofIfpu2M+vN3D8lAlab9fT36wNCbD2MZ5fqD5H/J/Y4rHFpuyVKo
8KT0dHYZK7hkIx2/DqPt4PjFFN7MQw9yCXnmdE3nvy7gHg2Nuzu12YTc7MtIugnt
4wbHc9Yjmh7Ox6lsYxEwIfzD1sj1j1lUs2u8h6hp/1nDUvklhOPEQPzU46RTSaHe
CQnlxZ0ecQ/j3ZWBrjt3bQnh2ItBL+V+l0fWP+ediXbbArvJxN8e5WsnNHD+INf2
PY7bT8378jtWSTsdTXAEd7ov0+9I3BqZcCujpCZsAQbcQiuBXezwNkcp+WaNnVVF
z5ap6koxdjkvjuhYbSIdOIlyhCPwbJW7oeZUoLJyjcuYuQHSvbpC9YQkXiB2zRKa
C8Oi0Sgf+5d8z8KCnP+ZsqXngTe0wAQkKCJ83D2vdj1vBDKVq0pxkZ2Dev0PIW3f
5qbKop3ADvd9NbYdJPGBZVE9VUoA5f+G83OMKKnKnFjNZa8qbvqLcfbR+KK6+JVD
9n9/wcxrNOYkIB7XuG47IpQQDQhlUQnSh2JZagAAuB9rCzT2j9/d4w/S2Iftceo0
RCSsyvavimb25ilZONNoQzlef8BAMcVMpeDEGJIYw8ProPxtOb8x8N28OFcd8lMu
C1URfV7RHLg1gyoxSm6BoDYKPPpclotbRwRwkc7f6TedebuS1WSA8/ojDKuSnRso
Q6dJN6+huA9sHXKiSw3prIkzvPhwXrcOULk60unvPRn4POqa07A1/b165FvQBb0D
qz9OUMVAvD1/753u6fhb7TmIfPbYbo1hkk9LpY7BmtWjhko8F2NWbfFdp2FRbznx
/Ih5zB5yizY8A9r1469kvzX4PS9W4Bqs6QqX/TahmRgJgZA/XDOQ1JFneRjTUZfq
jiIdW1/ubBaa0brvf+SHwW+wcJlMav/A/+gOG1by/P53BJkJXwvdpc3mz8QdS/3l
iQCSj1qz7yaJt5a0TZe6We4golnxDsQMIxJ82RNz55Oy9TZS8F2Rus03YkUd9yK9
honwxrLGn1Cslva+wM4f2FGItmf3DxvoMwstFPfoKjO8tcCcBBm1Zah6/P8vhZ6a
M2MqlQI2JPE9Yw85mSLGs73lHaUhwW5JFvpJulqNIWI9kVkw/H2KBxSp2qXj5l3d
g08CnGuq1QuXl5V27jN633HPrW2E0o8hbz3drvEkYKR+zftAt1eWnz+yWIM+YqCy
f7Th78PySkchEfPe310mKlMWItaGzuVQ/pKYCiqG06LdMxiQiOor9P+ChQBu+KUg
JUmRSbqsVOHOMMaQ6B5CnzmxH10PCSVCxIfUbHGOEH9CTEznvCQ61p3+nNmTtKBx
CGyQOLbg6Vtla2avrtVn940Sy8FUJNdefQjC2v2muFWfsbBV9Rg9e6+atH+YNCYZ
yzrtjp2edOvopHjY204fhcbblQtZ3sCxA3hEmAluMBGhkjqwnIRaJ2weIdE357qg
0QydRhD5yJmWf12B9hZ+L3xvN5c3QBGaUKj6E98/2FYh/i39Z6I21szQD0V8sDMf
u4rriAanVM4b3dpWWD+nxr9YCJpba5RS+TuTJMovyApgzgUdNebP6S793QvGNGtJ
wnyJ+ytrN567Ae48YpZfqv2EPx6lXUfXxrhWZnRpE9TOo0U1Qu/+RgY1WTsCX2sE
jG0OfI8+XLP00IP/AfwNS0nz2T9yStvqDz9dQn+i75o3vQm9M66BYwJ5G6HGf4Gx
Bc2KpY0JUu5JWDq5h4K3wtrsYCBIerP8We6i28Og6/NO+wgJ16v0Gn/oG+ZhcQkG
0ZHOM533ie/eytKFcXHw+y4vX28NWkwPyyl0OVdr4ICCT57hkqVPi7kLQgqEcHgV
v37sEk3U9DoynZNbYJywPog9B3Ets27PuA6sVDLVTfyDbKf/OofASPx76/+ntGZz
zKFGutgVHpB02/SPSUxEHg8O6RitX1OBgzxrwv7nGTlnSVU3sKI5HoJvcyrLFo7z
PRNQQIb2CxDwS8t2Afj8MXLFRm9IdvAIyhlRHeJYFowRDghM3mxLO/Gc+LzehMZN
lL2gLf4f+ehoPqqhqWPPd0TTdMkfCuSr4NCznwGU1Fs/HiwbmPel/89dkKITzfJQ
+PlY0jwvBbGQVnMAWGUOj1fIikgzinMBNAO16oAQcovAIEvOA2QoduJiQ1lIgcpM
0bU01WFRrhc4O8DVlAL9TBOHKbBKW4bn4381Vxq1lASOC0UO5xmFIqGGgU/thSDH
ONIHTTKnh/EsEGPLx0rRaI1luP4JCD2ewnjDEJFX817l/DZiR5acYI10wExJsxZg
MJBBjPAyOVTC0rYlz6gjfcDTAwIVdoh4qlAEWOAgD+eOnSwzX1Fyv0K+VmMRXYhf
p7T91R19Q6SnNTZYkTa1cRUdZ+eKvf/UF8A+6Om6zE6pYegTNhTDTTbc+e1G94+v
HLN0uGlGfgxk8s+A+fA5e4/M5NBtqAzUPEhfsKB5daZREpLimPTlTst4TiTMN8iV
NdHwdl3NP9OVLfSFt9CV1Dmrlcuwgg/yeIhWS/I4NJ9Y6unC4lqqsmSd+dNoUttF
CTv9hrRLfsEaGNZB19/4/I5dOfuZ7+YwMJvOLWogdWcT3js84OEnXpb9ntPRhFY/
YBI6mOfRztB2/d/esTqwuUo6AWYOt0WoZwcI02Zgi94UPjVqEDT3FP4kCZ4rPgp9
Vk0wnM0GzGD2Sq2RQ6OydIl53q7nfZ8jYlVFLXYPUqnv3DJKxSuI7NI+kvf6b6Qf
qx8SMqhdK/gcnUiURffB9V87YQl+YBrT1ne9QqjMtImdeoXu1EWdWCg4ZYa84fr7
rhjYvzeMrssdnENLdRhinkGwcTS0h3HhRetCTqehuI0khIAKK2Y8qCXvONncdFtj
bEdO70z9Iv2rXjYC2ird1VbpImecl6izYfY5e6YePUg9XccjxKmuDv4bD2ik14xO
hrWx4BDwm05c+fyqsioKPBniRaH9TyMETgtNNRnQIQhlMlo/04lOgRJArv3Uug/i
uLkitjUH7avIOocrSmvslIh+Z4VCDVVigH6JSIzDkeAZnL6k1rrkGZ6+l3aghP7K
d4BxdoWT/UO+Oyo1GDH+tRLx8F4CULP1mZo3g5GAJA9FPICJXD+ykt0Nt/cgQEMa
vs+37gA0/ELKChziGPbg3ngrF4L+B+TJTob/K7GqpG2RHI7D7AI8/szk1BSxJg1z
bOi81xQZsGmP+r7WuqoSPAQFC7Ad2DnD3Q1GacjCXZ3RvCZk+JgzlMVyqPHWBmo2
I0iXeTte9yGc4XP+IWmGwFn7PM2L7/TDhpZ1P3mRkyV4wSMSG4irREXsf0+0A2oG
pi/O+d577whWAwzWXHxm1I1dyUJk90QJ3/u75JcViuOoTXBew1qdCE6mOpQRpjYw
3bNL+69WFRckHWP1Q58NCnncnzdk8eGUlIBTQHDbLUr1zB01/iFK1e3f1bwBHKBl
EurOROyjMDlU2eLWTHqHRZvVYGk4/3xTqs6RzrCRweUrpOnjE3xHi88xmvJEl2UC
IVTXTTeoljoTS8K5m8ulFjxSG2pDSjXTeWs1GloGK1IYEKlCkT1RoR2leKiSYEFZ
Og8QH4neA8zW42S6J7tm5CLH4XW6rhCF/d9ygDyDUNZJYpKThO/Hs3wImjFP22f+
gR/EdKDwQo+ZMnJjLxhcEf26x4bgKIwTYrZK8uoGuiPwKS+lUG8gGq0e/SYVfsJm
A7IscMVyP5lB8VzFKRogSbdy6FEl3y4KK3mqcYGrM1rcNQoRhPd5Bl2vYcBolOaR
8CF0KBmetipexJEAmfCTlra8FIwQAARCZWVrf2jKWQw4kHcLw+BylCXncCEUV5kL
PgAeUy7z3m9gLfr7IJUSHR8bNT5dmaKnkwSbeNCgpUlEfIRgd16OCJV28ByKxSdN
seN65OpHncZjXZpMzwyLKusvShyrre1lxHEUreUnOQsGhYtkFOReGg/izz8Qzcyc
ZoYVrCemd76axojGtREI5uaAnWXWi5PaXlvfrgRWQlRdJFuGzSTtamVLtMTizRnx
be48EbSI5Rg0Y8lE03xpK/8uyickL2MkrX7proUugoERV8j5+83zb/SxmuCKGwgy
/teCCynlZs5W+E4rjLLnK7rX1PCxI4xuUbDTJFZCBf9tTIO2JAz8OtKb9cjTVGiQ
eJCoCsGmgfDK2z30ZvC2/K8aOkY4w28FrG7cUHqKqs62cQX97SYssBHZPEtcmXzT
rimAUXR1e4OXUliqH5Cagvmwews/5jWPvWJET2mgde85lVC+PpA90YC6X7kRQkN9
atWAhTwqQ1G0bxVsqPL2X+kd2NXmVWEZz3Pe+DaCuFkNfKDsiV3tJLaSVgi1RIVE
vwldu1AO+pMmtI/7Nf+gjmOhhJgVij3grfcPwVrC18+42HR5KvH3L1ELNaG37kEr
YuLeRFQEB47o9tKHXnaUFE1FJss5c8+uJ11HfrDZDO2cQtY7Y3qhmVB7iBG3LbKd
Z7nk7rpIfCMu/+Ho6nkCITeHRANJjNEXwHjQHCd4xVRajgcHxk8xmG4TycjfESiZ
oMqcyI/5jNjxyx1+XsbPNCWPoEJfQ2KfBP/VBYUP6wr8eGD1boxps6l0I2MfxV4C
Og00kviHrMBOIEEAV/nnE2HWoPcuNr44PzAVBnFiSVw/UAxCy0IM+bMg2PfBuz59
9yA8H+mSM0WRpvXSFW+vCbnCfptfj5ukwSmmo6FHMDU5cfsIIus+nVG34nLtXhqh
glRk+Xr4aVn6GU/rsJ1BehmMOv/gevPxo3BYvq8+3cl6Fci4PzrUKFMVdGFwOiH6
S0Tovw1XoYCvDdFLtLVCVrkWjT7i4R+NCn2EW2QNXSFZ6+nlBBGd0etSFjjpv6+8
ygNRhp/do1B2xPccc1DlXH+jpKwOd+9h4KDQMJM2f2Vt6nVFVG/3zoFQv0y/OVjr
t5fEa97jrm3/04QMdAYxHK/1HbPaS1ZUHhPFo1b9ZuoLnEuQzLyI5nIaG/9ueCHM
HrIXVhT2nj2Szi+J1oFJ1DKUR4mWXruYaSPGnar7vmx9PLk9Gtp/u/ZgKfEVBVve
HvurxD1y4/Fqt0wbTeJxo9utmxih+AMx5ArXtfa0nI+UPgmYgOtVFI5UTvq+/ESL
vlKrb9vzw1QJj6Wg0lwmq4Ia7FsXm35HQ4wGKj6+qragFY4+mw7+3hJn9OI0AR99
la1+fKxFbmcOZ56nEZNo49XkeNCpVorGydDuVSaMAhSE3v2do9FaVgtcVnQ2kshq
QQFWBBJ506sYCLcvD5wcPdCOGj8nwiD3Q/xOrjG0k9UOlHFvcZLncd2llXCHtgyo
ey9HowyWhiJV2wILZbVTA6TC/zncC/i9TlvfKdDkYhDw29TJnjrwX6Gl5Y40E8uB
pJIVlWehGncgerdJFYMZuIZYmM2HNwWcqu21iy/qkMSvG1sbpyp/yBF+z3MnPy7B
RpVhKhfnCwRYCFCtExk5y9AOELaUhiQAmhY/ZScHuw1T+FCscM277TOaLeates8p
O0T9xeZa7zc2BytBy393YoYlwNfQ4ensfLTATB16wM49Td01Mk4SkSnURvcUxOGq
GAwYktA2C2rexp/bcVBAzUAOKbuxFwwlMNOHARzq3HWpEvT+g/O+N6YFwCUyBGni
9a5bwQyk21b8iHyzKiFnvVRy8OW3wskadrpOucVpfTBmQsPNi1iTPYqP46TWi1yW
9M1WlzdDcxj3tbmq3rxFTB/7x7WfI0XLCipVVN2AMKN3yJ3gcNqfIfMQFAsuzbs0
OpNn2MjRz9Pxin0tNntaRt70juCUJH89gHGPcy4hm2DWR7vneCnLpkV8kuSY3q5Q
LDCq4LY2Hste9Zu9g25K0HwdmUs5W7CYdu+UOKeUJr3jVD8/EsJ/oXYCNI5G3ARP
37/yY5HPjPSvwk8greGyMhynCPAgJeCASYjrAUdCdUGabcF9O4UefJez+f+2jzeS
G7GxTEUV5jn7AAJwQIb6dzyi0fwZe/noYt4+6KV7n85bKXLaNpis7nIgRWMyiM8g
X7mAya0unw2zj2RsFAG14ce1eE5uxgDNxHQ5uThkNgeyjTDjSw/TTFoyfH3CUHJc
YKCVVG/84VYR1vx+famAHcbNhgrgnsdnWo/J5Vr6tIxVVnFMXKmGDKfXxBvLZF81
33J6XoQF3nuIyqwZg5lK5+S48c9b7hMuN+hzxBF5ygt94ad+j8K2Bdtcz0ii57iR
/3r2R7EFOiLa7q4cKnKXrpL396VIgIEqb/FQV+PVpEz1s/29QJZ6/b7JHO+U0SSB
z34B4z+9rJRaxqR0txvL9QDH5UUtBb5fjxcS5TP1m7eH5F+eMeoYsVaXOikupusQ
zC4HK6/bPRma29i3El/DJ7stHcXgoMoQ2iD6++t90LcRg0TpEZlCYKgPFZNoH7dy
PBWbUADdRXzt8f8/7p2aqcOHTTFG1qRq7A/bWginJx6R4pk/eV9tY4nzU0n05FzG
TvfNf6lNZd8fdaVDi8FQcWL1gtllBi6T7cq91d3qU7i3Q+t5wjLoIuG4lCr/fgNB
7FD4/70aX1Wtm8yxmW1Upgz0GR0RovZcL+mZmLndYUpUeyMjZGlfuKlAyu3wG6/8
JFohNm6gzoxBD5rTMNwwWE4M0uXsjEIg0cSbt1ep1SU5UQXnEwt6Fo1Bsa1ef2ta
bd7zYGOPLgSBEg4RSTFfm/Dvex5HEMXo81Vy3NHBLN5o+/iW8sosx2NcAHk1jzlV
H/pyWBcRiB/VConxJETTBEdZXs9F2jXnqSggxgKSfp75sF0rZcWaBVcDzv65mFQ4
DpV3ebxCWc/GjcH2X490BrsRJb6pUUzKNGnDeq8g6ArQU7KcWmSO0s/V6DIt4n+1
YH9bUM9GlAHq0GmuD+zGds9uWblgdUQf6c7EsdhaJO0kFO1sdbus6SoJYe405gj/
/3SUJ4pDwba3N7PU+CLnRFtUaC4hjnRokb9m6qusIwdGehHn2T5imF6fkHejQ3XK
/3ImS5rl6VdQl8Tj5y9I0Qj4YYVm01mguFCWMzo3VS3sxoeGYZdCkFnUmLhsv6Af
IaYJAa35LCGGWiyNEA48eCa0wBHeXuL6kh3KQazXz5Fc7pMtZz4pp+dsMtzDzhns
Jc/YKsIBBeLzzwoFxp+P6fX84ZzPgcC2+41jkp/LUVanZWBhyLIfRLgO80BPUwIx
fve0oA3qUBzJkQxHjTEM5pnxD12JeucrNEO0/SoyHW2mE8l020LuDSB6eKEyFeCl
5mS7RgrVifj5hf40JccaAm7JWDcAVWDH37gKRT0n/Q40pyN5SUk6HG6S5utQjZkA
1NBOfz15unpOkTSzc5m9CBHzO1x2AISIIDVAyxWDhFMZmOekpelWMbabxkCpueZ/
FwFzk9RixTrBwAUIvF77IB68bRKYtxu9gwsTnTvOz7iAseWwxpSiBzQXujazWCA+
CuhtvPEl4+438/T+dUT+tQd4zgWWHCBdcYLNB9/oc/bfnNUihIfh+wRb1FMJhqQm
qFgDhzQzQW6yMih007qiktn+y42zyd0YL1I+vbzc8ZO/7vpPQgWASZVmSsqB1+PY
4YT4d0HtmVmc/cZqYtV7ycU/CkTduHVQavpVSFenIV4gqQuX5rl3s4hqHoJWTVaM
Dp+Ld3OyAE0VSWFWMupARCSeQgElSNrwpFTH+X+PZZzAi9EsJjRY3KFjuEhGhzG/
GDwCXMAR1khO9JZyKFpfktrYOVpEyq+QgFEZvxJ1EXb5++2TLtxXmirCUFQK26DV
f65ILgWcU846Mor9aOkDQgrGd23zEatzlrp8/KrNipm7x0GPg7XRosJ5bXlQACEE
gYbh3JoPno9GKSa5QX2ucT4QmxtUtPJCNIdInw+ULishmDO7hVf6KqSrwcEgxae3
bvnVMefdLRSoKAc/65XTo6dQvZG+kWs9UG4O+UDp7SIG+Sk+JAeYCRdHkLwaU5b6
5n8YOJF0RX216fdVjBApFbmXTY3/iMEEpMErPFw0uslBV18RWSEbKt9R+L+SsCkx
aH8s/G3VudBM4yuYUuvRCIvp5H2MrQLw9S9Y4ZfUYtRenv+WYVcvyfkbHEcPA9ke
s2cOTj6GyzdbsjVDvzg4UvCWSC6b1eZkVuwuAmDzlCuCvTMJVEnV0+0k/vmeal9V
CVRBT9y6HYVhbTWTrWeHa5IfKnBF0VOyS/RlmaLQN1NT2FPlt9dm2XHUDpILeMt2
BuGfZFGDGSxc/JC3jgfDRnpGonovHk+m0vJgcVa04Clsf1KBOX7qIQkLCdpFvBgx
14hX8b7oQj/KqDPcN0HwqOUNiusDVdLdngLJgZNMWDJqo2oskXIzCgNARIatDEOP
CoIqZzNhz5/ZoCS9e+JwXxOO1LNvirHCsDtZqLL/pGyhX84J+K4CAb5pZ//ZFZ2v
L5AONjvUzyEDXNaA+zTIsXN0/sDdwlfWRJEUPKLWrs0XssRJfzJT8dWWKsxJypru
g8u04Bii91f9ZoDU3nGqzFZ6zpnERw3XBo+ZEFyO9N7WnJxry2znOpVWvm9f8d4A
9h8BTpOfRJTkKVaXQtuhmLmvlsfTFeGNOaNEs6yhSiEg+s+YhPDprS3sxHpSG9sp
9paomZ/KTvPREVxYJA/wxhyO9qfJVwReDpPnxsffhk0H2xtpp6S6n0g2nvEdxe9Z
Zeti/CLiuZhF3oMhRyc2gw==
`pragma protect end_protected
