// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fqBzuEqknwFJsnvJOanFvwxQcXFuiumIwpusnuNzSRpMSL6cZG40OfmOi98o7VO4
dEWdaXC0h08z6+HAeZuW6k6Xz+rnT5i8qYBD2jZslltCkYPltxkgUZczqbT5/bF+
jc6SDnloa5w7nV41zIA6LcWCKB3gfFP9uZrfbx/NvaI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58768)
NLI9c9cakd1c9BpZ3FnuyYGUj1iUpEp9AZNqfGkrJvUhSN8V86WAr0VmZO9xvvg+
S4PQTOMTxB8J+z1IXmj38wPTPWQveHxhHOeNRZxwkEU2Day3Ciz4uyoFGVGE2pZK
kLpbtR4ros3yP2Xe1/kOUo3xhIVEZ4W0oIKQ15gsSzalhD7GWfUzIvzE1lI74qFD
AfhF9utexQk/65NLnF+96OxCZtVhUgjWkzpgcHWuBdWUbpqevc0WQFziAYiwqOI5
7dfRoiKADjAcRNcBp0zt6CH4ntnYgiqNxJwurCsgts7GboSFYVeWPmI9brKe9QMb
fl86K3VVM0vcrUuZ1BsDZsvbXCRi7T9RCzkZ7O4ek/Go1VL1eRCuYUxUSAjk0eGF
rVPTLV7qYKiqfzFN3DBReHooz8lYlW43/yb9Fp+6NjCOPiKPvNDz+duA0U5mXB6g
RVCq0AdWB/noSofSExKpywK537Rd3y+t7mylUDzpbysxPXiHXtLm2LJrFAWpkFmm
cBgf1JwXNiy/x1jLvvTM/3hj9z+kCKTz76/dbo6W4VIx/pMsfqSm0lfH7hXLkfFl
1Y6/u1P/EfepUbzrgBHb6MXDBD73FlNkqvaKoZJBIjXqC7UFgiQPbyPIB6ZJEqBp
DosQkdfAXS4EdPYK/37BtZ2tbsSLvnZG+e/Mgz/aUqUSxt+Gt8UAt7itLBpAc2Yc
TliTL6wStvRh+NTObKqmOTS8s2VQGaDrGU0i422Gw4Z7ZYyMry5QnA3LZtsxtMap
GSiVprQQNWVtbkJ84SlHoBf987Pke47ZCw533SpOExdwvCzMvfwDPHAKrYl6jLyw
3usApGeoEnzCkWmutSURHDAOdxFbMfuWvPia8zqrjKgHQU04uK5E3sr72hstRj14
k80+InVHFczAAqJLvd+LvUsDKQTP/LB0E/jA3lyxp/4NRJ0zsJ2T+Bvg2JcJygDM
wvshJtaTH9yeOgJIBQXPRW2277AKw1eC3UvxBSIQ9R8EEo/2AQGBZctEIKuzguLL
sTaLf01YbKNOpwuoQ8R2bBmo7K/GHXemQTTftcZ755bXsdZMTsIL0qRLM1Xfefm5
yTP1ieHsdv/zNQUjBJXDnJZUzDaz6R6z2pgT37tWury910NA7hkAMCLd1u7dzPnY
ibB0MEETvDHZC3gRqvkBUj07WYuCrWAilqwsex1uwP6PZzltUXC+5DTR3JgClX+7
KDny1jJbwt3DBNNW92p5Ki8+rZ46Rvh5fg1+VrxljYgXV22kvn2e1CPUdo7zOLrR
/sKRsP8vuRsdsLpbzv/5It2XVEX03FT9fJW8YzI9WQSzla7sYVq8ZcMo/zz50MDf
APaXModRkKxYsMrl1SsE2rhXaQO/wMPdlDwiTBT6sWJEjnBpHnbcK7AJ8hzPnEcz
h3YJgd+czp+HJYzeoHdoG10sNidHP6tbZ2Fyg2kCC8D/e2f/3QjzZDjk3eRBxN2y
rWMyH4l9EHDjEuCkCsMltqj42NrMT7xfeBxf03mB5g+AV6e6oE3ywmbes38EIARl
QB7rUVNPzD6jWAbQc7rRTfWHRhTLIBuP85ipkr7PHLZbpsHNzdQQH/BClOYBy3sa
Z7+o3CVIkYohmU1uDUvhwr9k2NAXe8cpyVNB0fwFXbFlqAYIUcHT0RXZGvvqvT3o
iQljzNewi1Zy2qKV0lWCnDCVlsT85seSpSICMuLjErWNG5vimaxb9OGtpjw8gDBj
bVE0R87RDIGaKQ2IrzqXq99h8oCrqXDgo+mB/gJkywAkqwF3i4tE6xwVc+WIk78Y
KYoYLcYF5gGVV4dK3zbRtuwV2pPYpnkJxYBJk5fXSZZ8EWE+ytjKprz3hMfnqWr7
36Yv0Zj7oQUBjIaiH0pv/7CZPu7/ShMBpVe4F80CN9aiA1NtBl85/AR8FaqHTMRU
H/WlcjO6kVt/KZrDJutMQzbjjFnSwAP8+Yty5LDnYUe4PmXqFA5hapiOMqaNXDQd
g2TCjY0J8Do11SI87aGPecw3g7zRqKNZSs/ZIhvHaXKxMYgcT/AcS1PkvEx34v6L
JQjL3ekmzS/57A8y5k4hn0ctyEy1AIvyAEztGwZafCEsF1bSW0JjG2SoZD6CK6Ur
P9SO7MoiAIcvq9VQC5RwF+sv2l7Sbrftx72OggKuNF/hRM3RaSeGa4kWxTjbEVDh
dZtb2ZEAOfmHc9WZIyIU0cuAoBfQRJJxVmUa3vDCcBWYTiz2Hwt2rIVJSu1GzBUE
BEq0E4chxsCP9FkrJLx5/blw7UIpGgwoD42j/1+mPj/nOnNFrtIxoOYRV9e5SZ1x
Ce/ol+kVtPx1LvUEC1oeXS6KmXbN1fjJlwfB65hmGAXtiTCqDYYz8X6pKxi/fO5G
vz4WZqi5mgfxMUIIVRut5AaqrMg2RbZv+eIgUvAW8bwK+8LIYBIdMvPrUDVHR8yL
qpi61/V/f5aRyiZdQrAOhD8YuLIU0ynDLsGpVblJsfgXuH46gTpFCc6vDvYZpg7q
2HtamEt9uPieDoI0sCHG/3808rash6tEOc5JkZKlapp5TS2832bjw9coEeQpzU+l
XBhkU6QjeZ0hqc4lyWTux+FPK+LaneMkidVreHWNGRjHoMArS/exs7jvTPQXoR3j
eGAxvnSSeiNKU0ois2Zoyyf6KQTxG/QEcxsEsx9qvwUpKBMQM+ebDXuPGelBCT1f
1B8ITuB3sZ/bwiGbef1H8Vh9DlTkNMvajMp6SCDVm7TpnxJPaDdki6V0jTzKu4Eu
XT/gS3L9XCKT9pUpTvcfi1W1c3X872ijTYMKyWrEoqD9QiJavwlzgXpB717weClY
GtoCClTk3bGJe/svscCpslh8wrJRp6pa0NoUxdDdT6aR2LTZPlsEyiw70BOwKvhg
2bGl3TPC87dwsRCr2J3Vwi4CapzxTbbWFp0JxTVDeEMA9LREm2vVINLEQ4DrF4+8
vy22w248Ocf18ynyeVYKWOfwugxMRclQh9zGEGNp5k27NaEMmFik9iq4l7M3a6Nh
0F95w+lwztTYs/fcU8r8z10JRUUg7pyAF8vAE6YKQu8+cMXwwbNPjDivYJkxUp9d
haQ+PVBRaQaWH9QYg1s9yK9PzArno25f4+VriATaKpRdwXZHGh9Soao4btYPfx3f
6H8wXdA8YBFvdhXDTR0lYriuuEEZtoV9ub5U8i+j+Cbrt359egOYtWF7S8NW9THd
AXo0w8bt01rxz+HpBAUDbOJRo7+MlanVEm4smTcl23lv2+SzRxfFucK7YBUAi/kr
ANF45oJnf35vnPTflfA1PM+/wTaaaVz8brM4lpAk7KnVvjO3/LbZ1m7mROyJ3ldM
ybP3lhBCAHX3cyFge4N1jZ2eaTGT6SqSG1vGvkHl9ZnrOXXk9VPpGxpf2BnFrYs7
4GFqur2TL1h/UmL9p0YiqsCNwM19eV/ATjOrjXs2onfcSDhDJk4ijqzAJ1aVCSqD
Ij09mSVbbfgS2M7632B3D6aXVkIJnXEIvFKi/GNfNcqqVruSuohcHgvy56vTKPxQ
X1c/HPr0kwQel0DrtKy/OCdOPCfGx6pNs30TfxjjWOii+y1h238QLC3QNpPcB7PJ
YpHb/4SrGhpfk9jSYoDiN7g9rW5PsMrJ+DnoDY+2AgJvpjoOTj54u5FWXAPWIB8l
mY4OnJtTkY9x4S4R5SYCfVc6uTdYN44ngSEXuvTAuPHxmMx3Ks0Qtg++v5u5le9D
+3Fqu0fsOm8ZFCe8MMrrxooDLhyaZTm7GTpl2BibpYoWs1JCxYGT6bSjzwt+Q5UE
v7St4liHTssc018mo485vTGvuwbLsKprnADDDxjS1wsVxFHOA0wsXU+sx5zeQsPk
ek+99L9iozz6qbpDpkYHlQDzZM7kLcYAjrzEfnUG8kmwQOY7x3GgM4UalwL7UR4f
gQpAFLG/4o/dO01QWtydmDQoSwSBmmXW6yiTGJ7WB3aYUU494iX/XYqTaj75hero
XhCsYetoCSIvkKyqLhM0dXuXcfcoG+wNddyU+d0bQqGeeaLwAqdhaU3d1UT69j9h
Yw90cJoevWXGZTbvZIDeX6PYACfmpWWfoPWLYcL33zN4r/eAEJX6Ub5NMD9PhnPC
WAd4XfAywc6Z3c9A2p07/aYvI+Wj/FMts6nWWQBpSdkBCpIpAAojoFBtP8cwSgZJ
oQjlWZFZvh+523kh5GC4aAyQSalWIOvVXH7WF63qZ5efTrSlhFos4mr274AsBVzT
mN1w0sVz6WOnOplbfTurqkZcLpTkPF6DAuKAYx9N1sVgLlk43RbvnmWwdbF3Otcl
6U9wK12KOhzGR1Zq2bv7xCR+Zj94WK2QEbS44RJ6h0fjj9Insi96a4xPC+XcZINR
5ZgibnvuRG+DNSnZ/3sPErh3Nbuoif+KiBQ0jvbFB9OlWrExic9te/wY+Sy4yZXK
YS2TC1mf0qwHlxQd/E2KkdNKbht6SckZs7QTyP1mw0K59oBJa+itDdrc4JLISpXO
ogWBlXIAlbLfIZG6ymlqYqosgAWt1/tSE2di5F3NvYli9A+zi1c53dOKwVp4gYzF
DaPOuslMp/Jggo4kS6pCRrjZOesJDp4Pa2W31F18Xiv3Cbt8kuy7RRY7OlT6DXbN
D4JQB4xuQ8Uc94m0QcsEUAITG37xAHUA/5JVLFkU3kJEPaqSW+Lwbf0p23UJLxaB
udgm0ju6sxkrJJa3AnM9z3h8Cor5JS9n5lA4wB8OzDlP7mLsoYBIFumJlS60gFV1
Zzcz7fKU9kuM6TBXO/901vOAMQwuDyGBNQr11SQ/8OXSvcCfggdGJUxivr99ofUi
jEdB62FC4ubPo9KdWW5jWn3sUo6Ob6ZUoD6OY9lNFysZ79dxYNAVOyGu7x/iyFDH
+uW/NVpPt8zeqtKIYg/FXLFsUPav5Q70mtsWEoIizygB7D9gLw+aXhXeH3FTPVhn
4cCRCiNEqFLUgE+NqcwxDpwoxR9lm6HvzKph5CVU1UCHyGrEYp0ghjpjNnxsLnWE
Yu5qSC9SBVemAuz50IlCCJIbZal8K58sHjOxIkfASDKkHCtfsRGAwfKfFNSy3KWB
ICVqVN1t1m3kJ8atmQ03UJYOCmcQETI8mtp8WPWW1qTgY+stl01gt/kCmE5NORLB
cXiRbtaEfxcI/xfjJCnXEl4dodBngvj7wnMmsJPRdqv2vg7vODuvvLrKI52Cs9ae
Xxk6eAIY/RDjJTRg8RQSZRyKL5myxNu8wLIGRWedQqEdu66TaGe4ydxZdDhmmK3t
Q/CWSX6CNrQBr6+lUNcjeqSmDfQjKXLUd1CZNjNdbkX4UhjiQs1pHS/kR93syBYi
RduZnAa/2JzaTzAKEvOgplep5+uqO6+Xfec2ylMiYWEyxIwrwJfFBexoPvJATyvt
mcGo/DSJq3ZEdXpuUoytULxKvQpbVT6+u0bzCPTFFDqLIo0lGJTfqjfrNjhsFK3F
lY3AvhuHWEcRGzq+JVvEqckyyOPoh5qpc9RjSx95zlEVxIhOosMW9G+wlWPmq+iL
0gOkf645ei8R3oLaw6UXbTcMbBk+D8hDeL9+OCW6AtXci5u1H5dOr4Yu/Jn+Pc/u
kBXLQ4sJWulhNeKBzqzEt3TsDjTrCBqkzyC0dKeQ9W3vn1t5FAA8tAhl1M3xd1aG
a+Yw2myLlH8Sl5thMaE38AfxscwrYD83IeWJfhtHMTmC066Shpu7EmzFPYyTFYT/
q7Nlo94tu0kbjk2D2pLqAojwjqqgxe/xFlztXVtH/irK07lEzJICOdNeJhvDpoTA
HdoUmkjtCxuEy1vATHwJRTe7wTB3u1mmb4voEQMZ2XlzbIWQ/1wyOdYCLh7v4MyV
nGplccOYgJwuQCEGRAbxxaoiOmFLmHauE3n0N+RakncPSv93/6Va/vbqkLHR/bAC
4sN0WN0/r0OImz2/YkMq5dxhKwNScK4pk116buWzvYYcMhlCSfVUo2o8kMVOvmuJ
YvDahCb6D/ypDiZ2exjKeH61A5ATJ03uTqupKB7Y64iZQMYifnEtJsALbYzabmic
f2G32Gh+EC2Ki6zwrhRq6nSEN7O3EOw+LrJDwV8jNhmFaSTnKIBuWuZtP6sygy3u
2SaC+T2UD7MXvB5CAN+/R4K2AtxHgtF4RyqUbb9XeRND8LS4+G1W6GZngnc4FzIU
5qI5gwgrqOgXGkQx2lGmAxJnHTqQfsnW+jndMCssSYQ8vYZbe1Ck1jsO+7nsSuTw
ZFCLiT1lb/FakJmAucccZGTvvNlLplm43xglRyHTaZdyr5OJm0oA0R7c9iZdb1oD
FoCUCIWcO5Q1uNxgX6mLkNQRaDRCbR6COLjTTWaiS/t7Sy+St93pelPt7v/GSymD
dM9t1U4lalMfZZwBjDP9nIO8Mis+BBvZBUlyQkklarAfWlAHp1rXPyJ+g3j51Nak
EdWwgfXE10bne+nzJ8tGVZ0lEyWxm44frd3Ht+Zgp2wZRLIpVnl8pYH7Y1vqO3Yw
/LG/CuWjicdZ1zNa9HG2/Am8Aqy9nmYyHst4dDRuy5myy9BtLQQYylhM2koznsVD
+9oC8vTD7sP1Mkxg/MTluz9vt2OBPko+GS+JKhp0L90FA5ZL99XuwYUqud7mi+O1
rWB5AeUW7l2yZeCdMjCkQ7l/YjysUGUfOgghQH9eVcwOL1KNUk+P84oDlR5rsCzO
W7xYrvk/1zDd9EoRld3p8Kr/u9gKU10sWDR9Bp5tmXaUo9E40AvPCEjW36yxRgRA
ZZ/J+mYUZthtbaLJS12/31YAjn2BhjUbE3nZqjy9wM5hQGcCgCYaQJAauLk4kGOO
JfJhQ4Dya/pTG6OOoZvUetCuscaEl2WP8iakiBBUjeBWjxz8FgTrKwASfZ+6I70o
5k2bazqb5NV9bhRNqQFprF5SGj8lH+LGNTUY+HN7SujCCrDaru6Exg2byuLC7vk2
JjOgyuYzHEUSj9n4324VUSiLsm9roBZV/sQmDEMTAD7c3C0MkSKaWKqOdSlKj/kU
mmDWsMhtWCP4XZ+YeuuoiWw0BxdkmFHKjP4cgm8Kok1L4L7kcZuYVmX5z6SGiTT+
+HCePT5bDm67FFr+kUV2X1XVw2kK7iOIfMal5ewDpSmLeDd9OA2z53MRYe5nU5mz
TQoe173ufKvLQrU6Ty4n2mN02NDhYFqdfSVD7IAgbBAAPVqVBnKaymzMC3hXmjLZ
Pjkh6/rVJaxe976pdDrcZTAfmQOGZZtpgDpbQXAmASnvZ/qPmEyYQ9qViQN4Q7xd
TUF7MPjH/a6xqdpuJWfGaF0w+0YuV1Q+9xRgyFgBl+4BTD8kPPSrBaPXLYQeeyzN
r3d2WPLKqNf1tlyq4rHtCy2YfFmPMoN3SlT+/P2EyzuYaMK2QTen3iC2Sy66WJnp
gbqlywWz3bRYVSL1JHZbSBxQcEzL13Y7q1y+1zZvVfE84wVALWV059y7UGXdoG8S
wCFlrOu+cGfVz0C99z+UNoW8aJB3VG4utyApuYGPONODedHfoOIf5WXswQ6aGDGv
oxWO/k0kqyrPTTYcPvfSB0oLDll50QyIzvxC25xNX0HuSz5UEZ1wwWsJkpvJNrlv
PG6DxIdsXEnE25Fs5Jve0KRSZ05Pil+yIt8FGX+0qXqmj2e8RuANpVVR79fXqU+M
0zf87X0OE7mUnHKVvTPv8juimKWx3CdsEp5g4xPMMeWTM1/Qhu3C/gQvBwz4Tk+7
kmGJVlEFOKEo9R+IPlcKGz/jK5RXHEssHzbx4NOufmdoF3rWelV7y2m9bHOL7Hlr
z66iyvow0HQqqZWJCJ0Pfe1ke1vctNxv3EwymrRCHD9xpbiFcCdXvAJkUfO19sfY
0mFQ80uDFEGmfl+q1cyYCPlYUci6Vzevx+Wvj+Jzg+/96LBNsbIr0QSkdmrkxUBQ
z+eg7tdSf6p0AVz5T/Ya9tupuhAJHEe7gBT4gDL8O1QL98BVmVc0LIgS2RA2XJGg
HtFYxXcl4i3H1F/qqdw/ID4p5IoOZxZByEYswlemr0OB48cEOrfWbqHrENS2IJf+
dpouf3ZvyjdQmfRVJKYtr4h7HYQIn78aj+Noe4A7f+rn3iFyg5xtGyN/deqBxvU6
7JE9mB7tZS6FmBD2mLLGXeFvietlBUyaZW9wNwtxG2zwr5pvib84UXtDL/QNtM16
qI9pmIyz3nm3xaRhr5DJDlNK4LcVHYEyLuwtMWB3E74+on8wdiB1KEe6CzmnvM8e
9GmhZDjI6kHIIQpp25EC9obzRZE/wEWmN1Udey2N2v9RU4dkaRVOBDkuTkpDNvNG
9lzz2TaO8HSjt38e4hj4gB/Z95FyfG73Oa/vakZkUiTXGzIDdHJejudvX1VjYGrG
rWi7i6s930XQ2xeHILU9Ollg+SN24ZWJeVktJKngRxoQOIOHMephjq/Uk5T3Y2ue
p+gmsK1GowkzDZVf3NZjynI5PPcy8o2Yr9Ep1z794AzBeKsIzgLT3Kv7DY2LQFtw
fbhYwKvWLNGNfZyFUjckrlXBFg6IInszgqYsmN0tkHaAW5rggVwvdtFNJvVxtgex
naB4w+i4UFqGij+HpvGXzpGSzPxr4vpTsEzBP/xgpQMBTkZAYtrPZrxt3faKqnNa
iJh8wAxti0NhDVXXWZXogBbgCjF/omVbgHuvolTSHgj+/4syKWmFeEFtkxQuY4i2
w6/XLMEum3saqogTFEU6VoqdykdYo2amxNu8nX0b4CaSlUXugwak0cJxYsVA0nNi
wxpzqJOj3kQa2cnU6C/BjZRBuJJtdr6MV3xtm0jrzL6ulraVCAX0E1q/2R1EKUVh
li4w5aqZMfjGDVQHf4xFd6IBluJrH6Dzf4AZioRHdrqbZFNQQZsT+N28ge93FzRH
L4jiw3AQZraTd6XZTnYvkvQByvExv9ij0AUVdOdli0febArG80kHT8K2m6CYyqi8
z9dt+Qc7nHNJ7/YhSpr6Ccw7MEd6toGZnJqiC6+B0WMi0Iq8zqVPGXSFUwYYqRZ3
eDDhH/TtLTjruo8Q8b0n1F/SF9b3EvZ1hkQ8KdB6HTgc5pFcKh4sILqSKwja/isy
zh8UcCYyta4isPoJ8UV6K5/dXRa0FAG5s9qCERRUXRff/Enehfp+tEOhEebjkVyN
72RBp4tm4TB4AF3VuHkzWhb83DgalH+QDOGNPXuZxtDM7YphhQu9N/HKx2ce/H5h
4qBPscy5IoM+of3YPZSrU7G3PyMw3YVl2Hx8Gmmx8IlaqAJgpDc6MnWiGDESDhiA
FdZamqceWrEwRaL+ZmtUNllU+lRKguWa8vcF2migFFsElO5xnlaWeSfMXY1Nm/Mh
LS4BwLUrYgh1+9Gg/I4f0tFztTUUiFICnq4DIv1Kx4W5s/5sMikEonGk9BzdqT10
GnHprr2XZC2Kc8gSihvbz53EoOUa8RFzW+g0Nvew+M+v+GuXrvVRRpifcV3uh78X
LahiGJ6AFmbbvAgGY39OQX+2McnCoN4qf9/hcNHE+Kp3Jip9y0c3OMo9uaYoypG+
R8Efuq6vkw3njpgtk345INxIRNH2IxdOyOrAeeJA4WsQ6ly5j35aYa/gnaeyWaRr
YBd3pl0FgFmQmnaNzq5va3Vbd+S/VR5ItyGd/FIqtd6XwUTM1TzXQDYSbDl/Na0p
OAhu24H9xRxKo81d9mSbNdvIi6HJflxgXTnM45C+uVJx2oD9P7Io04exDBd2GdM2
XZGH0ahGROK5TbjtGVSzgMAsKiB8OX2OHlv+hoh+S0lJ3gHkSIlq4dRBuTPXB02w
30BoIVUze9a3HTACnNGWoRpZ1THCGCm1PexmO+ybFLPGrvuLElO9dwOG9scc2Hle
aGPLF81w/6NtKHqhwJsNA/6qhabp8/U/lvv7eqLd2ns+GD/S2SGIkxfY0I86tawz
g1W4oQjhvnKIEzKzcZw06VtFmJAI0mG5wXpOfPaaBMK7ck97G/KGOsDpQFfaLtZ4
c80X8IGmkSHUb7t6a5mXTdx5NxKdZcTqkJA925X1mUvV/L0w9FCKaaAp7GddESUJ
n1LLigvrUFx41RKh9AiIaRF0BC/Qu+RTZ9vIB3PC3ONa6KBRl2wVhIQpPrPNpSmg
8k4X+3o17ncC5y4V4hHP/+QqVl0SVXrg+9hcI6cjhH+HaybmHNH/ljjVj5c/wpa+
bWgTQ2tZZvjR3+29c8cgkW0EiITJ5UpcewkP6q/NskCtLvWT4GylJZM9n0bEuc1Y
EhYGLXUUwh+2tjHznf3Hg1Lj49m1uVIcd8HwqMqMIXONug98rBWZIQB9nV8zwRYj
EAX95gebWEpjqDP4ZuXc9fNTnlxfESfKvvxQb9ljntU13OluJBwyBUnhffwemGRC
83WmmZC2++kEOPEKrvKbL3SxHj0bQgoMwkg/lCXjRoTRZ9HRANb75vorpuXP6B+K
eP9RqTpz43jseUWaXz2Fs4QVNtLIo+zydisNtrCj+tD12CygGAUmGrMwxrMWNgVh
Symd+kON45U0x5ZBGgJjZRs0m+5UrqUuL6csO8UIfP1ceMWzZ93lqxqsj3kcNjbM
NGhQEoNxML22e9JcJygjls+DS6F2K9x0HYgzSpbs5B5KgK/EEFbIOiCdmMzow99a
CHLbcW955C1ziWwSpU2Ami2AuhX/oPyD+B7ToX+WVyaIoumqHzA+JmAjifiPHdIr
X6/MJo9/xrnKqjlajiG5M+uXjQUsHx1x5oXzQLMQu9E/InkSerqKTnJCOR7RsOdK
m6NnEwKCwHaYPNnOA7U9a9PWqkcvKMbgtGqq3KBfX6CnOmxVeQyyHVARCBK/Z8sZ
zb8tozyQ33w+CEkZkLSonYOsz7Nmad/nMUbRJXSEi9lPYA1xfvPf1ldBxztAUdvX
oZJ3YrsI9gjxIqpd715RvO6TNY20B0piSGJ1tVzU9V/wcBeDi8HBiIMwhOy3gQKD
tS4p2/E6qIGB6IxqGN9ygxYlI8IU0PioyFRE8StRNqxkGxs2azccFqq9V33IgNJS
+oApZL1ApR//QSQF5b35tJ8eDlz5hXlvDHcFh5fdyKMxgzG9w5IIW3WLN1hvNqUC
T2rHp9F1yxKmj6gc1ZOd0zwxtfjVqCkmmmvQvZVIBDzQ6LaZ0y7EXMXI3OS0vAQD
VGFXeJ0BPHBGBFVQHbX73QSV7E5kEokjIh7S/DyvQ6VyLBdHdCaiylxk87ZOZa3K
1eRRwtXrNOz06BjqimdEjesfxZt7Ukk/y+KTITlMlsrvdu1SY20NvwCVg84qrZlG
JrjGVg8AM3TR2mY0prZ+fjzxi9H3tvWmlz/oTw9U4/quKTjyMaBrkbEeWNarCsU6
NAWlGE98/fLhscosiwgwUJBPXQoTVAenhIDegf5emLYLZLOnebkg8WZE4iY0NVr8
8vmnVoIYls5SDVqU2Dif8lYYBO50fe2xG9PkFnfrhqr8eiBToUpH7J344s7m+DMm
5SaaO3AcjPQLkRG3xUqL7QLcQUuC+HBRIW5H6KooMWOJluZLTIeSnpoG7wk9DXHg
6yRnM2HRiX+kya5T5RjC/gvkKZvpaDCA7/6jnvT0cgjhE6B/bNavUFdd/tS8YaCT
0F6Tg5LUmClighyicoYpFVsxxp6GYVVa/CH4HFZUcSdlQf2uqP2TY10apk7OjBFj
ZHEvKx0Rhuet1S/jjR7oMHzQ+W2lR4u5eXx3xCn7LOKFkCoBL97CrnRfZx90oGhS
v64uYTP3dnqTbpkG5+ADM3DxPIEa2OzqlbGjLegQ4dkVgUtoie1ugOute69WW/dm
dHKMNLBO4iDpolE7F+1z1yRVN0/Ygx6e2eyb/vIsWHdlzlB4/USDfa1oaxgQoDqV
yYNKyfp5NmjJU2TMpwRqAlwFTAKBecCHxGrAWlINN/Z/DUts2HFKavMj5GO8YpFq
HW5DUrkVfCOjkXn+63wxyUI+hNLe/asxPGCKH3nesqBwuuY4be9REnLeetOdxGGm
GxzgCFFe4wGX7a7+cHB/psYiBF2tJp338trKEQxUhPyU6/DzN6KmfLy5Me2086fM
gbuu5ysGs3hwx0HwS612bbUEMJHhoAtmFNf9zlJi7u1xVPwjG2CCtEE2GWMSQbdC
ywpAb4vzF0YX+58CDLQ4m5BtgGLk6+Flj+/lYnfLTlZKhxwNL+kPRBTjp9syjl2h
coDw0TDCQ1a/FTMVIxN2/BLkyFnW0x0vpm2zTyKK/6CJ4+5TlBQxa8oEl32dmSSn
GgiyZx9f9kL6iU9gjDH6JoiwHiQqdfuBClmXQ6X3NmBypbqJ/9PqZQUDSa1RPWf+
Il9VeazwLYjCHmTifPi2YE+q3fgLKMZLPggutLP27i3TMBfWh+oKa3MHLIUq7pB4
4zR4Yq3vTJteDYDm9JkQ/8CAMIvciRpieXYIOjnYWKAoD3ZJTi2eoeXO1dK5C3oC
j+WvqEImKrRYSlsOjfMqxulDfp11Sxa+7mSdTI0lSfLS89kos3Rd1SBOBGDq6iOD
gAw1/gLsVwmD+APMS0BeDi14XFpgHcn9gIZ6m4I12ylv2d/LtEIaFAMkLVpHYsSa
TrYOnyvsA6nchwdh5y84G5fsJywg/XwiUintqyIMtoQc7t3sETjdHUj0MFKBhfoK
dwAUxiERzthKxz4atmVmegbRy9WammnopzpGU/o9bQx+4wL0UAPG0I4G4omur2xY
IvgFmFEusW0zjsBdIxRFvxENduT4sxuuklzcL8rumqtnqj4wqOA+d35ec9IcOj6d
V8NuvyC2BtyA0NGBXi6KTqYRDyqg2bvXGHvbAqb7k3M8JH3nd/scOD/AJI3vAN64
XOQmOEKtPhRbJPrI6yRi/jXzDO4jDK0gyVyQQFNE+Bc5toZSonWLaaQj07cPODFb
IaFEJzdTud1WFznZhd15vw6NZ3kxiEAhnes58TenHLucMLhjq3Yk/PpL++zzystj
Xhac8PM5r9u7Sl7n8yxLPEVhlVTpMzmfAaCdPlmwdWP4Nyf4YKFLQtRkueuktOcO
VxUEL8be9tEhf1fD56MEDHcFXYef/hD7IfHjeDpTDUrUa4P709VmlkbhW80qRyw5
NfSB8mF3UmBnpqtOHhIJgV+w8EXfYXv6QwLFZgHhS1IOVRS9VzhSp4V8MlulOX7G
lDavljLgTy35lLQ14feWQ57ivVt0jvLras9OQi8qWySyV94p+p9uEdXPCHgtzU7g
u5Qa2JqZsRdgHuJStNMYat/W8UwQ462uq61CDJfpyjetrONEKn4g8o9uJuWvmoDW
Hj+v86iKTUgiRKdRqZLRLNuzRBoHd43dfUbDwcWxVrY8WzjlyOYIfOmJFfi78/d/
ksMZwcsPTVmk5DywErRfrcIWFahsSaQnx8tpJYi8vx3dwcIFKK1ohtOMC4n/JBH6
kYu6wl9pLAk9fmB/u99meOOkIJaSemsukLX2ZWW/aqsa5WSvtiDTASKVLNq4PLua
aeoN4UBf/RDjv6DEykNtY/YNz5U2gRxrW/pRTEkAxJ9ecHf44YCAB+mHroiPU6WP
wZreJD/7rANsvBjsseigPt/K7yiCVW68waTvCJq1S5IXRi42m6zrTkZGIJROgFbX
yVMoDEGqyWMfZ/1lXUZTCtXVtInYpigi33kjDsUmJWuW7Dq8V4e2mshqreW7n9yM
/Km5jqE54+wHgP/JURZxExthzYxdilS+naBIwibt0QZAXI+s4TxDaUAID7x1LG/u
1RCc39F5fuKgCX24OPV3zRbTAV3q5/D7Kdh9P3BhS+2d2X7ltlvxrWaHIWPt9HN0
JEfEi3rc0PKm0cfPAyrcZfwANZ5Zys5tMUrYRI7SeJFvAGzxJJnPw7G1iSaey9dv
OiwEvdJPGdMa42aqhtR/Ee8oxbhGfMOq4JY9B47VrC66lpWQznsMPBNFQ5oDUOaW
CfXFEDfH/qLoQTTM5wNXifv1SHgwphHprK5KojjXou2IDMJ8STvy70pLh/5+C8H/
Xch+fHaoaPdcmSSMcWFDIhb+8AnWaYmzrDDGL8hTCPE9A0tM5iWcxTpB6DYNxfNd
O10e7PtIePbzc075Zq07xPtZtmO92bjF+E1t3E8hcXxLSDrFlcVsQBcLuzzeTYzS
JghZ3VJ9Ldf8i8AvI5b8bJBcRtJ6Y/8sqJH8lB4QqWGBxM5V65FxwLpQno0wOpBT
SbFjtT2HXq9r7w3+K4s6aUftd+1mWQcMeCS9BM7VHl8ppCbOw0EKrUj+JwGc+svP
vQ8xwAGU5Prvpv9ym24m+3uw4ABqTwfL4qJO347GqwFSuVJ+p19maRiTSroXirh4
B7yr7nuOiBERqMO6Df8TvnPFdjvsOzHYO6APp8PKlFNzoHTLKdwd+MgBjqiaexo4
uK96loR5uCopqsn2bWII/a2E2us0PwK7oPEXsSQ9eHBo9AVlj73qyA5rAxoVdps1
04XNp9814WjZpfkjlRau2JQ1cwdsDnwRMRbxjaEJSew9AVeUGOBvZzDK50yryhxN
m5Xz1aOAC120o/iwn0/QY+dY12ISEGTr7cey8nbFTT2ASsevhQaGDGjEFttcUPb+
7oaT86t5Aft/f0bHCF7QbTanuKd2HeAaquKNc8GylDOzzi5CcRWAwJiGgtle1KkQ
xjj/a49vemsO1h31MDccgLwJ9+dhZmaOtu53kGiWuSXjUIiyFeF/iKYGY9nytDlR
2HKHlSxlnhU0XUIVVK6a6oIcB3eNPCiuD17VUgRST+BrnWBFOK6I5KwaKcU4qIdu
KcJKgPC1pJlo7+UD/FypVL3C9Gza0DoyDK6bGLyzfv5bSuDYg29/ychv/s3cOYqh
I/uRjNseMwewD7rf5EKo7g88/7WfrRNu2t+yAq7ouFBMUvMGjVRZyeMsz74Z1U1h
Dj2eIZqYJhqFu9Ioez2NB1Z4QWkm0D1LLvQGAWoLexVPbzRcEaC7rKYknVwV1AmH
JtaLh/Y0oWqkhuU7zzO2CGyGAMttwG6cjhVKCkt0VlEzeZtdeCmVAeTrTKFz/Sec
TaDUK3Be8FOIeFMVNM0+YjlLZTldsQhvvA77UoNoViwtAoLKdOW4CQFUWZgf84d0
ifie7LRnX7WwvVWr38/GU+fm3QB1dnaCBXFCP5qCk/QkP66t0zZndijruAJboJtu
A/gpEiCxZCJZLgfPNl2BxqKAp+kvLU0FGr6Odk3rFbkpTqVpIkLy3WrSW5Xp+61/
h58SO0R3A7ywcxSIz/RmR7gyhVpQh7BYzfWXA8Jgxj20dJoQsKbOyMDA2vg6tGRx
3vp12gUpxcVB+ayMJNly+jse74n5a3KEQIZog44Q0sCGct5tGcmDFOw5Cl/3oE9m
qZ/njNKD4nV/uqDHdOlEm75WD/OprFxNcFTXpOJfLDrEkUz9t9PVRrbqkgAeUICd
rSq4SxP/mCVRavHu4NqP778l7nkvEfFrnAsNEcm/7BTKaue+3DNIk4gRvbp1Qt2j
Lbn42zjCyWkPoomBY3VdqbDJa2FqbnY6cTucYcLbwaC4Epji0/52zqks3pAKbwop
1svm0lcaoIXCNMBPngOFt7lpUvta4ESISA2NB+xyeZUz+HJzBEdFKe1FcWxxgLEU
5UWv7FbzF4wvK3EoxC6eQyJnqixOHMZfNY1E/PvIbz4osde3jUCtpYNx7FXf2iVg
Mmqw/eKF1GexHLiTz0qKF89iq/DluCnnUMp1aQCRTUdFspdH1ZIqwNqBMhc9upvy
bpZfTCO2Xi70+TjWLCDl9Zt6yrUNMfg6/EIM+vFmBbvJs0KdPo7AAzkSAzoRPGRQ
/rEMJ09FznvCqc29hVFL9O8LvyJilSAWQUVJdlP1kIphTggREZoi7upfuseSsv/f
ru8ayCMtCG5cVgXmgvafsUyZNlT+ogAQ2b2cZZSOjiIK0Ee0aW/9Cugl0BjJnjkS
1XA2PPZq4DEQQqMOnwk0s82CxYxm8M6/K0qddMMMBZBaokbKjKoFWfx6JZkfBdsK
/txuWs2rTf69Qpz2qw8TP5m0XfPbDivyLg4XFxFWVI/n3rQEolpDDlWAG2N3fcsE
/Nc+C5nVO3RERyhq+XVDBKUwlTPJGcjqaqhxPFQEihLryJ1w2GTHC7qQpUPdvfG8
hyFu75QUcUqkVx7P5y/0yBYdt3YJDlgZB2Hb4rf+dIaocJ3FvaDCtMeYPc4+UQEH
ce0eqoNA52Myl0PIVa7sSW+WvF7SlKQDxvkJH9Okvk6dWXTyWSUsaywluTgiuS1E
2pvgnrASVHxw+xLe7WaWGMDfMpsrtQUpr4Yb8SF11pmoYF/GQq5JMVlWLBKQNzlv
molxPGOYz/ewtfNohYrFKdGQ/ClhJysraMtVssekwrapdOZEDpMnJYoGha4SKYnT
q5mkfG4jxZXRlryGb9z6IuelX051C9Qozn/Ul0RqJkzGKDjopiStHNyF04iDDO+J
xSfTuJlohY6Cr9x6sG122JMPntpc7gMeflFYs43pGERek6IWZAb54aRLY1vq0ll3
jdiRvMCS0DMHFohBZwhKBGC38+iYAEmHIHWDAEOqKqQxOJuJO5tAjQWPD4x3W2bv
ox14DS2r6H84AZUSuv9gGNWEnvds49SvRdeuvOo12QPqn/W2coueHl8Ms6QoNhjp
VhCWA2XD8TivRef3PcGtnOyMzJYAHVM6mYmBsCZjvKO66ucEsUcbqq4rx826BzX3
3kncQrWQFHn4R047B/TKAvYybslQHjnVYYs2cZuNV5Of0HIv3nJtTo5wNC/BJetD
8y7PHXAznYBPzXR5dLMd6QQinCV8UxP/tBsL/D5b2cwVXIdyciEjHkPBTXheqVND
h1pTZJz1bD/l06poXEdaCLI/tzBwqDAkVySOy4/TgBI/uyTrGAzwhQwa3stWC84i
oM1ZeMBFfpSzXyrPQQF2qblVh3va6UUcinl3K2+9zuheB+ysE4Uzxo+ycslqeJul
aQGZdrFaWKP9lg1rKGeWMh0awEz3NGsECO21DirycP6zzl1SheHBdY+OINwgViM5
hmyCzHTAUtvkqsNPBnKokzJYgREptnPC+HTcWusIgDBx7r8hjwD3YA2FAfQYlf4p
903+aSZf7sPOzqprE4B5RCoIEidiyTvigLskwmUYp9oK4jFC6gA86WQevyERPYAw
YpLrNz8eCWHS5c5aApZ1NWnoQYf7nBJh6907eZk4sToKOowEOjpMgZEZDal6QI5Z
5WYx7ee5W7rFMuIwRWTPTeaH1we21FR0jOuFvpSydAdhkQ/VvJMxwiYP8xg7uzMd
e/Pfzoc3C40cMabguou+J6z3kEvFVKAEm/4OZhuMBrMbvWI4KQy+CXYDCg+xiIBi
skzA+iznywCx/rVyBt/TXiuM3RzucYKzLGVbbFUxxBMISjr78ZZfjh2hyruyzir+
lMrz5N8u3vl+ZXYdK5/V5ygGLw8jGTIbEe1IWjr9cEOJ6XL0sVbJwi1di8IRcBv9
uIeQ7AFJBPSoio9zH6gSv9KToRx1C6BQPZujur2Fh6u+WnVlgI4SgxrVnuiKfABK
vuGUIBw2q/AWAbYrxDqkMFRSpopc+OchKQGzcSizjigpZ+fnIoI4ylIM/kCxSzOw
ihLUvcIsM34+Ji3/tkVwXeTdPbwX5OwV1neTEmHDsj2D7xWNKF09JfYMEIhQSrOU
3878keQ/70RZwZlnKz0JAqCzQCZ5jDrdS92wYxZaR+uA4BpE3qBGUj4gmRyg4iYD
o01gHksjUYRq3Vrh9nTx54uUMrfFE5rvulDp0AWvZjtEnNL9EpqccMCFfHOnmf4D
bycPr2rU6aSe5y9yx4nlZ248PkryHLdIb2VojQwIjGP/nSyM5Pi3BF02Xgdjup2U
93z5Dusj0DIMdoVMhEb3AFgHucTQUei64jANurgmASvjtonmJDmYsPvhmeA3YAgf
0d+Kz9n4m4Bzn+QIBfI9G1i0DCoehqKCfhOcZdaPc74pol+C7c8jjJsQABirx7vM
f7NAvzYqUNWaSS7A7I9OztdpSNFqepxdI62TDP+foM2e0bzbW8acJ+U1oTNIB+r1
YJIpI8J5pFBQMcNSr+hBOw7dT3XcUGOb4sjxnQbDQYesv5JMnoM7k8ahNDMIDU0s
yfF6tDstOw+Cejr3kdHKTomHG4xnxSLfI96wkr4wAqhI8TZlQNe/WSQJj3Y2BO5U
Qvohf11pUU47BY47uls9p7CcaGSjEA0PeVYiCZbEd/UHBUQ+QiRcj7hecT8XfQsr
6jfpP1wKErla1y8TC1eNe0f+VGCHbVRNHC9E1N1yAvsbOxgsWoQ/E9gotcIa7rFv
SeeaZYdvl+Y9pCu/13ishCPu9gndGyhgAIlNtZhvXHQXRGXDTcpXeFgIJxWFW40E
0c5zACowHX7vt0yszJ5asnPg8N7TTIju7Nmpi8XwD3ihbo8Ve2Vj6DYVDMH0bAaU
FbXOTWLBlbDBIET6MzF7ZhrvFZAWzWxkBfUkoAOo9OcXZiBaCRHyppymwHMKsQpU
YlMaEhGxJsxsJXFBRS0AgELfyUW/mq+KZc4xWmfbyH3k+zNzk06Q862CnlQX9urv
jaxc7AFIqbRZGtfOvaNyQS0nKouflcNN8u1hjPrwMdaP+7EtTdT3B0hiD9Qs364d
WBV9hjzdJkrU1SCpwJN/Uz5BaPfEJazcnlni2GBd1CYFWxSDBHaK/w43JtqEMcdQ
7SfC2FOMaPbbKb8S5Mw50qY6bTHc61cRz9ULlaEHElxoFl7oTzjFnKAfoLmdqFGj
qbwJNFcYhthyXOUylYGeQD7DlMMPTfSO/bM3xw23xC9xOL1ExKxnv7DHE5y4qG94
OQ3s+mfl0IoorGQv6YBJQl0wBFNW/PQe3COOiWf2TQRwlteHJ1cBLlLzn6jcmktA
lxw8vWXFDlvGhLtC4UA1YRkP9JxPzExjj8F7HPUdyHLnGBEdCoAkVKyq7qYwYvIe
LCkAv/9urmeF9yCKiFY0xwjPzB7bKNdMBF8fsV+jSC9bKzcCVXnpt87t5hBG3PtV
FRgcBvZ9YSBds3bhZD09js/skWgXD2oQ53Wc1tM6u5phatUg4h1czVkPFkQXmRyp
L+zEf3P1KcvdDNa/xQ0fHI/DSjrxjJ7sTSW2FWGDQHgbXhJ2EgyAiPVyF+rAhLA5
Rifx5iIOlN2TU0FkvjChk++e+G6LdhVsL0wwZGdDQfbdwJ1MZfF4MAlDa4N+EGQk
P++X2dOR9vwbpVkFU9V21TsoNKhVz5LLgYaJe6D3DlGCD67NrgU8Vs45nQQqboI6
lOLbU5rR94T4jjPjws3b1EbaoCq8j0P8Uxsw2s9Ra7dyiaV6sgwlG2m4iflhBiNp
Ethz7VxyAU2LF4UGuqelP9hLjq9Avr+oXH6qZ5GVDphLIEcjfUGuAg3GIrQqMlr9
PvL9SALncEMCFIYmYfz8LfJ8HXPAe5bDxRXA64QtStjLmoGgUfmMcnaSWkAHsjEx
K41UvxMduHFYaXQEbHNDd67AWOiEMl8JSqTM1pOqhM1Ba5MV03wPDj+cbVaBs7EJ
0+DCWUyQFXjgFMuhhq3igC166UTKv+R4EwXl/60dtRKvu0zkvqqVQbAO3VJmq4w0
cuk0mizgIuqb0PNBtF2kfPjPUdSI+hank6TofT0my/Cxfq4+m7eIPo8a9y7Rp1v0
eYX9NdrCmvhd+ws8VDf+oZnn7zfaWK/pSsz41zqvyGnVHXojHgEWUWLHy/G8RlIk
/byETVbO0wvI3YSMEAZG7Lrzv2Kw9SPJc2xqr4GM34HsAgHGLi1UT6PMNF5+uL/y
i23A3aqw6733QGo6MW3Bhaj9ud69V/ASBSR1X4B4c8pvcf/daf3Jw52yO4g7BS8Q
hbvpP+om9+plyraXF2Qsk26S8NRWylxj036QFBInMQB8Dl0bFK24A+jfJeJp6dmH
GLvIMrhEKIirYbpcc19Bi46jagHAidAacFbSSfqm0coxaO41rAEy8jdtWdeKAeXa
h7Eo2REdpcFjRu9KTjSq7CPpQDCmqCUUB+A5TqBYcrji4r5/FNJytDezUZR+CJtz
lQU2WdK6rN1l6dFNUt3Ul7S4xzfwV1qXS5n8+uz363y7ClhjGNN7BbaNnYg/eGzc
2mU1RmsLsbbW1d+C86WzGPeKDGpRYXHLSTWH0ykxR+MYtN8UGPmraSbdlc8Frv01
opDTuFL601Vpt5e7ulFWK2xcSrM+DNntudJam6WCih+cY1RUVJgNpG9Yi3jFvaof
BC4FYwRrb5Pn4pkqsInWo/54nzOqb+Ao2hI7ERxTANKHqBz/BuI2NJpPg6/SV7KY
LETLSOKMMIU32ejlbXDXHuo12E9vBlUWh2N3QF185X5StX0GZ0rH9IybLqtriGYa
ribhtQ6hW1OIo+4imyTCViX+t/HRd14xsE47TyXTmS0vz1G4Ah3aO9tBgtTvLpeq
Feit7y18tmBRxvpWWNCkZRCA72o3BYmuEn0arbsi4SleiGhl5ERIgP91uEXgdRTK
xR27GbapeSKC930kdUnv513uIDahyo9Bfzx7uwdlu61ZSbYBtNmidb7lKP1c0UB6
FQlELefxdtusurTWmj1N1XvZUsKqgNA50x986gim9QvuD5zgDC0VXGKgGIBFRui9
bcmP203YEo0sHBP5RJpnV/M+8NEz8hINQ8rwli9Ks9Nvfsw3sT/DIHzXJ9NxYPyT
1tdwq5EZjPMgHdSDQYpoP2o9fy/crjxTTEuDZPjDLmFd3vDus0f2XCgQicT4F3Md
8Rib4UO4JFh2JbadSZsOUZi50IM50M69jVteXKzutEBJZIWwSbH9BOT/frajCtfu
Af40z1X8NXQgsnI8PVnU+XPrK/7tRIYV6zZnyvAKr1uNvIx3sZY1MERDUH3xjBWo
MPVi4nt2va4x/wXJwNSCjxLqPB0Uuqd1Y4o5fvg4otSPkavoQn0g/5wH5c/zUakQ
RqPjZxKZUU2DRnzyCiBQBNHxYtxynQxvCwjteto2Qngg0DW2EJY4IG6sCMdxH58Y
Ksh1hTTUB4y5+siRtJpIt6aY75N2SEFYYIiFQikUEPzNHKVMpm/H9mlMdJb3pSFW
y4uDNXm7SlOLf4pcZM0CRfJnJX2lYONLtHsi26MeI0I/Ce1gGIiaP7mykWfo8Cw2
FufC1fvsCImTioQeAr62YVhM/yQ1jqo8BTyqVlbQcEDPaFD2wRxWS3y+gL5h2/KR
UGpCYShxz9L40Vzsf4sqlKbpP/Kp1c1+cBDKd6D83Ds2fkgTEbK0o3MTqX2CIMuV
nJDwMxKNeMN01VqvMM0VulS5LLoR+MEX/YVa8ECAGugh2N/cCyhQOFW6iupefol0
/OpqlM3n9uacA7iWTooTQmrE40OHKkD0QVwqy5hkipRbUUbLt6EJqwAdOnBwrc5Y
n9qbEalfejIMS/873pA+jdJBolCunhIKNteYZUyNY5Q0+MhecB1tAlcXw/iAOBY0
UjVOoG6h0CQGOck2WYPSwayhtG4u6t2ybJHBQ0UEo1eu8mokO5uVCP5qYToiKhgg
trwMrC8DKmcMlFKgIKtRrpmJP8sPZ5bZrBHmp74JRXcIXsaDvey5JoiIa2ghEs3Q
LHvLRwqFeE5wREn+EPZKEGsBz9camN/3ojNp+P+PPTEtX3jYB0AGmFlstUqjdIT0
u0+y++WysRSOcyq0XGnn3BNRFRJNvuUe1usB1S+7YFZNZh97H8X04HGMoIEDTQWb
UKS/BMN3GDUWAqXL6mCj9SVeOaRR0G9QfX7haJJE90gHCynPzBIKGe9lm17pcc8d
FfB51yhFwT8ZKIjNYNT7YeP5Ixt4xMSHjUja7cSiB5FrQrL7zLB3gInxkdYip7Fy
WVMLAJOqc1XHHuPlZWX0nhw2rQcsiybjk4GboznTuLAZ/sDDlDHLt8KuvsZp+GH1
qpl3a7ajg21VoTqTNpaeUGqHyzf74Rm8f2qOiyh6Udj9tUOejhdxXAGnx1UchK7n
AIeit81/fjcw01iiLhrfkcv0OmXgJ/QEZgMbRaqg8H7RcS02mZlOQdLY9cVZ9JQx
hYkBiec/dbP1TZjlQSGxRmZFCM1Iyu3nv8xquFdFOtco7BMugLWZXl5V7mKslr3g
cXek73rsBOg772NUjRDE90S8kwQOEV50NIri0B3W0um2o9yQVN2cZXIeatg9xwyP
NB1749IWvfnuEbRaDwSWPLs+cO+Su/fCghwf1oGbqi+otIPFPKJGRkiPC2I/UiNT
EqvOHxSQF6xJcMdmKoDMyk4NvDlWCkMhIDLXZSekIfWk/WtyMDmBltM00B9qc9Hp
0CDyjd48EaA4UO5qFXZ7fJj5caBc5nUeXXOAqHbBFxzcr/KqPss04/HoinlZ064v
FfIZBrVkeXR3IKKtUveMf+jTc1s9KO/MgA5MxJYMcnuLw4C5gLCI5wrdHj0O2Tz5
i2q4MHUmHouAUU21deIjcwdWvms8xzCEbbZPI5gEXKh6kDuiSY226o6uI7ufjqz/
lcUtC1TcvWzD4vWizPr01keDlnHanYnae4SiVy9gW7PVyXFUtHhf8FZpsYLQdq7E
ADIyLZGAcGXjwJcbbuB1dinL8tMgPcmIQLvurFipavZy8/WRs74Gi3SnL9ykT6yv
P0webqLJ19XVZDOyTlFkKJ2rAjTPHFcXjGw4m463jono5j6kN555NdwZAgyMfyLx
xBeVFcohhAF9vY/QqV+exXM8qVY1WZi/boW+xAdv09r2TShlDtf40Rq1r6wFvqwZ
ErKRBMw09JxcLAn8OX+KSnG8L11QAM44BYLPq12KC3OkIsZqHxDXUeOEIcQL26uf
qroGnHn4Ax9pOjWW2zPhxi6/fRc1SsqbIN1FTUPjWEaR4ipuWpYVelJrp+xvFMjP
pMix/i8Vv2tRDY0qeVBLUrkPMeH9rvYV5mUdBM0BrYGv47YV5jPjixyHhVPQ4mVk
N/aWK/HaiH/p9k8WEEbdc47J7FmNnhTlZMcFDCOgFnXRt85ltj8vn7Gu/Ij2UXxs
LrKAn0PcxWE4Bect+MhEeDbkUWaKk77+ftSrN8n07ZvQnGAISMUA29q2QeD9DZvV
VAWY3nXJeIXnM7kgSVKDKFCRUTn/nlAKZc8O5gqoM5P6WOa2ANjmEt7+qm+nOvyv
ObsyspQ8Z+awfI+/mmCiMVMg01p0qF2O0NPt5h33rNhniOEn9H6Q7/B45eXlJZff
EU8HCWZYIUYpwsWDlVWk759viCE4Ein0C1EmPgQYKzapeKWCyhDKOW9Lp2e+HvAO
sYoIP+1ZUB98zOnuD51x+Q+ROOx1+q/BHGFVFWxTjTWJnHDx1uR+SeaO2FEKmcuU
nc/nYudGxR2CzMxuLTaOXmzwSBQZ6qOz64bIzVCbe+ET4c3HZeUE45TGuCFPmpHF
PbxDx6cGrOO6YpQaCq9XRUE6bgb6MmOLN3/D1SbOf4mgOIkP5bZY4zbh0fFsq1lc
QOPbQQofdr0+HshiethkrlozLhJH+KuNZL2Y9c7q1zq0p87FaWwxVdWKtNYuAhWt
bxJ+nZsLkoFstSWgd1sNs1TZfVxvWzittcwVds8GuyrVP6Q1ZbP8iZexYdUxYFq7
6xxw8jIkJKEkNFF61a0gDtdG5vDK+kwt038Yr52aNoxFEQTQSgagNBiz4e8YJGjZ
42oCZbon3+o76weoSrmUO3Z1+wpKr4E7fYXy5pTO5c7PZQ88whs8OR6B/n88Q9qv
y3bduvumQMFQOR9T8cSY1//GivVFA3tDWAyDD5FlBtkUsnECO46UaSwAsdOFah1Q
CZnCFPjq9k8dNoyR2UFWBDt/3S4rkbaSi6Wj1uqX+LxoUBvmGaTdUZXJ2vsNRDw+
phavIuWMYe3TQYd7BgnA2kuMMxg9nsSCfchYbeN7RkrJxqJA1zuS+nn89QWXBTgc
Ixw7yHvn6rbx+i4g+WPB5Jgqo4pfe2YftAwXcg8ClpjweNvFhrnJu+TFz8ki8ASN
b7nlTi5gXb7s48UMcN1oGOY/k3P4EQ++YWfXr9A+ZVzGP9K9rE611LWUCzjSpFpu
/1P8gCCATSz8HFT+4BUZK08waDin5Wib/yQtzsTV9wQTg45aiCqnAIln5gBy2KXa
jnY6Krzjro26riy8O9gi+xSZMfFNu5qYw5Z8Z7YS3atLbjZa5jZ3vvbv3Q5QjHs3
9w1S/iLqpiCnCUqqlKaTAbkk/Cw4H5+j9OT99rNG9U1kBbqxMQflr1DxyDa0whEb
N1Zg0ViMy6Twx7CXXLlf87wNpVSRYbOBdXDRmZOVwucEMz/T4bxk8QUu6TimXVF8
7+J9Sg36aljTS+WETjEqyfYMbtgJUD1k6O+/x1QsQSrG7XSerR5KJ5HONO6e0lC4
wHbS2BJRzYW+q/TSGWpZ71lC1+uM+oLJdxkijV/itsljNyMKZYgmcBD+1PM2Ij2I
uRcl9x264GShwZ1BwoMeblU4lkC+LMV32GI7/wvMbHkoAZIUQXTdsX/PdUTzH/gF
/ukxsZ9hYagNubJFvqH/Gy1IHXLoUgJEzsrcxaulBgLyBKQ7Ek70wFgWonO8DptZ
1PBrzGOEcYEiTmMDlhgci31C3YUB0mNUSqyyLH0556kaiR2s4jzDsg8A+1QmHw+7
KFd4OJQsk7nJ+evdMsB4yUEINcpDjgVSz9QOHW4Ty62/ILU4Aopp8Fvjh6caevV4
n9CFC4r7WH1iVpCRXJb0q4uk6zfGOGkatwC7R44jVkgaXhL09DyIezNNxoC2lMtW
vSSx3dgW6KEMzWYvDP6Ff1njhrcpUmtGUGRd0/RccRxVR/uh1O5GTn+bfGWmOxZM
Mim3aHeaCKZ/UsvcNJuoTXy78N0WMazq9eOqKDZzeWsfafQW1eJDiGlHuTCRo7Gz
t+LCjWILgyppEbJBG+N63xzgc59y+iTtIyBKHUzBjVt9Ww6YzCoGsmEin+0QVvfH
CWpJ4cPHhePMeaZDqYvjRu9SrmsL4ZHZ/bo0N6Xx1WHacXZX0h3B4SPsfSyFdxYo
inIKxHKk8+27pDESrR49iHPapjb0XrHMFNMbNANRFKTMP8jZ5hjkg/QzMEIQHcZN
zwOGKuT/F+2jkCIOM9BavIaTEfp71cFNDzQPqBoDVdPO9a1Fn7WEhuNfuPaiuoTu
4+myZ79ykaYYa2Y4RLTnNAJ73uGCiRuoEvctOj/+u98iQS02XH44fh6sF8tz6Wn8
QfHJITdFlcd6IKoUADDpVuxfc+tQ9OIBEO4bVNVoZjnfbvXCqmB8ym0+85JTWp2C
vf6XrOFLqHNeoI6f1jEw5DsmZQEcif+JtWi1EHrfPzZz47UHd/G6XH2Y1OgdT5gf
y9ILQ09f6JoGf6fcItUViI9J18U2Dhi5xm3uvKBbPpijNE388+UuJIdcp0JaZ0II
L22dg80Y8CmDURFx3P0YDbLv74EZZZ39NbO6nVmy9+UZ0zdgK0jSytxhhC9IQJdi
k2xvvrWpOCfeYnHI7fPdWm+3KIrFLdaK3IDxpxAcwe69xhpcl4uNseaGzH6egPvj
hRWlamU68AIe2APFiMwbr2J8nsHWAJzs7s/9HExN/jR/IYrVzIsvJCRKqT14ArfO
h9v9rVawdua+V34g/Fk7PLfzdW6Bj7GIQN24kFedaoQJUGU7oWZD8jjeU3GgEepI
W7D36HTL0Mjs8LlESc3a3Rd2r+VWE0W272ek0bjJcdsOFbH2i2u+8kgpsta7LkEt
UXxKnjtEuHklpuhOTX8ni/8rGss35tU6degiclqjvD3oDt751sj8hlSrq3heT8iC
Srwkj0MO8YTTKH1O/O70aZhFXBsmQuIfC7B+rwhwAD4xQncZlNdicIHiH0SKyzfK
VWSrhjo6FQrHEAmM/2Qa8u4z9ZQV6ZqXJVffn+rjY3Pd0qXRo8t1+j9qGJo7pWm4
pLChXFUD41/92tX0brbdZPG59DEeApvTI+VWwmyFJSPBGq4GM+23pl7uLkn/6+wE
XN8O6tQ8Y4kN5FQJvHN9wmNeOgGo8NndF+eywZaT8dWEsBlFY9pUo0WvWFZhAj0T
saJ7RNEsYntPsPL76Im6RXW1Dad4enY3kXlHCxQR+4CQhvZF+9ODvolps4IPd88/
zMC8jBnsaliluLyRDbsyhWA/js8BS0Sk/3mHe+0sZ185FNZGdDg9i3t4jC+9isbD
wEUrak2inuDpo0jZ4UQ8EfM8lGL0ecLR1nk3OXzcZ73RaiXGpe4wFG25LCgnf4XF
D5yS297Nik/q0cNkjIdY6cO9qblhRBHbCiLWhi6hswA6sDC/kAbUZOLs5wh5KWPQ
VQxAUqnGGZMnYKdEV96dhNgGDhBZUcCfr8j/ZvhUATkXt+NC5FCE0IzgPBT9TJRj
CF8s+y+kw4zF31iTjMWAqUPvV8FT/Gb3QmIb5riK147XXAVoYtojgRtsf5a1Uoff
ha50cmWmfnimvxUu+09AtprQVRUkR8VF/hf2Be0TOlj4V16zSZsLzs/PFN6KP8PI
3N1ELKzDM9osQNJHDijSDmexUzCUpeVRcZxntFQPyrzkW9pRW3rHsWk3muQ2Cdgw
jAzg0twvmaQF5AyRsMB2gXzig3ldNSPwW1WcUZmJFK7PmAmCsyEu8YO7DDaKkvIh
amijOsI/vGvIfGqH8BLLyukpQu1ZiHOYhfHzFP/4u9sAEiulVykH0uFrYGvf/wzf
HYE+1wBXAP/GIcz6rOAl50JL/4vPMwLts4WdpxMG647K6FTmfsSqfOGwsTK8iDrk
L00+DJypHPMl68vqF4NupzHY92jPpFr0s/5nMH90sgYvYEpgcm8fEryn5Ezmkib5
YBublxn0ylMrMhZdW12w5BvWnqBvhTZZ1OWWRf8N/NHmM84iJf2ZAwCzJ8qYWZo9
pw1O2gWitC8QYO8y7Ilhf4tqr2Zs629ke0tq/x/0fS4TE92+iCAKrpw31Jmub+Q9
nRI7EsHlL2PDgw6oq2WL+IBtgyMw5qef285xHHcyYoMQcZRZguKjhpHzjJj4MkYW
aQS/t8ZAdAWBHCeeKcx47upG0scbaHP7tpGH0L9jZYrK8OBes3j+Gbjc92XEDw2A
9lMt5my5R5hg1XNdexZvOeLkdIk02B6Xo4Yl/0gB6CacCh4mjbhf3lRw8ioD2ORu
TbXTE7bl4NncTZeIBG56b5MQZcobFKHIZjYmVOXXi07NDVrB3t1hXtJNuAmrtyH2
N/ZMFR2OqolMbYzEIfDim0OVM3XIr3peM4aGhG5ea5rbSUQayTcCDQu057GmW5zH
+PztrR8sGRV9KXzYXUcouDtf035Xbt9a3lUuL5cbSnJmBioaW3atZZpFVpZbXDnf
LSqqcMnSm7+dP9EQeUS1R6pV0jFjHWdCCg2+GTlcos8Ryt4MYgINJi6FII13eVC+
o7vLi7iERj/aak30/fouTykDTmk8ZJn27j9od6bWdajwGAjL3/u2X9vrTsapQnXE
y+VnrdJe+iejjCabxJnJv0Lev5HVS8MB8U0keS34B8x6cJNmnDb4JNlJ47z5Ebmi
pX9riu2IrsosB9wZ018pXbwhgZ9zpDwkbXoi76pM03qCXCH5si5N6CDh3LahhrXy
ZipLcLgRHVnxYoMazqgfSiVcTcpNyVOpkitPhbYjL/BLGeQlMoQ3NqomerXCUqyZ
Z59Q86RpsIOoMF+UQzJZzwrEhACivr0DeXT14ZzJpJUrDvQGwvVpgIgPgufPisqB
x4Q4+snJ2RjJCw25fRLHaIp2wFQat+0K/dVkgin96ac0yQs52oEYs7ZblJCTx25i
5+YWcY5FBC6d0q0gXaKnqTVy5wtuvMExt5dAFMFGt2/7p43oeiVxs43LsFcPSrKS
lbYFRlUcSrR8yyPvysWV2XOBpJ55DNt8UI17Nmp1lDafgaMSjr6cYkatsXxrVsvd
uPNcVoNIs9ItwThjrci8i1FK5lNuKbVYUiRgx3cJjAzpGYoPCGZC6X8OzyzZ3TyR
xgQl/FsBf05Z0QhTC4qWfxXav9EwR199akCAAoNX6cJEHvDMSIODbHuTeBx9MVhF
iYgCfUVIehlPezAARgRKVDoRwFQoHYq59i/9qTByGINS2b54nFRgFeKHcamsbHrQ
YlBvbvwY6/fXHAPSpr2y9NArwnQTNX9LsujxSjVEqZBFqU1ZSCMBaOtF7y8ws9Ju
UBpv6yE63KvUiMNOEzrJ6TiHvKNFUajl2jyRnx391bP4dOYzyGCkZmD8LVZCgaTV
Q5H3ssH0J4VzFlY8YHc+fVSU1GTyfc7BGceP9z6C8os9flkGAklUANap66B6EviQ
H4z5m9pIV9PlFuJTpjIrH9JKPuefi0M3x2oUz5uLDF8jhUKKzrmOT4nRtcZdZrXW
JAPefv8+WSS6aqcUVrhnK53awCYdTsoZCKJT7KJILQz49ttpWv7ooIiU7evB9Hhz
kwdQCNyFmCpvLUjaZQCMmzTQFp+1QfY4BNeX6qY8peCfT+0o39qwHWqWGYC4zZZk
YmyK+aPQ+uii68YeLog6hTybnfO/3hpoRk43FGK1ED0WZmsjsOxPd0arQ7Iu8ub2
GxlXWfh70/YgrVDY2jIQYIdEsFmBlqMG1a4kI8cyOW+hdvUb28LsfklnPzBkc+fV
X6ozFCt5d5HhL8BvD5LbFM2hQ8jn5zDoehOeVQkiDhiR1JjG35NfnIydkSwbxlyZ
f6nWk3ufSysZ5gTH12nfQ+HpcZuZcOiefgX7pueRJTPWjBUd+kEcrzBlzgzdu4Zz
zbn4bx/bZma4EMn49LmuHx9q8eF/SmoXfQpHTb4iVVjhy9QjSgSHondT5pNKc5Wb
yZlIVoBnt2sn46UDwrXPGC3PPtBktFg99jPZzOICFrJoHbR+PY4QBhHMScYu11Ja
gSjQW6jpYYf17+C0uxEHHED1iHJlksHEHebd41R9cCY+rV1Nk72lqS5DiSib5Mab
JcFfMYihGJhivv7NEVbO0PlH0A2hBZ7n1P5pgoxY3d4lKeaPjCbHyiTLQGEXvdn0
OwawUxsol5qRNcKwZjFJ3rFD+yxOb+raQmjPi3mKYDpTySBKQaOyMa0Y5jKZJ1nr
ziVNnPCQ1o9yHhtTKEFqWlOVXYOtXjtZvJE43j9fyDnznU/ENiyygAqj32give5p
NI5/qiKWRbT4qmgrwG7j2A+l85eXhbolnsTf6rmSV3fOLdBa09bpitp+1lkYbvy6
PaOOhYmeWSu79bzNjCwGEnbz3+xIG8WsBgG9ouqRl54z2xvfFSVPc+A5WNaMKOf2
/H/sgk8Ken3E36LTJGwkC4LveVonMFT6PxCMAfY1mfLamjYpSH3rZW57peG5waAl
EAUeSOJwey0MsDKUZWEl2KFVyc13AMVJ7IZkESIZILW1hQvWHbAAj9darxc9Y7Bh
HIjU8/XkN7Bv80oJQljvtLbDD+mPmzef4W80glYaCfIBiW9xmUiFii4Dh5Tfj5bx
pMLwBA71oojzpKkcMuim0jMRMCKF8MfPTRdhY/CD/gFkF/u28SKA/44mCD85ie4b
BNeLfHlH44ErVSW8Jy4xmDXFa0jGX/2e7fVyYpSJN4Unq40fL+8prae964yI0xfI
3efXAlX2RKkI95+yPSFyiCNxQmrnfLsD1u9pvfaWB6D5nj3qZGwehfpgterFxV5Z
Geh2Be/2LJNJJX5zykLJHQ9NyYQ/Q38wAY/2WiJRpVNLgdfZS9TEaeppNMmK6eGN
PYcDaJMFbtiKccEJRTXC/SL+5urnjJ/MfH0UwQ19iUF+yqXg4knysvyIV2Tppoep
Qo9nGEfO4pNGnpmlKYtXf+7byx7tQUXYMQZwgDLVIgxZWgil9HQW3S91bJtKfSFZ
dfsKy6tmlJNpykw/2IM2BmYDoJx0EAD4BKtWZ9ff5VJL8HDyKIt+3n+nZUlMhKHn
/b6V7Mm7vUYCf7WaCTzYIdh8ku5obqLC0mjp/a800W/WUGUh+AZYGgUv9mdIQDN4
U2APv7YRD+nKddAKnOtiB/lIJ92F5GQIVNQ/O3DlNRZJCGNDj/MkRLyFmUtYkLvE
fyeWb+jCFKiqbv3gyKwVZOawcsRyWOlLhZ868VoPXVc7kdODepO22oPNwZ7xupCJ
zEWxNWkgEi3d4/WlBR/geJ8larrTeCwKMidzuGzVnViTV/HCVifL3XBtLyqQNeP/
vPdCdRgxgYRDMFUx8IXMmEIqrsK8OEqD8a8d3Je8OEkyfBVD0mDJhm1pA+k1r1Pc
LJ0l43/EMvP5nEOwK6IFjpV28T/d8Qrcd7UzgA95Zh3p9rYvAVJKi5OHxENS7SSu
LqjShJcxY6Oukt15jaB7Sk7NG7wpERFw7PQNLyJYOOtlmuqrk+zPuh9CTBuV7Z+i
LJgf6wdq0H0LMLlumzer/0oCxE1XZ7JKmD81vKxzH6wwvNcPfJU1ViIJ8G1Njb8v
KVmdSw609F9BAEKxSTsJxWahVc4Mfe4aWRFWw13KeqKGgJr8y7kEa6w3Vte/1XKu
WmUQFXxWBo3oSX0aL2lu6GYYjSbxmtMN0bBac2sZHxE80HnUlLDdtiIl4M5pe9dB
m9Kf5aIX12numSQjsUbzyoQ8EsV6rZaktAd04BQNYQS7UMtkWL8f9MbXRoGVoD+S
qdfLrYVimXAZ6bTRIUA1ou9ftaELF1eD3FdjtM43eJoUI/W1m9ik7dOWRTL+4ILF
16mWrTLx1emrgQusNxcDi27wyGD/HpbTGL6bkWXeCa4Vbhe0cU9Qqr86NaoWIFnn
0dv+JvvYiDELGk+m1Olx4Nx2e1tIwTPAniMsKF6sI3vHOvZk72r0vtyq8wFz84TD
TgOxufXfjT17ledUD4ypdKe2QpNgAP3fm0g9/ra9+UOPKJjCpDRNX85ow9kxDXIr
ulG6ptG4rwNOO5ulm4RLuX4HiNjrMzgn0EzAWInelCQUAori6AO+B6l78ZoAk4Yh
zQbcFePNJO/G94y+k2NgRsaVhkjtGZ8P9MA7wVxqTmXE1o6nDcB0m4a+hZAxwDcm
iBHqNP2TlWonezhNwRUdpg04DAeswMF/4Wall1RwkxL3+K2EZOOyL0BbJiRyxqFp
7Xgm7V9RfwXkdmkkM6WUw9dcfOkLIvbAbXq+VD2YnI0GrgAtyTpbsx2Lcv8TUNXi
FPQ8DJpQKErI1vHKcknPvgze/DUt7yJa1zkqvu6YCpaxde0EuKz1zkMwqvJa/hKO
eCBGBbnn9lYpV4/ucImWs04KY0pvl/DlnGVcR0uuEnJT2KmlTCAY947yw7FpTvqn
v6sPouOxHuTDcMEpRI8yrIvrZyMtOT7UUk2Ps4q1ddhblnTJKs95eU6XumZJQHfE
p/pmQhVf1Jhxl9WPdiK5h/poaijJkVFCQhqc8OiDmEGaz1tc5vu1SnmfoagC93CR
N6suAxwpo/Y9x46v8WY2Ipujp9dbLbDM7mUUBzOyRsr4omV6OeMi33xjyZPgMJW7
iEB0X5G70P17vyVoBd/dv49l20JbpvX8rFb9Wrm9SmY2lxkaAVy0vn6gxwACI/rx
lskEV7C4qCgxl5hh6ynTrwbfM7VXa6LWICXrDAPANb1o67bi4BiJCBqBAv79fPh5
Cfros7oXkNFausn7uvYgu/x3IMsAZn2rRybEXPdSwVx/QiUneL9754VGO8w0/m90
KH11Tn23MWk9J5PBh6J2zbErFxEITYR8CoujDi/E01/r/aw9V6DfyHd+agmeKKdD
18ReZHzOzBTP3LoahG90txucwJJ3b60WZc7Xeen4nD4ZY8HwHpK0fW8geVSN6Xrc
AXcY7wLudb3EBjjuabJAdnPW9uWH5oedNtJKyjhJZ5TEy3N2NwJCBhfEblPZyklw
8xGSaHViFYuJ/qo+9rN9yHl/9o67x2FNk3wApXIzarAoZnghyGK94ykY1bxR7LFA
CVuEU2BaLnrER95u3LRsKSiJoQfOPkF7NeUtc94s+1b5Nra314XSKp39GqgQdjD7
fQfgdY4MaoAFSeoNXgMuRy9BB4HlSl3MqXZdWAhA4wsjAr/43lGnDtypI66lO6q3
OdkPebTqGg9OJ6mOeF2ih09K0wPs4aD4z4datcfh4LQ6zDBl7tq06deoAqS/NAhj
yoyKKdTa/t3PP/Y1+f7Ncpu7p5pVE3It/XDb75ahbxpBtvcXtID4QsVZVp0X25Ep
+G41Rkz1xjW7pqU8WUY8JVlrG+HFkJFPm2BIguNk0SiVjrrws/g48W+7cdlcvvW6
b6TYcfZFdUNAv+JqevcooEVFDrFInDfn2I91cr7eoOZFGI7kG+gtIEXZzyHlLPuK
7iEX4dwsg1vtGhbsS6nAQjb5jNwSZUkTaLf5Pd2yGFTvH3mLUCxTC1SnviMeKXoD
TwTg6WzGUeAqtxGCoRIBIzB3pMCNhMpV4vjvZ0vpMi7uDHdEPPUsvt12zPwIG/i8
RmDlAodEd0dago798wZKOEJOG9avRSPWdXekoTerrIBML9yFc6KehFzR2O9UvHGg
oGTr38cj7mkTljdepbGGRHRnU4wVQd0zOOK06EXDhSa6EoSa49gszN93UZmvyG+H
1lfoqlORervtXh9fY3WyE9zwMhN5A89N5qz++4YdsPZ+N8BwIddG60Kd/wF67q2+
LMQhIkNbP5YUDrkYNxekjmRaW+7lJ/1xWwgS3WpxZ/dkZdfkY3iXL7KmAvh6ifBK
kFpo3pKVuHvLaL3C1C2Bfc8Sgxz1HYhKG15/vDgvHMXVMeMyb/3wgH2yH2uSHXTi
bB4IOez0rQSxGzMEI+EZp57nkgffOC+uXnTY6mrrh5ZgbTs6fzEI0wQ4n2sb6RmV
Oi6cixe0cPk6KmLYoTNodTOfiOsgyAQZDyDYDgjo2ldlzUBA0Qr1SmH2ILh8L01J
oafOxWJjxFzcmv+kqah7kCd61q6dBDpAeGJ4mXiKZmDPaNgapXvOkvYVHlbk6Gni
oH7bEdw/fhNrqjePIP73lvOJ80krZKlIliPgBCUaXf4qldkSrG3Z0FXfViHnfBZh
Op19nwl+szc3KhuQMesSdhSXWRcVKaTWTyOBnDh5yxkyTuersrItxfubYvjr/yzj
VuUXSF2ULpst+fKDv/pBmCbWEriXcW6cMe1KQikEtD5OtkLVmn7rX+XUqhIEKoFy
eo8xLIVWtr09XE2ql3dajgxhEmu1my5XF9JKAfwBftTHScJJ5i1r8SGz0VwZ3H1J
a6VLJnHcYS6xPGRVE6gPe3Am0+nUCfXFnAag0M3EEgn22xnKvpJbu04Pyf3ky811
gGPoIz2RjMHfMSfw/l8+Zajw1+zfLqLlAY6bhNClOHNowZwhW7rztF4A82Ae5rJy
DRk+owBtACIPRfB2D76NDvdijV4jZaRzd0btr+7mF5hFEeV6n/p9xbn31A8uE49o
ILRxzaxPvvvizSPsNARRQdoVrpYqqgJqcfy1tTBAxjjAzSJiqWsBPdzWXVESqNQ1
tKWmjKdZCF9DYPSlCZ/QaimR6nwiDcpvmyQZa0oynvqN43SLinXzOjyS3mdHiIuP
WA+Ug/Ka3r+TBS0n0rP2aj4mm4nUVPNZDO96XIY6cUyngOprLA+lqTlbW7SpQUXW
8MpZI35eWXWaxhs7e6r2Wkd2JpxB2Ed0o0YvscCRrCfyFoE6UUUfKMFd410pffxV
KgFMkQkVCZH8UwpRZwFmKPyBrBniFFwFlqGYxqiGvsITaMifvbYJtuyGOS1JszcQ
IYUfEJTxipzx9ar2fgi0BUo43+EZZxSFNe977Q3rWYIwaksiZNW4DXuZNRu8ZgpS
LN6eO4U3lFSzkSVvItCVYBsSVH67r0jJFHu5QznZPseU2BpmYBgp7PFHJFxBPkSP
rU4JJdjSHyMmd7xT5AMCBaBcXv3n9h+fdxwXQYEcgO32qC9ETL7MqJROVaLfAoBx
kO4zg/yNZnqz383D3fjZTUjGwXsCwDGqBWjgFIqKnUsEjOKypSjMwOzt2tyDT137
8OE2YNcW3nSipmykIaVt2MaRsBZDnt0VxH+tjne095YivK+0fwY7yun2fvQrzZFw
SFQod50CFCq3yf2zCogkABVOMtdKK3OigVJQyPUTtGhb8wzGiCbYvnldShQ99ivN
DoNkimO6qd+m98jI0+L4WVABjjHqX45rMr6uaUYqPKb473E80rY6sIbb7MWEXVut
5Xx963grRNJgVUKgCq5aWuEqAVV3l2c1P0fl5rBSc5cu8bhtoLfppSmW/8ERokcb
Zbq9e6n6Nl3Olr0FTFwSppHjc4qSt6qQsUN3g1wVsTAt29VgTLGbMrUJEvNk/kHz
cXm0rsjeDfGZI986/P04tO7Vk0jS2Bz57YauKN3SeTo9pwo2HxZgFhDldgkASkIk
i0h/3l5hfbDK56xKY1RYUkZK743GLedGQa+OztEjB4WmJMBr6vrsKW9D/6lWtu+K
jh5Pm8sNZxyKyRbMOaE6S+AMUjm4nrRogIzC4H3ix3gH78h7kfAgajztziAJlZh+
OAEvt72vAewQEGa5oDpMox22Mye7hWe5EAfNiBeOPF3rVzuA3uL1LZ0a7FdbLvxU
h76Gb/1hs7KYRjX44qZYtzqTl6TvvEzhfj+w+2URRtIIumUMEDg2FnkGZta/7utp
cCv7eCSD7zKSKmucQ4ohu5zhrPZr7YTzXqeiFPK6c9/SMYC1EhkfJsRvyaHqpdTT
2lF/VU75JFdNRugSmk82lBoDz8h8Yoi1ufJkmC708yANhgpQOBW/sRK2x+E33f12
MRtgp9EI+OpesYh34wc9GY38zLa0OZNaBusDtwFvh4+IiJoswsau3GkoN3lXQ1Ah
XogTBq2WiSXrGQSX+BHZEuwvOjvWsLozVepSdJ5A+Nx1zRUPYkW/s/jw+1NIHkaq
QgDjHTmH+0Chq7aV1/yIOCsYdZ8Uca//cbhxPXSrmNydlJEvNO+FMWTwO7D+GViJ
M9tYNMGWOw3loKpZci+zdklrWU5w/7iZFV7jrkCLZ1+6f1yvCD/ftYd62wvgwXkY
+yWWZ3VHAPjnX4QQy5ReflwPLssTtjU2eD4QjtF+Dwy1qLabri1cXF7E3luN4X2p
d6uokLh+UsgX9HHA4CX2oWx79wJBWUUYtA1F8BIWz9wyAMIP0KgA5aEF4av5D1Xh
UYdaylHbQC3yp54eXXiblwNVmoBhv6iYVz0oSD/sYtFhkMppCjkN6qz8ctv5C2Gb
2JTC1fnVd1qkfQw0ob8P/zYq3oiFReLzldoTL1KfXyZg4zn1s0gDBE4A93dKTYxm
mMaayP7UAZm2WfFj9wKl5ay2Xp2x2MqLRISQnnvq8LRXET7PMVgGhj9Pkju8bAdx
xq+EW0bxe1iLAoBd1ps+jyXFwU/ku/NxtSDcqbF+Hli+eDReL1FtYhzgPI6LpeEG
JgFJ6GrdO4MzZm7iOj2xFMAIQLffnZpOjiwyxAETDqleVAW67V3rBaO33G2qOhHL
HgXlOCF0RJ5/Jb+e6A7Jxsoi3dJSmNeo5ZHehKGWI9W0/b2ea9GBqPXa1cPsVFvi
LhUe49cX7c78JNsJv6DFahqd+3r+yt3dEe5nNXKL1zwWSgNCL4EuyfXwjsxWjUze
MGYI1zGvfCD2quZguIzSreLMRoWibXiH5r0Da5cY2JJVemtvhBO+jyVULEHmMq+y
08UPM7BciaUjoPmoydEv2YKSGbSRuYeSkNDUNxJImAiboqzgAUos086JqUIFOP5X
1Heui8qJF14N24etnbd0S7lrZF2IGyBGTEddUTNOJ+G4a4KzeZ4cf/AXsE8Smxf1
m82blZTrWY/0wv8SrgtH+n1iZeOURcOl3n7M0MlUoC9QdtqmhfnsPpuXhoyxVPQi
dLlPobOnFfapOL8U6JR5eVZTXRW6NwdRW6pAXb8DIU580FIcKFzBX5071lCVPfPl
91BPWPHjpAn9g2/CJXkTSS33u9HPfUE23K9jo7wcNLvXeYWvlOBHRNg90KZKz+4E
9OAStRZ8DgahIXgRt6wR5p4Wl1Yix9crjPhPfCbS7BUDuBAiUVneeh+CtlV3YxC9
i6xKqVsX8Xi/FhgYMLNZQSIHhrPr3GbHXv59fO7crdUEy44MGPmHx2riJLq5MfZf
TxQfA/PGmomq2rh7/aGWZOpk8F5l2rx4Tt1RjsdFkFdb413Bab15Zc0dV/9YxH5t
btBiz52zqSlgPcl6ucKYqUSmQSAFJkq4kHxiFMJ7uB5hL6PAR16sOBEoaiAb8E9k
uYgQ5SxU+eVNFvcn8xB79h1YbKupRL1Uj1TzQl53aGK+srAv14czWwYv1PcDLg4z
/3g6g91b9/Fay19nNtCd4lg2NOvu2HEkaWMm7s+QgvbrC5rW0aGJqbb7zcj3rReJ
oVADvIWBhkaqbV/kHqn5gr8RuF8tBUHJQfa0A/q/qlAUpiuQ/NXDToPHTUE/vVVk
iox+dje6WRPXbn2EX3ru9KXcnti6Fca7fqm+11cHOw+CA/vG/hNeb+rOShavoCRF
B8KiNuJpm2AWSAiL1mFy6uFOnjzVPfwWs2Ub3BsHxBqP3NHj0lC22Z4yt36XIc3N
F5b5D08PfBQYEaABKUOi0ZrlJBS41Hff4wV1V6b8olbtb9FkukC3ZeMkeDv29kDG
Zqi+x+Mqfk6+BUjBUzuQgWn+8POS7DdlOlZgR6TDASZFirT4zlwoGk/YQd0L23JS
Mcw8pdpGzq0Pi4W25s+MXJQ8TJm3oI0QWpFaJV81yyxGc4EH4AGrAaHVShd2knB6
MF1OjcKNgJ4NUDmoEZSeaDFCxutHWaAihqUBpoqNsPRtFiRYDLBEUH+z8y9eKG0p
eMTQgGeHDE6v4n4L6RUR6/3J0g1nh+r0mIUzoPaLMhPnp7CEGeZNs75urSdWHIO2
HSeEJNldpuFaNqRFhGu/L+acxLxaFgV80ghEViTasGmNjEgwOqRhun41y4aZ8UGm
BJWQCnGbBHXgMBzXluAPn934theOpnKPM8LaS1NMD1mxkCJ9zSrZGlfOvGqKSOpO
XQNlkerA6vBDwkvbeMXvjLtFYB1m3jclHnhyBtelPjbWCqMBElml4zxbbyDuSFWs
9bcs0irZaNaMLHrnmw14dWhYwNU+4Ir5pDEG5iwn1Ui+/K1i6pfcGseKHUrSHHl+
p1t/MTDC9l/bybTtdfzICKWFD9v6RAR235KuMy2LMHT3OanWlydNRISrCMYLmo6u
/sExGMvtLVBCWonN4HDCLGpnTYqpmW/Fh6TlRxvJY/TEUTgz7SFFDiZ4osve7aEp
2YF2ZmOFbb8oclnltQM7e+k2qV4sjg8b4ISEsmdYMSKOW7GOP3/Dhy7r+yHxKR3o
s0ZSfr4MjkKaB6GD/2GENO0I+9qpGW6sbRqeoPOLrrzFLXykB4uPSGrTuO/X2ydT
wKQ6492Ku2Coz+Boi86SYQNFwQ3v4jlOomZKh/d0xPS30FQ8mSCojUyo2zDo8cKI
A65nSe9lqD+hXo+Bdjww6kRPSdGeu/3fXS3vsh0FyR1YWY5Yt7n8nIx2mGgRX7BX
2GwfifjpV/vUr7msHwhF28a6L3UiEYO08IvEDWN87x45mntI4HtaFkITRLWhrDZO
NMTRLRbCyof0LyO1K7Zvp7T+pe7jh8ZDCQCcYkkDN0rOve7QdHeO3ysLsBpPlQR7
4Cjd1ZSkMy42ti8SnTqBkjuglJ8UKoouEEmguw+Xw+iigvjZeh4PXTrxMwGcbsTI
gHLK9SEIGzoC5G0iMEkri1CXFFbeDrWYWnjLjOQjveFEc0Ca048k1nD512h/kqSX
uhlgj/02Q/bDIexWtRyuoIjtpbag2yDTuVoU5amHvckn20+pJAUCGebs/QkWKWZr
/YOUadkfoMHBr/pZaqLxzWkzvcdDqNMdCgIYvvH//FIMThs/HzEVUzFMEvIJ495P
QOk6z3FlpODWF0raVd6cIsoXg8CrfzdB5bdaUh3+wYbyqJcp2u8lv2T9+4gbIKHt
s6KHAMoqJDS/K0hJsAqIUMXxyHV24DmjZBlt7Ytk8SEXrDkZhtYSy0qxTF28sMdh
NAoflIKHEYzTg2O+lKNPuuDhKZ9LWeqRLtaiSsVUH024r2PI0AvnDfQvi2WnBREc
oiqkyz//ld1PppHjhp8t/qWL6bCGCMGZU78BgoETsFoMnEesF06+0UjC+jVNSlMA
YprGDtc461YrxO78yOv9vCYwqZQSVC4KjWoNjrGSore39PgGMRYmmgwQFB2EaQ8e
qOEFnXVjLKPdcPZts2tFEOhX8sPm/L05ftkGpik3XFEcnti6c+Byh8vPAidb7iNe
IjcbQbRDULKFGE57hXoCibDsvGPr/QBLVbbM9eQj//cOzvo9iyUEZ6GjoR+Z/ToD
XG20pXP/QKXwUWOMYwgAmdOJqc0vfMLleUmdqqaV5rT1ejOWOrcThyUyr+MNk3D9
+q6LJxRTMQrQJsbtL1ayTEUzRaLHg4x+/QMhEADMGZ7Ebi5jxcxi47XYH3tnBnXE
8Gtfmu0I5KSFLm3O9bQqBV4eNxV7dP99ZKdVbGwhlB+TNLCzxWk6M5mFfYRZz/BT
o6kUc1w2x46I/PgdNh7hMiUonkBX3ZMZsyTM9XpZrLxgHotn5PpJ8UYXp3cm8LI5
om9v3Ds1fHSDUebayJKb5cfIgP97d4QDKcAF6FaSm8wCEwQSWUXTZb2UvhUGuA61
nH6EY9GPBwwcr9JdOq1bPrxAQSRfSJpGCuYZcTVX5JB/okzfUo3pR9BzNwGoFKEN
wsO7h9O7ujutxZbdYssotoJbWYCLXftS1H2jcr+dBtwqBxIZQyU1pnrkr68TWiPb
kuz21QYWYYIaOE1DwNpsBofgTJyLu47aYxBIO4fMvmOvuIWaOQXFLI0ChKsW1woB
3NcgvvEqsZxQF5UKCwUW0SPBaDxZ07t3AB2J2pEYCSvkDjlBI6smFujRolnVJiK3
srFbQD3F4Hc4orWYqCUqAyNxbGA1C0QzwmQBa3zYy3JuOM69squAPIj2ZpV2gU73
7UdVXqrFMin5H55KON7An8vjTKVlI9IYqn7gPN0d4JQPBzhCWJgyXFLDi/7mb+KE
cAZzOG7/nXFZEgMDriUgbavLIlNVeahxBQJ7gGnpU0ypHCjsHwZoFHr+6A8fKKBu
QX9ozw8AdJaROUlTBC4spRqkrmiR6VySiOUMkrEe9iRvIraqSakH22dFR/o9fnaR
6K1dMy0PFFAYPQ+UXz7Pt2nzjrtInyvmR36+aWv3gSLqtOgtCK/oA6hnlL8clPmJ
VTUb+MzTl6gxhqLIZrM/genxkswCnqFkMp+rRavXzzAVIad/15KIoHqg/+ay2TB5
r1daKZb5IBG6X5gI0jMQAQLP3/HO9N+hSoZrN7Pnwh27plvLDZ9tBdeEnvx68hxE
YWPpmg3YNnAPmZE2P4pLl9QuefAeEez/AWxcNKwHuW6Pc1/ebPG/Hfr2m1YtBVyP
aXmx7O4GNIsHd08FPhMDLT6WnbT57eLACA8PAFgcCoPqj64L8d/ZCLOixlcjQNZU
XI1Ui1Mwsb6wHS8nQeluM0QyLSH3/zEsnQad8B/6gaRqxrkfBqlQta0Hs809CzHu
5wdKu5S/urvgQS22BPYsIkl2sFu1vHoNUyd1Z+DuI+eYI9nZMspX9tMPh4vjjtxw
uU60C6GfPbrgwopdViQatPKVBCdJN3cynxa+Tnf+4+ZxwBl6u9lMkXvLRlLwD8mC
BQO64lXt1R+yx/4fRHBhRTY2OTEIqmykLI8pEjvvdR4tsx+UqD84bQTqG+g0kqvJ
BcB+tLwLHPkmJVRKOWYprqENpuTw2rOT+cbrFlN1T6dxtQiE4u0gCYl8s37R0emH
SCde7FFIqF2XG0yiVD/l/UxJa8G4i6M2+MTzOeN0vwSvLNDLDuydlisGDsyqmjn8
SjvCKPdRfBkkG0zGir1p6ta+rQBPI1Mnyx8hDWz9innmA9KBTsBPNi0Z8kA2MoRO
hOW2eEg8EN/wIMs860nR9DgYilZRuZY4WMBql/ZK242CrqXtgip5a48OruY5oMoj
IzYNGs1eB6b7Y8Cul24P2qGJ7F2A34ex3Dl10fvERJGOnlICScHyT0dGeCqgIh0p
Cx9lwBPHhm/QIOzzs7uMAG+nAh42B5DvnfnpCu8H+gEHmEeeGtV9niWXPXOhpJtp
P58748Z/O9UhziHRQAksyZlTXDZNWFSd8gd73qeRRr/qTB/NaKR8MFcgAq5/KvUu
T3hkeDl/IFVHLdfJVJymPXdjoM52iDlggvilgW81xBC5Pjsq4hHi/T2u5ou3xY1A
/+4RKb7aVrLLIiEuUL4afLvDzGAcXPq1GEmYHnEqVCOItVJvHn5zbWz71/RCEcd8
RmfetDdyhrBjm17ScBkYcsg4qs3C8dvJ1qEPHhchOyFslqMzrUVdfUHC/gHtrX0J
uQRVSac/jCYvYdKML1SqeX3VNImlvGM7FUoHyxZsAZcA2Biv2FtlSUzPUuS6sLRc
Owu+ikG6nunBJIJjsKJszdUZejIFh+GG+9oJI66Km1qG73yVSwfHH8wyTwTaoNop
bGOFbjXyk+w0P41sqS8l685zuCfkqcsTHbo9m2jhFcVpssnq7INaGUpGD7qGGrGQ
UwG7/NkcftlJdinbrrCuo91td4B5LW24P4pr8ruGZMjETjQp2+MxAd5OdXJp5rtP
lyAYOvNRUWPFavVtJqUxqReslgdGLhpeK+I35ghRZHJoXsW7cDRL3MmYXBA8S/6N
BpZC7SWdXmtlm9yCY28HmQs/JB1ifFHvatoQ5yneb6BiefGU7q/e4yvpnWZWqnbt
6bSBLLog9xJQkJnBPj3nrw5nZLRg1DpJMKcHRAeflViYEpIqgDzv5BAzzE3TywEH
SOKk8AeZwdzbB0nUcmorIhg0/J2G+MjmOenpMnzYNaoajEH101+0CZwQnvJbnUVM
s3SMMdxjxI3145MP4Wf8glKqje9D3xxQOhxZboCHGX7eNIV67p3ogb3VPghMvyYi
tJF8mrvZh39oAkTLlkbkuzIX+x4sjTdPO3rpqLOXMfGtgE2MwpeKea206M2o/5dP
xVAIs2UbFzJtOOab0MogJ1e23Cl8baOByq0nBZTj0Uzcu3yQdhkaxVKgZvYNUaYc
96/m/UK55E9l4p+jQrNMtNqPjngYCfO0EUfbctw1VCfgdsq06yunwhRIDftHDZ22
5TM1E1FB+QniovRAFeAyL7P9/QE9OFiYRPgoxEYmUSemefAe1jJfe1q6SwkmbiGO
bHd/xpaJvrYTFbYeutdQBuywa+sEfEgNWw/EPCEatwQQJx0NU9vFxY7BZBIGjCq7
AnpLwC+jXQ2DgVn3AytXzxYOjmRCLyYIz+X+VnW5z649/BZv0uz5z6x52Hz92Wsd
kLbl3sqwmZm0W1qmFxNm8eG80L78BiTWIOjifvnmCU8H+sv9TLfIUwIvL21xTMYw
VTIF9teIv7SvlQjZ4qALszEhRhG3qlPDl/EaKGC0KBJzDnuM0XlO9ftvJ2vUz2xc
TkRajk+AA7Ph0hGNiuH7rbWK4HV3xBAT1qP9KmQXf9WthvFntzOCvP3DDLhqHMhd
HrIgg91bipuDxTF3RlMqSRVPqaB1IVG1YAV3UO/NikurARVvEtQR3PEqV/1vE0fS
WJu0zYWCHNJROVjEMkRM1lDcL9/9xPRx9cvt5bnz+mjzCNn/qGksWPd3nY79h7G5
L82+cjZE9q5FeaWnfAHRqVIrZ//e78+K7OtBTQVlOTPFWndfFU5L8kBjcQZ+c3ix
B80nzrFnt8qJKUlu4B0vmTMvE5IVdZpRE0Gm+hhL+vUQ3qCRymI41jkz4f8kGORf
H6mtQDXJh7QBkTig0Q7142kDnGZo5Vt4Ix5kCOZThAAZmNc4QZ1ZHeiFxEt8uCPL
PFtJvxH/hxRSGLmL58DEOrYZHZ/8AlAu57xgM3SdbgzV5/1OTZRSAJGwCo0u6aSa
h2oUxNzxLJeIR2fOygZceZwBRC9uX9hKKadRcM07kybcuMi/gknlfGG2+EZ8TgrX
TmIiVg1H+IJ9DGL80exL2OupvIGLN5Pf+6O80La7LGyFWuH63BnvTBH2kfHB8A61
KRSMayUy3QAKY8GrJXYaWm0bLnvZbfFg0/0njM0WD8FwZqkTncFe9SAC0j7JoAVb
b1++LbqildZykCF5jTusfqs2a3OYgLeZX6k/HkTrn+siC8i2wc1MMXzD7ktk5J89
TUOqiiVmxEVUurpu5F6cIxKDtGgaibi8bjr9nqQLgBdwCPH7Lgdk81vDAkdMWELX
OafrzS2sjpKIeih81UV73QWbL/h4/hXlfd7NaB2dGj4UlnalPql7Pmfm9TAxPtWc
SmJxg5r6DPF/TjRvbFaT//pUqi0tD0o65d1EbLMfhjs4mw/cZZh4Z12YfQnlptkY
4oG2TWxeA7TTC9AyP3zg1x48hoSbvNPXCHVhTfUriSnt9tgy+YwzPigv4guj36Rk
uslVnuPhdudLIGi1cwFGUoqMufh6fQgcWLZjbYzGr4WzQ+PD/j/M7NizzG8wF+YA
OJQT/V7eIGsIHcRAJ7gizWnXi+0rXrayebL5GKuLWLAKrYHhmIRk/hd0z+3XW+xj
IygmzHTiY8wh22qN6qtKM6ZCurAGY4h0NaIIYeLfKEC3EmGrXDhML2vngC3D2lmw
ozrhXT4+TSvmh/e6lMM7aVzmzYx0JlOu4/gHOD0y7N1z6q+eCo+SeyErtfBdrbE5
zPVcS+hbG0ExKY0QcpR0vg6bu3+3sCMwTKbXpJs0F4umbSl+mLBr256KP/9VKR3j
5RuIVMY7KikS+E1XBkEzxeEru9bkwJriKiUyF6n+6E/hy9iV1keSHbzwvZzoQVDl
blCAVqXwZq/cX8UFecjSJG7ACeKk2pWQyYBhGAzOgAUx2QLE/dsfhey2Qmm0Escd
z+hQT6CmkhZLM5wuYpIFEdDEoXog4jXfmDc9ko+d+SZuF4kuSWKOjwP5ooGa2KRm
UW/r0DJTCckODFGoHn19Vw3cWyjCoE7yj3b84PfkCIGl+RSRxND6+6eCCIWe/SK7
56ebxOmFx244kx7oUCvKHUOUDbGYuz55X17orh5huFWfkYy3uYIbWho0+Mn17JkE
6wsblR7pfyIP8Q16tIh2uYqCn05YNKRRMBXd4X4YWcRHglBWYVkX88VQyvRNVgRj
8sDzJulKEN1g46skOmQpdCBAUCwfD9YJIF4BqUYEMEM/aMtO+jwro/QUPE5yw+3C
WXaGggn8Kjjy9wgDtbKzOmW8ZVUmrmNzgPNCUTzO7Th8KWYFfhlAdy1jDAi0+U5v
xWGkt8/vQQIwYLYvfgQlLbL2wTFAs/9hYTRr83krHfgyo70AquV4Xo90ODhdFAaz
8WxT3C6A5rBWPAHhOrJgiVlOmujP+G8B0d488rDOhTMZ9Ts8YqeQUAGSiFU2VZcc
6o8qBkrmEtIuLlnGI+rQ5OKz2u5pp03hTmMR0/bJ/1Fr0GYu2hGOGgVOTwPRzSYA
LDJEeLtrVPBn5KPl6+mMHmJcvCcZ+BGSQhls0TI4HnI2sZH3qmo08PWhWorCWbUv
QYmwVR+y26bNiJeiC31wS5W6+3HtRZagizXZA95ZBQ0vKvWLDBczEIb2ur5l0WaS
wNt1eH0kwsOdPTaYFOWKY+Kt8LF93V6y8Sx01kE88u6mZCVktr28RlrJ/PxeFH/C
6hQstDAGzBkWSrxyBRCMc5EamDoKkCNsvBhyq0R/VQhqbZGLc+BZJZcajjTMCSTq
0xn0OC3UYDbAFdMyoyheUndlyP+Rhm3p2XxbDTE0WxMPz0iZm2dzMnm6lGlfHhW0
DJzl2yZnxyghDKi+QoKFgGSA2ZvMJVmYseMA6XfUBrV1mqtmF7tQu0Vjhn0Q6H+u
6Re7yosUg6HA1R0GapoGkNqwNsly+jbQHo7I7AQXdSlRM9VvpVJgLD8WJfkkmfmG
eV4P38E1bBwYkoPDFwQFgD4511EwfVf0iw4D1Q0aWdWbesKIlx4DUyqHz1Qh11wF
07GmagffCnPM1qeftBvYExQUUedgEAC7POzqY9H6UVpManT88hCVzxsENJiB31lN
OjuoZJqdzQo0/50tKiXyN6gav2lzuQYK4yPe7i6LMCc3PKR8OueyyZgPAoNAYiSV
lbB4cqoRa0TxLtfeinG3ND5JsvD7FvuW2GvEtmet2hNr29YiUM4AfzsQUe28LHW1
Q15PdT+qw6rZXCDFET7iTYhtih3It48H5cB39HU3aNH/C9sy7FqzfmW+u5W9OrWp
zJa6rN/59MQ5Ll+ojeQg2xpLkOr4ICDjQFbeMO6JcWYJO8FHuZZPr0GXB9cSSFFA
3pHhwTRM3gedp9nhb++3PXmv08JZ4kxLUdoZ/rOqvrG2cdqWOSUEyrpqB8Ta5lLx
H5I6SJHGr+fUfWHGt8vXtamdDvM02qVnOF7i+hivc/7itx2LBOUaC9FgPNqIr+LE
xlNrsW31tUkFxUzeLzumIRpzd02mgym5+hsP9l8EuOygeFV7RxRh07H6gmfxyRf8
kkGjSN90K+k3WTRlYyzFgB8rBRdsOrRTTBIihxaUOXSQyqqNsqjPK3QhaqcpsrjE
EFNFG6/DDmMDJOSNJXf51WGjHCEVNf3D2cb+DzLjA68YPyK/FUxggJ2AM6d/F8Mf
Pc0cq0hNJIm9aA5XXQdC1bCkNoHf0W6QH6t7CK56OWyl7BPyL43KE/lP1mfObRJN
t0/TDcq6dh+hPJMleIs4n05dVT/MvPhT6U2tE/Wkjt1hrWkHP6KYF3Chbb3csuWk
86OfqISjU1BE7spIZMmNEJcNROKDvJv8GaaMdSDyz9v96kxFPCDQ1YUZi3LnDkNb
IYWcLlZTjXiYOouUNAKIDR4WmiWxqnURR1DRuqV07RbaKfxpRKNd6SVNNyZVoVpd
FcCxl9qpbvLfWn4woYGtHYlK3wA6GpLBm10DJoDYMnxKqyQ3TJfnZZW6dh7Nfaih
gctzbW1I1LXczQoBjP2NF1nZ6evgDDAe4oY3ZmDGrsy5gLYHs8gXpZm9IfExMG89
Hzj77oM3ANjWmEgDn73UqH3V97qWJepB6QjvEmafkA8HyZ7j9e5S8RHY5m55lC+k
0T9FgCIGzmcsfh+mYgfqIzERpaVaH79k1ohmCFbDhj4raqnFH5MB9rREi1DthTCx
exnJ4BDigEdz4ek9rJHHJLKDv5g7+xO5XqfU025BVNIwtWZq4lhcBdZ7Gt8P7RVP
ggw2EZ0q3jou7POx0E0BPCmoh0tScDJot5dpA2MVNwVU85np49MPR0GoH96cPAao
iEOQ7H/tpUvNh13eVqSAn9Ag2ui07L49TW/AsHQ6ZRRmf5aQg4/MN2I3miYLqLIE
Q/e9Y6nPF+V/kbKkehCqQRY/f8KMvkE6avHK7S7+0x5Px9tCd6p2ZNyIergeVcLw
DTd67EvaKF6wvQp+toB2fHJECAiyZzXxJboyXt+Ib+ASGciOHngPmLVxUbdY7tLm
rxMbiPhB/3taeBcotx0puGWUQdiC/xlCG6wWW/yuMKIeu5CFlQRg/V3JsdTGwzt6
6NrLL1TH5EkzOHtHmJI4HW7cT6Xn6m4CRlD6k4CiswK1Mt9jnsptttLlWkK3EbWo
xrcG1ZpgzjHqWJ5SbTXxxKfYX11C86gYSvIXrJYxyDxHS4ZR2Ffdm3VXMJQuTn2j
Vum4JaSh3+dk6wCUC5ug9xc6JRzch4spsVDUjBWGjW8JhzSuQiT40kMjmZdFriQ6
cFCMFkSB6PP63jJWJEHoh+S6KBWttlHjj5/3WFJR76jh0NKX9Y/SJS8Vzh6LnDnD
GMUWCZSC8Nbzj/2pcKLmeY3/ZWDFMifZudCFiUmjAmdYI9CxboARXg/sltety5aa
rfMNI2pVthouM0TE0egEglcOnNucJAThk3D/ex5mamSf8JXnU0rqgN1B7QY+d49k
hMHtqlSTrf0FM4zQ0+eB089F1TMq2GwbXO6W4ZT+bURPySgrB1Zi7NyqSclhhEfs
AVcK2dc9jzYipB91/7thFslEycQshdtvgvbAFIldhOK7K/eo4K+3rumwVF2Vk9GW
8Nt+1bX+Adc3i9yeI78yWn/XkKYspX24Q7TafChcMqEmqelonmCZCYZ29/zFPkXI
r02eK0aYER/ucMXgomlBViUAWP3EK2hZ5fQaDlu6I1n4KACUStEB9DctG7uIy55+
jG8QYT5eVd87QlcFG0igV9tBbD+pTeF1fGUTkKGwCYr8DBo1tr7FR87P1/1wAHcB
+SVDs1YLMUMw/5cr77nvpskwNkJeRorpsGlu6ZyaLSCDh1MrqVmj3FxHtTMyrIMF
NtQHZ6qGXygFrPUFp5yoW/eDUDvhdv7gfMnxXW4/zXnECYWkl0+TbikNd5ndM2KL
cC9zepRR15ZhlM/o1M48zYeEkoyB4PMUjPR8xH+asf7XNVhXlk0EAkFCNkdQ5g9H
bS1OeMkqxlaemhM3yEOTGpjFxvagrVKh/jz3J3+SkCC2n4QVxYV3xiP6WHht2ic3
fuJqnbVAvnbTm+ixaVN03zNJgiqcjZ8VNPfKhw6684KKZGgZRHSz4HDdqwpmfjOr
NT8v5dpSg+f9DOAmBDzU/k9HBeE9WvvrTDpMU3NGeXUG2EU0XLsrUJXAZymWyzxY
OXn4r+YJqxx24lJiFDsDdp0iJmU2iNEqLt2cnbhTWYyTJMMeFiIrJxLz4lv07ZJ1
k6ZAJQhWZ/lB/RN5oI5C8u/+nuwcZhX5NLN/zyluioQekseuoS+XYrr697P2ysgR
IGIZAqvqW25gJwwiIpmuD+7BxkJAZTOX38oL2BOwbGrmDqbFthPLzO/HicIBO35w
fAB030Kxebj7fwKTKYwvUhTI85FmWBmJ6mRMBUrACE73/9xH0UEzEG+/KjMlMkZc
scIWKry6qoQ4NO07dKbeGnDogUK/YFwN4nQSZAByd7IzPLoEVTT74dKaHA+hbvEt
hCjkzISA509eU/AWFBOStqqwC2co9+iKpFlX5sX5dY51YfObYHVkakDC6hEr3NQB
izQTAiqkAlTM9mo70SzfzNS+yE12wLiXVuiCt+9+co2I4vNcDsHfpkFXw+GdF3z+
FSY5PLyotjYKF5WqsPT1Ixcm0NOJ5M8QVezzQZG1RsU+3BQWS9moDD/FG9tZ9y2I
Tp/pirakkMuiCDxqZWDQl619pTqk/RRGRMqocLjERsTrTwhYw8WjOFC6t3pq5uqo
cOg5czmPl51dUNwuBzSES0qjpMhP+u8I7f/zw8YH4uv7Z1rZHBV1mcLyTe2TiS6q
R4snr9oucAsR9pt5+ErrBQR9BnatWA+eU2N7nSAuO3k7sjXzHhKfXj6UAmm/yFxI
1Jc5JbLyYRP9b5WHDT196CnflfFuEe36O6KnDCygIFGL4n1T5bWZYA7PSvpYpn4d
oY3NA8wOtCneeYxkcKPbxz0jjZ2xCe8L1FGPiHF5zX0l/6GCy+5tn5o/N0jGtXKu
fRrTFtdkDGM+YXPTGKmKyLBs2k3MTdAY2A8lNK8Hws4O/SrFpSfmqmJ86xdSf9/W
xvJaRhycOHDJW+GOqt11SSiOS0R70hnhQXrBnEbFp5UCSeFB7wFsL6OifUSZ1iBF
KLZ/ptp65qgKA4xrfgXTlZ+EvZMr52vMZnE/cY2S9yk9c+hTHlOFe1oac1G3mVw+
l8wimoyjzWKNJwhXtdvfX981eImI0Zm23VP31v2lEU3GayBmn8D9DQk4H5o9C8Wm
OeUm1QaKMoYQb5QoptYMSCZL5qr0THZO38u1m4LhkUcBEMMpVLaOQhxMxTTgnOyJ
EqsMl4bOvrZQuDLq2sHBlwx2EEk2g9eSrjo0vd6HbLlPHpT+LXlTTtihuKUEZL2Y
AR4uY6nqwx0XqQ9J27taso6jvAHSdtE3fSea1FcSz2176NzZ/6XT/ufQWeCenx7S
lhoX01qDqw0RHTv3WNaG1VuNs4+0CXEv/wMuH3C3CZ/Pb0nDIabScAqFEft6Atpd
G5f9V+5RzavF0gRb82gl33Gh2+Gipayxj5aVuYkeIVfCj5xxEeSCUoHVZRfSdz0T
iiMp+cY68BFCwyQEs6tn4r4Y3Ad8iMB5Iy5jeLzVS/O4LOvgSkExspX2PqPFkQjX
X67W2LNwdxpYQUXYRJJnZ2xLm/OpPjBNV/jMwefO3kHgkrJp0vbDVEWky/t7PmQg
F9VBOOnULxS858CCj35Yw1c/trZ/fDiLpCa4KH/a9jMDWhe6d2ANszeIQgu7bDpy
oonYRSCyYCI1oepPMf9hsvc4vhggpI90oFZig0wZ2SJv7Tj/CXv5dFD8dbmhmO+q
L8yxMKVCSjxM9iCR6qHuNRJkcMoJymz9p3C43FcjGIY2qSv/m5o1juWPUkAcHk+3
6JazlME13y/CVgQn4D4Qbj4KEI7qH7216Sg1TxfRNwLsHUCMCH5ENmvPHY9tRa0C
W0w7ywVRWnVp/g+3ybT6PaBo7DlCGH9JEZI2p2migAijdEPTVxRlUQt7WBrj67ll
rIXaoQn70y/YmOzbp+IH2QAiHmTB8WIQg0FowuIhqxUCVopms84sXEcoiRxi8BMK
mYdbBn/oBSsyy1/8tfMubI5Ob9rhNhsn5zzQ/7ezfUPKU3wVLje+sq/1med7kjEB
hY/clL/yPMZQE8nXqz7eXwUP1Rb/hhU+Y4HhEZR9xHzVC4ILBi07ZqQ1q9RcwfFt
I0H9Y/UWp3AaHaWCMRAYXcdZMiN74Ogo7Bp6vD0motsf1RNlYZMJ39z7AxIAGnEj
SLLDhO7j2tSxgw8ZdmFZS5k1UqqYMslqSnBwe9eyfKYMvVVNGM3A4UDqh33deex0
N4HqNVW4lfCJ4heH8qoTN06sSyFjzH7FciX720+TyOwqCsceL1qChuoMk95ISk8g
DbBv3E2hl5le7ExRe/cyQb5YnVwuJ8/jH5RBPUyVHUCMDcu1q0uWtHBAFXyH5fTc
bWwpSNJZMrNMhNAhL4nTb/rEmWtYwwVHHv00x7p2rKDmynVA9PLKib/m1kYrVKtc
SUZBihRPFzi7JGKL/GGB2HPJtxUv758A5xSmrqP7XHVQQ7jkb6FJHYNwxf80BbE3
QfxiwzRxF/51mMJl59AjHYsj/TGFkKnyshFPFA3+MrubDf9VzIOAaXz8/ZuxNu6z
s0jBq3qAepC2/ieKUTXnLlMebHT78PgXWSWpRtFg8gG4P4D+bw3YLoHmAk6X1zd+
WVJUqf5IJjLc+Tp8kKJUvp7Q0NhAp2M61v6DfzAUSpejC0YajY7eMmDeRdTtlMpV
c9wKsDodKv9oCGrOvReUIL/Unbv2ezFPbD33Zb4C4XPNJVNv8HV6SS+bYeog8+Lj
8XJvFYCikoKL9DsJQx4VcqLNjV6rgN4BlbkqImPBo0VFqhtC97DQnr37Av5OwGkf
4w5v+iWlu82srNHpjlaGfY0EFEgBnMvVkB22ssMKkzxVLP3Dr9BJY0Z8r0/QSCsR
vZ328fXvUvK53NeJrC7QkkBStyDhCcmMweJpXyz3EHP/BFQbS0ZnaB/iPnH/NRCb
Ai+r4Npjw2edpp25gj9gLfDLVypHwSOLXaJ0F3sFrfEj/GrIPAU4zeg08PFXAzi8
0yCshw1nogPKpvyCszFs+yOoJpqplL8LIH0Cq0rdV7YeXjwQWVB8Z9M/fA4bbfLl
gQJkPzq72ZmC3YLlCSLNvHZhzIkC4U0pXzVaLZBE+YHtF93ejwotKyry5ipipVCO
rrSkagNStrf/AL5aCqWUXpDflwTsjvFZhFwuiVQ2OL/SRUQAuEEZNQ6ficzvNefF
Io/ia7wfO/dPJBQ24wDLco2OdXLbMlnN/0jX6rgrVjHTLuOqjo7SmRY+DHzPeArp
bk34f84iurEVHGtqYpVE9q4ciHhNq9zVD1UrPABOUwLc9kGKfhK6YXpF9TTUFXf5
zgRoVEL5Vnn++gWrDDJyEjdghMQpbDFSlrT5/st/cfHVgFvzG2jObd9dHQM5USRR
bpvIUllWmm9dunDm5qY1VYmJmQsbQ+P9LAhkaGXEPbercd/LV1n+5X0mq72wF0sU
ECiqpk0Chlm6J7ZgkubRAJshrh6+KRyHliWO/MX6sd01zMKgHYguXGzHGPHwuXZT
9rC6AzoGVEm5JhgD7WMHKwaIcyZGJGeMZBjv9cQuQXd0JMzZ6x+MlRsxUhDobkzy
1hrH0fbtARmgeCzpsLyBFSaaO/JuY38nPSBK5QE+Wr+Ymve1YbIuy0PIRodUNKrU
/WereWbh08YG2Qpjm3mXxLxpo8Ha0LHeL6qvM6xqLm9D6FzxRQXkFjmY907h4AlE
CCDlE7JFvl/JlcviJnvZpMLko4Yk5SLHquOS/RCIRh5VIev5EA4bSgrOthJ50scG
vND5wHVTUqnzshSQ4yYS6hzG2ozJEY3jwq4d7e1Ec5EirDKkNy8ZsdVJkgX+fU/M
hJSBSgMIZaxT1iwW/LbMpPQCYTG7CNx+1sN/M5fsT/v8xIkmlOpu5FF+gH0jxTDx
pJpn1E1EcsyROtec1Czb/Wy/rWvqJ0ZWC3PwKxoq86FI9Ww+mKbZLkxqOvhXC2P5
idEDDwOLLPIq0kZSojNreCT8TxCuIaP7guU1alIOpnFMAmQiSmjDl1voTS+ktC9U
OERMmaI59ZVrbORuNHxt8zQTry2+IdNxlyHxlZYhEghP9QinDUS1Qs+HBrEDIKZ6
7NhNbRdIuatcYmDFpds56KS7zxitPXXDma/c81LSF+6BayuQVjulKBr9TMJGD2Xy
ebjHMnc3zzBagNqIg+R5hw8WeRltcYQggTXlZekGzzbeECY1mwuf7Veo+T/6e43C
KUo6XHIF4BrN4rC08ytmKXnnMLuWhJB1HmgCdIXzyx04fEPke7HJAT9h4bJJ03B6
muP2P1hnsC0QJIzoU2V3ArP2n22BRWz1V5A47fMmfWvq0DFKimS8XeE7kAFuOxxh
2dsZWKaLcNjtyxmWFGnkrBqQg2XTRbh/5FBBNnMx6MWCGGovu/gopxTcVXbWcraO
Dl+e54/+vercgSG0CD5zmQDZ6FKoQcEkOi9AjKsEYy5NNaT7joqTA46u7o6EfILk
87SyrEJkeebKUf5f22lSjvlHZh43lL0QpCg4S3B3ANcp3wZXkBnMPi+c02ABGpN+
xKhbDogi7b+lRMX2BGuC2kcf5ZujX1HIsC8hbfwrn3oIC7dsgCQWI13iEaKGjGi5
YCr9VOKiwGERaQu9q9SeByiZhM8z2xyNfpktQ7qjk0BFDiTzmmVEjWjK1TsIcShK
9nC6EP1Z2ukzHaYAreIx1DYKlJQXeavCAvfMBtqS/X5YLGxK8dLdleleo6AnabVR
RA0JOnLnU2Koq02+/X3UyvrQWSLeCt0xM3atwpz5m8nJSYR1P3w8YG1QdQvfZyyv
7LpUkaU7mMYhpKsh8n/L6ZcyMVNyUCiLYa8jIKWeZd/LtUlYdPxn5GmTbGtLEEEW
pvZDlFb8zfkG2Qzl1bKhERCFa/zqIgBc23J0ZbSpChJ+vCaNNm0+sCkFTGNsrRu7
ygWcwqNB/jbpGftjB9hq6eBDw03/iaQ5KtZBh4X7oXzOza0zVv/BFjPM9lDszNsI
dYbDNovOw4IRzMChpaErWuX+kQ4IxrqwfLSAEKG31wSPIR+HqstfQ0D6zeYlm1tb
7MEXriMukQOGLRoq0uycWqZ70mZYOJLirIgBBEdXyqelqHDx7sfMagBKiICIRxII
WJK0PslLL+lEvw7Kqc9r2s6hcZjhfy+Qj4wYGnZ5UEmjt14U4PUJ+vnc6IAa8PFj
gpjkm6Iubcl69fZgXB4sGcDqe0e3qxE3ztXehZH0CnT1JyO29Mz4GNbiqSQkshOG
890l+MfwDf8RuAnIw91u7GCxPrcEF28bcOeU1PiqNpjZWwfEzhJSdaCam0Ld/ptD
r94MeOJ6iJAezPyMlg5p2tT2JotEmLimNZHhqFOhTNUWbRWNIDxqj5fS6J1Cb71a
wIOWfl/mgVKYJhVgdJZASFJjYbSft2LlbLtrOUIAJ9Bpi/WIWrN2lTRadsfZAXvm
BRcQloHbAIP8cizyCH0DDPLnw8ONouqveP6c4sR2B1C40OZPOsQJ+QWnGS1bQ0Dq
Z8qXTWN809EOnXpDyOpfiNnJecd3DGVNfDDBvumKxdSm6rsbx2F2CgRWaD9CKr6k
7toYIc/dwjIAKULrBGEFNXxvngzKRv/vH41Qn+pyopg13R+rRkiKEDCRhAqtQXm3
d4wy1oh1Re0FyVdoPJUo933KwXWLCCfLeIIfHbWMuB6ji7L8j8eq+4Bo9+sJx1xx
3CCE+hVvDZGucAusK5m33He6VufbCYuUKnKEwnO++A12S3dw1lPMWeOJjvQ4ghrz
E5dBrc0weOvhnLcH8yMreXcYYVTQyEjm/cVDDKmvp628Wf2jB0030lPTcattg0Oh
NjIvXbtVe3qMaZl83E0+b71sEjkVtmcHqEqPlWMCpjhggxPEVkhS36l/G22gqTN0
9BU+9aa92P2PqWa2hlg4gXmZVken88dgs3ROkKRAjUP0DlQKvuliiFoLt479xmBn
NqXFpOITIAf2tyBbbRVtZ6eDam1PISopwt54FN655N/nhYLxVlbISeaAIHJ25Ulx
uPeKqcPjGmX5Cz/gVuP0VrDzy/kxV1UYvSRls/Q9acJ80x1agWdF3jYiXlGfui3X
YBdsXpgqhoRKCmmCbAANlcNdyW0F/ansVEzUiEBRDMEbexOx0uwMcef4KQL+48pQ
O9ZWMnqzvdiUtGhCF4ysqfFHKlU2gzNiGz15GSITeF/EvI0BIG6MjqVuFwYsKwSk
WMKATml20AUVg44EKum5WJvnmRNdFvQjjQTvTfpgkRvl/gh1EW9nwWwtjH3WxG5j
+MHcxzLV0Adk0w6yg47mYzkrnDzoTeAm6hc+esmlfYeNEwhipAhb6/0+AJNzpVVJ
eVv7/biR9owvrPGjjbh9SEB8StHgOuPBfhyvWZ6xrVPSSBtjgjEeH6pzLTrA9YXv
YvBhC5gRa80hDQAr2ljp3ZHRxHYYA5GQKzb0XpAsUPtSdfkzBBna6RL0cQk3NcAO
B400mxiMNGQoDjlWIcqx58wGkRiribKrgp0CgQX1H0j3ts7QH4Zov8b1IMY43CpG
VxhL19Cc26TnSm4mjTBh46Ngjad/X8/m+/BY8dP/PsF5lHv/9RolbiuVc1Zwmlc3
nI9kaPY9jVGc41YHzZkeY+m8hGk0pNXKksHNnjgs45hJRukj9yVKV3/7WOXR4kHF
u+CuL8IDBnPI7P71mRnuLfm79NbFHlYWaP5qPQfeV3SoM5wab8x33tJq9O/F92Yg
Dy1+pG+FjyUdkYxwVlSa0LB/a9HeYnW8Lm1md/vnroL9y0iPlIyWwyb5N446vIpr
DdbhD+UI837Ee3XKqxogGnuuZoEYwWqLUV94pYO7B5BZJMGo58yJ/oyxcagk48MU
1jvi15Id0xvf63Br+z2yvXDx0Y/jSyH2S0Wad7eMviYAaGtE2YvRuJ7ukY8dzApY
Pin6oaAjjtFPY6cUinnqJpIDGkVOKsIZAKWamZQBES5uU6Zj1Ob8Kg44vz9E538w
8UTeg/4J0yp9Bw6CZh0tU0jFl0Y2LYrbch1pXxBcM/LrXDejZRPnN5uTWGAn+ha6
WmDguuL9usO5o4OgopIWu/tE5a3PLzUIicyVaPFzvF9h124tben8h9Ipen8te87j
hnxbZF6bkxaLrCX6G+6In9p5553a84LeE/1TTusCXJESSUbEChfyudrMY4D/IHXi
VBaQuMPPNRSKb5FcILcrsi0R9kNKfQKmmsAjlm/EeRTU8xvfNLLogOnD5n2+PYZ/
FE0gWIjnEZfFcKp5dTMqDqbNz6ANFXUunlqUTKR0ASkAjGWBngvFdMyGTbaVeoou
lyr4dn8tf/cqGSHcinew3Geji1wVHZdWvYgJsczXBl9y1YJt3RDN6u/KIBsH6t4Z
MiDbm3aLvs+k21fU8rMGtMRZobRP5yrDjltVzYbzDXHBAok553wT3ZToAB2l0lrO
NsIo4dF8VHGSymzOzf/JBuwtJpPitZLYaKIFFB25qzhNPTgsL8LVXTapmkmBffhy
+AprrOQ88Zr+OYgeggKYvUEqQY9r7LnqroxPPALOys6XIOVfEat7H4W6NJoDXVop
aQCmYbTYfXgjVkW+lVZdLX67Mq4PdTmlphm7ajwY6pQlWWRfkzkvZWgfvUh02xHH
kQ4gIzrWNrtk/W0KApOpwZaSRNRG5uw/GUT+G/C06SwBUOI4hj90e8U1af1mWbz5
qHJ0xTQzGoDtK2lCvOyTLC/bv9rnNqR6N/YcoKj5oE2BlGkDNxi10KQfLn47F3/u
ApkO0BywFFzd1nPMRPYVNzYOmhqBLcWzGL+RMBskiCB87QgYIdawgbcqf9Qr83Ey
ET3mlk1SYAXavRjt7LCkZS5bsu8OmxxCtXuwoOX/DRyxWADFnB58bxZrMeS0NDxO
oLBza5XtM7nkFk5+qPxMhl/Ves/qMwDnsHo9B/TaITzADr82Tx5PHB2pVWFK/rl3
lkSqup/TDoZEQo+rerXS3ONr+38a0HNcMstienJtRLZi4GOTexAFxnX7CpxwRUYE
MNOSufnCIaEXrpF3EWrnO1gZQqZZAyNk9cRLAoi3TGIHDfyJfJEX2EZlYS2E7TMg
L9m1TVkz/fl1QpIeQ22cq7YUonkBFjjYJ9eJxuLDz1s/nPiuF4EtYSnZ6n4zaT/r
ws9vdTl+2TmPYEG5YkYwY3Ml0Tldf1qkqEEehA6FsyGidS1LvA0/KwLcsCqqkgOn
A+btSd71CE65+XVx5yxoG6a7Gb4kBJcqr8uPds9r0xHtxqqBb9blMmxw27pNgH0X
U2arIg0e4VY8Ye1c9EF8WPbg2e1jxyODDNayqKTCxzrlxa/opDogmuTYAoqK8Qi1
uepftPanpYjfArC1uJzj3TQv1iptIsR8+ZzDRDyWahQ5E2I+FthHGSyhsov0Shxh
ItgeNpO2qeJUT7q8/u8JbOwPUUqOnsFVqbW6eFOdE+WjwG+OfDJkvGTtFdyJvcvF
yu1vDCDMJGLENv+Zi/bA9ZOWfERVieFJxEc2rTgXwJVCuRqAQ9PMbPasbKFnX0Sc
4dEP+dcYx7eRPo4MYvJUvA/p9TYrMp7dqyL7iskmCwyQZCCUpynVeYLyUb7amFfO
y9xCyR2wPsvYGmh7ysZxFb31ab0UNjzV/5wRweQGLTpGavOnUcXCkv74kgxxZWP1
/zMi2uR3nnAcALQQI7RSANzhfMYbPiNSWJSHI0m8PYl9oC5mTsORx5DW109sAOap
sMSHqwGAyOavtLMWpSLsDoI/vTP6gCkHMMyK7chacyBB9wKBFfc25BTDRSZ1BY9i
kjEbfbgTW/kMfZ5Y89YQYDS2eWGrwnipeNcHJPv7gHM1sxAFjYujPV979hC15FwA
Vsucn/9VJjIC4A1IhmxmEjnKWgORD5RVviJmuP/RErNK+/MSUVEp360WeiVCz6ff
GV9xi9ntefdz62ARd03ve3b2Ot1fbB3ysDgtMsAtbtSVOMovLQUGZbuL51+MwxX4
5kYl7bwfvqwvmEDzmQTbELB/ONjytqMw1qVLDnf79Chlt8FOlDUKzva1y/dFDL8r
6L/gUMaiXv0JU03NsJliPiNzh9BKPXB7FcuyVBqtlsPUI4/TqupNJdiuhbvSlzf0
qLGMgytmZvlV/0zKHnQhMWgQo+dL5CN5jD6m5s0k1dYOUj59ie4zACvw0wFmnAt9
tJJ8jjMTftD5BjY770ASz3vrHBc19AhgMzd1EooO9NFOHaUySqQcY+Vkk8HMxO4O
p++TSzROdkkCAL5S0GOwaZyWXgV7xcaBmCTZhchM8KAbtlXaDeVcZBSOU/8EFMKJ
ntneQuvyHdbbzHnyLdXx322LuX5GXtY+1N2JlY5mJGps6BXesOTHNtY6vdAAwqdJ
MBUYKV7L2pxdkSPUdKjHeUpP4UJeX3+a+26c2zXHRUBhBBHRWo5LueWt5bZ5QEKA
MkJgJ3zMi/ZtdY+AWP5XIpJSEVmU+1f+/eF2YMztEhHdHiGWn5hNt9b7KJeCdY8Q
vUdxFZ1e1/4Qy/eID7H8eI+o6bSCqgnXBPuyFEXsd4gXKKYhzoN+uLGWQwJf3q2J
iNGHBbmdQNh5B6752qlkki6h5i4xL+7XZnwdV8B47y638GcWiL8GU8SnoqYeZvgh
3lWucamW03F+3RDW9ojLEwY+1HdKEbpCp0PYYCszuOGFO44uSPPU/k7SFj/xBqM2
lrogE8mJTvdJCnwq3N7ui8ehF/RSUO09yTk+p8Kl1nlP+nHQV8BpOeC3UcNfTZba
Jg8/qB5IANov1SbWOhRvIY7jROybjGcgWE95HUwz/9hUnHswDxVyFpNwxjJWJP8E
YOCT32+j6oIYhT/zywRzsZ7sDb+ok6kJkU1TSsHyUcpbIH04WxWfdgIrGIVM9wRd
CkQF8uOBoPOmydehlZX/jTn9RHHbxnxKU0Gdan1EkDjyeQDUmfKlvLrRl4CSFW9U
Wxb7sEH0Ha5QgtXglpSlcFTUCuct4C1/Qh/HlHB5tEdc+KhXO7a368dmO1cb7e4Q
GE/0ocuakuBzUepv+BNF47VXvB59ibqfQLQuNC+57XZghZJlt9wsZ5L0Fvxldr1d
rNbgBcqg45KV7bwMlMEF/EEBQ+Mzv5Y8xxwW6Fjqc9zbKEYrm1KL+zD8Tz2BwFtH
twcob8mmDFhvX305XamjO/MBVrnXXvYITwVE83vAYWYDV9MhDJ3K0Z3YE/E9SalR
lCbfGu1paMd9wCMtJhofukYO0mDoIl6wl79kYPi5QhKEeAlYPKhFpul1nH4v7w6P
gY6niuSj8q4SIPeXf6PFCYTZvCXgucrkCgGUSG+PZ/91yoguGoROWBNXwrrHF7CT
oA7kG82Ewwkg0GYM+vddlXxrImyV829cLxbbIJ/i6E3CCRXdOFycnwhG+1jtY3Fg
eWJ6QbWDeAkdF0UljfGoaTe0FUcEmVzI033yme/6/wN9BYXKP+QTayOW49B3Wxv8
z1Iu/HIRDanwJUbK/StanVVG/BIw9dAKB+PciGnnmPE6cDSpLeK1Whu9ujH538q/
GH+rOzrpahcdUzvGVkRboRF4i/DB065Vz/gDHklHe9lh+mNdDf4z5m6n0lQJLAjR
Sa0Eh2qxTkSxesTeXzCLS6U4253dmUOn3mc1QzglKji4wsfZi1dZ89Z2S/0ub4gP
ffaQZYeUwDSOp5Nh+dy1lO3saqM/sQt/HdkKoW77BHKj1Q+iRpoCFlBm+RceKJQS
zQynhtedOrHb90yGu/Q/TtJKMKOIg7zfeH2kFbsUKxa06IQbTp05RqCQ1zioYbWi
gcIyumX1QBWxYe1ARI476Dg1vONXX4RMlg5Ug0GRZYA0O9kBBBbcmL4gFe1n3rCW
fiGvHYu8WVkc+Qbaz7Go2DnovjB81658JDXHsXxD0Og/W1kkp4enmRKXGeY/o8yS
iiCR+70oBSJqvNFFVqoSS3qhROv9j/4XIb0d96UIUpgliLg0L1mkg8isnet38/QH
g2mab4e+XF0bCx1gS/el9O9/BNT6EMNo3YUQmY0VctsdIqlQI/v9HP6lOTJXACnl
EsSofsA7X0S0M5quqUrOCcfBHE+F4B5224tPXmC/9nc9jSiDjWwWWH1SrAZEB2cp
TonD+KFsC6DXLE7QPGtYsUQ5VfRKV6UVqZVZzI24DeoEaxdCNE+8Nvh/8gVMR+iW
7Eu1V9w1K2r57pgpyy5Y9fQvLlR4ZUyfDxUTWTBZL9PAo2S7s+nJKA+anVfL1qR9
ibWUUV49O91PGCzoqsqCB+oc+yvL8Oh5CwGL6Z8FMjTpUMRgs4OUBZAasruBdEHB
Z9iXRaWuiiT22GMTHaDbWTbaf2rS3MRDmt5psGfrNJgH+GNzbL3u1vSlXku4iuB1
3WlF+lkYxg17n8GXfxqL8ZqsFLR0oEQtE7D3jQNZLOth7HbEQbXvz1SL/MuOOtb+
h+Oko7L00W8jfnXlnUn51AMAph4wIiNdGC5xuycDzEQmEtVLS7rn4vmpnfiQ7U1c
qzHbn+ViF/c8bM6+lONmGfElUaqpZpGE2cdnmksFL6+7SKoJgd/UydBBEQiPmkXZ
9kAXfook9aEP1sQXNn2hfqQ3pwdXtyIkQZkCqlBBGVAZGxqyjSy6yUZtX7+HuFAc
ckO5jHSeyHGT6O5AqEn5kKoufdks2CZUJHTAk1It3E3gh7DHzjprJXjEerAzP2zg
jpdSuebDca3NzcitLvIkVKBDGtL3mqO1zmPP83n4Lem5X6YD6ozNtq3hOXwWAW7X
6ToI9cXU0d9z/+QsXAoEjNJzJxj69o7V1VDrDbseLy/1VMCbS8EV2JbesPTFIA3A
Ma6ZyRDlov0KpuYSZBuHESlmrLNGCuoYd7OEK6DcMxMtLn9YGFBSF3jFRn8rEPlA
NVa12WQjaq+gztJGCkSNcVNNnxxacTAsdoDqQBSqjWALXS85H/aogkD7z98kPDMI
Y5KcSdQhFSsBeVEgDXmmW8imtzD5ED3MHSIxIEfkCxLvKaAUHKigEXuFIqqAdfVQ
BVkFiLujq4pGuuT4JlUD2XF2QcAgwZNHovdPy8veil5rW0SlKO9iIbaJitwKw2bY
2/vcMO/kfSsp8ZkLHnjngo6bF2EKN+3xGD2AL8awwuyTYiZnBdaig4veCPPktTGp
xSgLBEAMeoPtTCuM9zD1rDN+xYQm3rmvV1+SamtqZNWm+9iOM43p2qTjfsc8DzJh
dRpug2R0RrjIHXDQQT41Ge2ZY9PHwRfGxB1+2izR1cYEQmsQNqGIrbn6dbAcdlxp
pQALY57ErXYJU3Z1od5OwCzhD2ms3086AecPJfw1t6P1oZKdANs3ZnKeosiD1b2W
7AiH9uWaaObCiqKsltlAIKfeWy6UWv/IOGp+ZMT4jw0z1Y5sQwmGrKlku2xoR+t+
lH2mdH410os0r3oFfi8sqCY4BL/XZ+SDoi6XX7iziY7wsxlMv9EH0WwaLYYzbmK/
ebxyO4lXGUK1+oG8tF6/OPEpQo52zGoZewtz4lhzZy0tPIwL8lIcENr+s8UihMLi
C9uMQanOeyIT4ufsSStsfOh+25JWHsWxjoOStBOxNEHijwn0d4VAzhnPVBy0FNoQ
0cX3qnnK2OBwgp2YVseS9K0oJwRh/vgI/GqniRcKHkZfm/AbKIPDWF7/bb01kS7m
n7mEykfrVeniP5/qgR3RO127YyRhguQ2EHSWvjh6zz8l3liN3+ZEzZxCDSJfufph
cAwhEANf5kexP5+XmuCnD6SC9ZrJUDUFL8xYE/g+22mzCbMYHho+hInC8kzRXrqQ
L2zRqkRP9kMQuX5L4g42vRBfPpCIH18SSj8b+6jPofeNamuyyMtlNBAYgY4M1Map
qYQleEBKjPZ6WRHcA2LOtn07nCU7qmmibgBu66D58rat5bJoL6btx4WPWasWGg9F
9ADg+MTCxxO6exVM3081eGSnM09JmKeXp7rX2VN+77k7rxg6TPYL2tMfpiSSobKP
9YG1LHlkVAAn1YhJSaa36lEVn7XItlnGGvFFuwneb7IhWrFt6EPd+g8pJ5+8mroX
mQbrkL0mDi63882wIIKQsDBEZDRCX2YdooYlGSgn2ZPU0BS9UYD0rI1y0WbKkO2M
+ZeInCgBtHYQoGBPEQQhdpPfVyngEY3fbFledCJBUN93FofK2oa1t91WAzQeLNTD
SuyzY1zFjByBFFWnUKQDAmXw7QgscUZ/8lDTa73OAGAzTtLBtA6GBq87EhpEz/XB
gcR1OIqkpaZNf27Hr99zmcyM5UKYnDDVZY+ZbwnqQ+yWG3zmSub20U8HgBlMtjgs
soqsxdEkDuxhtAb3gEV07DLLT/Pbu8W8RLOu7sLzVldLqc7Y6QW/ZK/FvVMAJITo
/Z7JJorH7KpWBaHY12YXuDJ+xb+UM1McCFEwmPz9/OdyAKuHZhwTwHv+QftA4kMK
tE80rRcRJrsrB9yrIll0jBb2UCnGNVo144aVD9D4RUy1G24e/GQNufaWBXNrL3xw
p+pZ9jQofbg4iP8tL+CSYUu3rnaGh07MG38oOzcDJX0oRFxWGMGBlvX8yp1rbmxJ
wgzuptSAS1dCvEBWGg3WvGDvnImPCaoJAQoWkogr+eeYejwhYRINChGYpSZ8yqP/
g+pYXyOi1WXvKShLZXL3AvgA+KyopZk2gIu2lL9RON/1u422X7EkL3tTn/0oQuMr
rE3KvJMIJWwL1vkrcOz2PrKJyS0FpdbFWdqj1XY/BD2iLyaQd7dRQNgRkWHr8rBM
vEG5DwCUtfd/7z3/Lk5lRLQJwEcLFWcNXQqDl2EHL7mDlh1bUwrpuA6+lwFk1RCX
yRExrEdf014dOJH7eRqj0aZ8PYvDQKFYvHFTkTf99eLJGzjBqL01XGv7vgPMYAvE
CiWjrOWTwpLXqVT2vWVSZDI7DUU795VyAwQBJGKITnSDOphoA32QS+5hjrgvIPOn
yifigPRsJ+gwpahsRCss9811axktiyUvPt5Nwru45vdN77Az9Ayw2nbGxWSJ8Aj+
W7AdN5XwSO7bV6Xe5OnFBlyPnQZp4pWTh/QrEGh3bW19S5ZgbHdJeszZp4Jq71Wp
ky9qQHsi7OsJB8/1kT29iVGKIDVN5O9AOx79swShbt1OnQj7gHhT4qBm+z/3wbtk
IrT5/bKNzw77v+KWyw+6ENXiDOWP89xwfHOSOMS3rQQu1RT8ZBY8OBVHMG1fs20n
vYxHu6kSXa7WmBizJlZpEwyl6ED/fZ1ge72IOESpdsmDv5VC+bsThym3fP18rJp9
lfmsbgFpLuvUDIdX1W9KypJfSdPt4jUeavu3w5UHPr+OCTeQe1FyXiDm74D9Yfw1
2JTmhHY7wGJvzJHJ8l+80GHaLT5/zK+bh3aNfgLfqW25QQFqz/eqxXHsv+dBmtvp
9mMP7clqludV6h3TlNcuv9yP5xZ9iW2S5gVgMQf1Z1hF1riexn2Y2/t1wJlvfNrG
RU9rkG+7u5Rs30WpXefzEwNC3JO6JB2pE1PjfAypvBoJ02X00M3KUf61Vuk8PAZD
mRX15V5TQ56qqelzVW3r4rngQHaG3V/R2yQai82hrEG5fOwK5PPnDRiWMWDkAoXi
qjV48uv5VTBG71NVUJ90LqfwV1kgLpiziogOENZ920VHRLv7dur4n+qo/kP5KOR/
DsY6/glzM+i4zhCMPby2Ied9OkvLBxvTYdCAhjToSmE/J7kPL7IfkYCOXmjfDt7+
HX2KYg4yfY3K267rqR77qin8SV3QyjQN4D8H6qvIwmB+JCHMJ1iUY3d2BzzoqnvR
+HwT/35xVZbS1jmaMmJx2d7Fyygf/Ymq9+okiU7YHHEy2QsmuQpfr0hLdcS3mWm+
oAeimB/MoOfr+GwpZqhqoNPoXv1ZfzbF7lqv3GI84QBNmFOMBPNHlilBkdg9x4g1
rg17XhdPv64MRdJUF7NC8JHxcQwWODXJ4c3YLxGHXeiqHDBys7tTM52G2OkmvAwI
KUdWOoIzQZMC+FUzVlQVNSOzdldsi6yrFPZbLcYLG6TIYb0snM4sOlTsQICnKWXl
yXhjrw21nAyr34+3uwkZVUp00iRExT5N2KQxBQCkl09Id++ECGITjWn51APtBx2Y
UCH5pvJVNo1qc44ID1pqLNfIwdimrB2HYf48jWqwwkZW6hDdMI+pdaer9GZwng/y
gW6VO4pXvtkxGkQEYf0Ge3rlsAt+w+vFQ4n73c14G6A4RMfuS8+iGKg//lNop+LH
Bh70wR3D/u3zRHK/bX/y1Zk0LAQ4iUP7Pe3wlwv13Ta2mGo+aB5ZF9dEcrBFQJ9c
uHVwXJzw+4nQttHWfRnqhwbFWE7TvFAMH2E4ZGt9OyLPmMjEYy4/SagJ1qYHfMO+
Ha1QGUV0Y5YCkKmuUiHLhDKWp14XOrGpLNB8eiJxwGVKJ9fgr/HB4RrmmsA9xCm9
TUMfQ/w2I5LYWyvFk7lFaQZvwjuL0pFyHWw+gjxqI7o71ANHKugZXwf5rb030klH
Se2SYM0DhtIDSlSWnNGPzCSRnI1rqGP4ijY6qFSzWh4Pf3pgujY/6rrsyMgYaJAQ
XKzJVAK1J2ZgWsTonWauOjwtohwkZ++Xm3L/cZBKKuZFJQIN0j0Gx4E/d3ZXttYY
7TuYCxpM28JKQDj1uJs07j5DiSIfi7YsLA9ISnL36APMEudgrZ5AurkyntB+3kKq
NtjvTx8Sfn3XtoinwsgQuTgYuBXjCj6GxzDxgM5euIeHmRbtx4MKzyzhj87Zvuo0
FPnqy1vUaTewddzNFroCZC6MddNtsovXeGy/bb8J9+cy5HcHHSCFTExw7wUT76kv
L2OcmYnr+TQ2xhi4G9Dg+fNNTboPExAMcX7ffGxPs7zBuLYS43PDDFPU1TMHl5Eo
ErlWHAdDZmvhhFTo/FkKz1JjFYtJVtOp4M8iu4trYPMeU04v7IrBr7Y/+e1deN9X
W7cSKuMRePXhpx+QscF5PKjKOKSF2dqxRNCaaLjSruW7t43/btc3ozmGU1c9u+Om
7zkHcxPKceGaELjPwRrzmBtgiY3yuFiANdu4JCg7qUHQtD7VGixShxiimf2xHApf
bAC2pVun4XWsPU97SxVhLJ7+R4ACCxd8NOd4F7GqgbYWocRus1lZdHd9kmw4+Khb
+sAqig/9ndSYga6xBHCfE1mmT2YIxWmE6sSYUS8MmR0xMY3vK4G1BN8Rs3gsL7SM
UkRjFaKbZWxn5QAPOF2uaRjRTr3mzFteuVMZZMc8wK9yiBpzxn7wUTHNPkz3WSkz
HD45DbbOqUavwxM3VBmBnkgd8rK0vyLBS8s4H4yZNbXl2Ooscj+XexJ+PbQO0zTW
vlqIeuk+Y1/7RzSVTHeK5x0ZR4oP6UbYxF49pxI5rrf88Y1Ze+JcBTsJN0AhGdKx
zHbSKYUAwrWqsAWswsYovLIC2JwbDiXCivMjI9+CrESQA+RnjB/hLm3PfUJ5vwwc
Vt2z/DnX7hPYziZ3BjK8cJy002PK/HlEu1Tg6BcbXoI8vWG994qibamV2PC5OE9L
Dw054wuNFB2qjRwfoIWarmdi+OKAXJnuez+vgqs5Qwiqpi5QHutl4zbRTLNO2jpz
KzMsu9at1rf/p/sAIFL4SN6Dt9tkio1CR1KmU93uCwSI2KCLLrdgrJwaU6Wc5RKL
9F8pCYkKvdWOoPVLkC+5n0+2RMfpIkGcuBoUQ4qMPXo38dgOZp/B7qNYw2MR6eX1
A0we33wLQG6fUUwCdjqYRle/01hFI6ZMTwm+6tQllH+snVN1yNA1qX0tmR8nzDIE
1nXDPvr+tXYJkkCgmGK1Ce0vKfQWGq68fSQxduefkf3FqeGv3+7KykuBd67Jz5W3
srCWH4p2kDIUyFaHOmBhP+MQFVukA5C6Uflq1xLcDNPmXyTHq/jKQnsMTid4EJrn
tbG3i1JkbU+POnwHbWg/Z4VyPqvzF57ZsiPHBT+ahzj0sIb/NnOPsoQmnoOW/fWS
dfY3Re+ql4kc7YRM1IVS04JE24Ayw+fWSmumJTBlG0774jMhkPSiETujNF74k2A4
OllITpHpbGv8hfNsqEXUE0QJ1P41Jf+d833W6g2bKEqHGmJOvMDB0PgfGIdCTLyP
5+Q4mQFQU99jAXjDG9F7irsB+mdlsfuMCDxPhLDh7FKteIYMuHAm4L58/F8smcpS
TG4yh0uj3vk/8RL9TvyVaqC/WpcNFIIhcde+hQTCvQoHIMfzZig1lyS2O9DzihQP
K5EGsPhM12uNMym13pN0qxDKbEO83uAKiNBnWwd2lMHr55dnDA6/CMOdC7ZKN8RO
nN3nFLEP40HbW9oT3MRGSI/a/wuTU5EyRMGnyG3WbmEBZP95UPhS0cMwa3OR/d3A
h6aD4RAJPPfUpyvPhVbNr2tIi0lrp3RVCYTEHxsohAsTuLT8ppzX3mIke+r4cHlN
r5wwIavRsUvFePpYwo5BUdSaczm2I57L130Rx9Hd3ujYz52DpeSWkk9P9/NI+rdW
YGqBozkN38bAOSOTl+E8Okx4ssFgxMVkiFW9ko2CBmsng7TO5clM5uHCpqRsY48j
E1mprbWCyR7TAK79AlCPUMiI6GRNcICxS0QFJu/gYI9ElO3d6/cnjoSbtSXt3h+g
IIwOy+j/h0c7e8m/zEf3mCpE43+etvY2Qr+cmF1rNhGCO++y2ZFcwwsDnBmL03ap
aoGShLMWFXUjaDz00MUHdYiCWUzzrsJZ0undBJjtO70hb1mMAel7GnPIQRLVQmTB
Dn70omDc56hMKmZNy60LqXGbGDW5L2Yf+TxMKuxbcokcs58mJpdQG8NIMsJeQhkO
k1ct6k4L5qBYNeUSwxQuP9Txh+aDHy5m4gXfMGVISQlvlPk7ShC3iVw+C/BO/VhQ
CQyYwKcugWz0ZFY3BmU0/4wb0yovUnOu9QkabkTUIXtu3KND2iptqzHdJZqMIe6M
3KNBiUw0skM91FqToEqQ2xETuWr+LOi+NPPw0xSg5Lbh4Hr/fJEnsU92gL8Pixw5
QRnuS7ivAo25SE4WMx/0gJQMlJvQ0Jd9ijmoNpPv6EbX1tas9/shPIUdmoUoAiDv
GcrNG9ueGP2x45/0Mou4tXmVlFb/RUTRjkWPP1pIxXttsl8u/JI4/x+/hXGCMQQl
/SiEaJqaTmj9v4VlpP7y9QRJFu9qsG2fTzs8nT5agWQh/BDdwCFVkGEvQ4bzMw1/
uP+0w5jL8njwFxt4js0Rb/nOSWLnR4lw6KjYCJsdaMVsmtBIyBTO0rvKjc22SK1N
Nld6EIXTiM6ZyRMvukhjg7eEK2nHHI26Oy2iK0qv5nXnnFKEEoXkSwhVP15zKDb2
Y2vXDtv982qFM1Pq4SXsEnofzfGTr7D26sf4lGaFmVndftPXlWdh1eFpjW1rXVKM
rNc9cCRaMimGYP2H4Pdhtypo1TgvxJHKWOdINy4+eMyDiAgNzndfsc1QuQM47d+S
nuP5tdHl9jds99DcV1BpJC+lgp4N1M6+kKXd+6BqbpE/EAFKbwiGxN9ZWDmi5+HL
39p/SCMPzSpVS99Dko+kkGfE8/6v2mojVwDDgRoFLAxf9GLoz8tUdt5aR0MO+7b1
WiG/2Y9rM1B1htyQgeIWclftKtXzMZu84/E+sp8jxj4Zc3PTFuyc3BJ6qoTjvJna
i+8sF6jTiGhPsOaDIlxXh6jDYi59L+d1m14RlQIaKaYk8dMlpAtETbQiUMlCfddT
kq7y6bnHqlDAP4+PeXKQuq82mCyr2RdT/63yZCgdtRGHDziZW6QOZe6VEVcD/NhC
WPNEygftBma/VTOmFB1c9hhaWClxiqQgz9D9TzLPew6wD1ZdGKZU88uWxo/sq0tg
X+kkO8dWxU9jWutEV/unme8UrfItcHyzesGJJSl5WITYE7yr5nencIsJo2N+uc8l
Cw/LdHGJLC0x6pRZgg2qqUQfooNEdQrvDnUGnC4szGeQZo09++MmA7kPN0PGNFwg
LMGbwZxy/c/TnP+CDIGui+IBB+ecTgSDB9bNV7NVdqhr2+tfxANZuFFyPRTc0TCb
GIueeN5937X00e4omzHISUk+TwP9+rHx969C+vtCo7K8pdvGSojgcRYWg7bTGXa7
TlB2FEPTHhE8mt502egx0ZtwwMVhwGQVFntuBpR+NU/N0hQ1yKBXTHDXayM45Bfr
apkBKlKj5PlHfQBoafzqGH2SzMUwjhDHJ8xU9j6pn424y57kJrL5DV9roMpWSgei
yv8Y6swWAnObRKPzmpkPZ5HhFZMn+c5MTauxj+rWOir0oNHrY/s8yKCjJ8Ee7kdx
9ODfmDpL2iGchwGAgzgnJ5DIXR6dc7JqZueXB7ymY3KwW2mDkn89bdyRQS1wSuJn
+CAFriCdWc+k6ABDgenREgMSutGaCZBlTnrxkwl84AW2hFicXTwST5Zxro0PrMyJ
KiVNlzm0P5FLnyfjzzrORAwPbmDjNi0kC6OySlqhJpOd5E0YiydGWjxHP2eTW2Ik
xuy5J/n5MNTHZcjehnXm2MNYTKR/ICF7YfvKsI/76W1Aav0xpBtS+OilhslEbCVW
z3yLcXOV/qqeT+98r6WFCgSpn8MaMQ0K5Bzsk+tMufR57/EOuRmQXrKjS8q+5bgr
ow5GX+wUmVHIaNa9AU/VqGSzDFV2sBOqw6EUOxZGIaiwRLBLgTFvPSTQsDy9Rfp2
7pOI58E2VsWypSlIli1HvNr82hE1eI4eyShar8SMJkN/BDD0z6F5n6nYiIoWeZHu
Lt7uiKfE9+pqC2QqwbNSfdLu4pV0nIGhjuMR1BWTdwRjwUu49W0Bocldsjwumfp/
fzP5XPL2tHT1WHYqRbeuRL97g7iyEuXwg+aqJC/PGZmaYV7BU8A785DPS2DYi+s4
eOHbxQyUqCfrzY4VYTGMqVKxh/6Cb3vhq8oxbGx/yDZwM61WDDO9+iTWgklnqQ+/
xoQIqSCvHmVhWelUm8bITSkbvWU2nz2cbgL7/9YzkWd8jWHodstKgXk6E1O56SmF
5+nKak0buXhYGdLfeQRKndQlL9nGfbetUxVrY5bHWBHx/FKfhLO9PwYFa5NZqAHf
eCq+WB3ezECopwKOmsQNt/hhDklPbniCh66mrWOI8s9Q5w5iwGikaKG1KeF/jC5f
OWN0YGsN7j6rV598tGwVeC0dLR6fzIK2lnCyx67e4MHXsehKclceb862evEGbjrx
2eM7LG/Mmk2lAhPQ6FKQViLUv4W5ZXBtLf6BoIVphOCoIjWNrPvtnBqrJCah2oCd
d19LSG9D3rKtMvoRbChLligiVL1n+N7e+wIoAzhO/j/iJluF/ztudRVFALA4Y7Md
MVnCwdLHqvskapJArTVRoK6EkTKT6gzojtCP0O6F7TgTdYwhofy3/8rqU3vEaMS3
0ZRCG3T7pAd0Xy0+hi4JdoWK08j6+bOUCnwzXe5Q/1AbPMtSvoBjJYb3rvJ5kDnC
UIc1owdC0BsdCldwMYc7xrSMKx9BsLwJuKd6qtoweUxGnly+YTPND7ch74lwNDam
G+RoCcfC39siyVX182XGaESmxmOHu0tIXLy/8anCx3zWZZGK4V1KBsw+AurlAPVr
jmFOO4g7k2f2fW97kL9TbHsxICVlr57DYxAeMIO8cpl88mUEdCwWPbo5hpDGPXFS
iMSX2TX2fEQljORMJW1mcyFwydGC1emp93+91Hqp582KMJ9dR9gNlmm5HwwmEFX4
Hjwynxe9jxJR6fWkqkR0IzAhx9UEe5cWPsItaDzOYOUnhcZKnENiavnsqurQxt6o
iOIKisMiyE08BCcGQfY6/0RsaSfSoGmzK5bU0cPt+P+ibtyS1ANbmKhljNgZ8Hch
DNjT0nDzamKb3J4pwK+E846Yvy2fCh4kCr7zmrsLyJnX2oUbOXlXbjjO6Jovgz5e
uXiydARNE9RtVElWfwRgLBAFumhLW5cOZ6BwkyYpp5rASTzH9k5ym9KIGoKx2Nx0
Mx+UzjK6mEiupNvNPDKTeXhCW4AxItHFMmk3n9zO5tuWjONVS32vHgM77vzuAMrm
zKZCIW485L284ENk7hQanMzqIa/+4/ucatA9XyDJ6GgliQ0+ry+p2N+A7o1dnkqS
PNNS+v9LPNc9jKWZY7cHBusj0YnPUk1/J1yn6SRnDaEDP+plLMG2dYZMWojogIHr
kWJ9HKnkW1IApht2C59xRj3fLWnC5z8KnhVfPvja9HE6+/GlZmtYAzizkxho3M8H
rIOQj1ieV1YZIDB/bj1bVF/+zYNPRQ3U8wE25bBm0VD6PCJW4qXL1N12T2zdmgcf
BXmg9XGUkg5SYRs14LrI77bzX8QtG30vNG1Gw9qYvPnrsJO2sTc8OlrmNaMFIZPB
HfO0djehorJmL1bWoGotyC2NZk/uFvbdb/Fp6VRoiID4YDkl30NgHbGtKHOIAEK7
1f1XDsQ37kpGEeoo0hy2mPzWrl6t7nkrXnDI4KGZEZq4GL6BIax+oshcVQWXK12O
T1qrxvNuoIlJyIGJ0TdIIZuMcj2wAbM4X+U5mV630ca/nEXf0+00jC+AYgWSl/+A
AASxZDSyrLIWI6Kip99/DPXe+d4a+mDU8tRsRnLSAo80zujMasnfrLMN93nyHmT9
9URTIqYe9aFqQzdg+ahcFieRYCO2HT5kac99UP9j04M/FDYLCIUlrMi7FvkiSSIh
i1R3sm9qfceEe7wbi8J1zekHxk1h2IZ+F6DA3ydSgwYacdMyOyQ3aO4U23WJu5oE
IX71gxC4DO/oBqXgKmRy5VeiYLK4PYQAvR6vcowiUpHcgntkWU33PnGmlRxZtfUz
CRpK8ddP9BvCVNTcilyqIuysWn+gewB/ivpxWS7iiEOuFuNZo5m24PUyTVMjMf5Z
nLHvuEMRkIVCXWr8/bT64jssNdPzUjV3eXqStr1mVunfI7XxuwflP9tqPnnPr5o8
yXrhVCwHaf5wt+mydBaOF92/0EpBOAofTF+RVD0i3gaRh4vcLFB9aWdHL8GXs/U8
ypytHBYsxGrvx2yE69ul07CE+VHR1rmOsyfuquSJwlbA822PQza62F4/UoHabCPb
DfnnnYUG7EyYLaPkw1vcPijLy8Jck1xUhf0qLBGH0tMgV42BmHwxjxMXcCzyh8x5
b+15UG8n6OxPFw30xFdO8gsDrcxLbGzk7bKkAn5N8vc6syd/g0HJPLEiDDaawTQh
1u/aXsUQ+JYpeFOJLx9VaVNCF5w7OelwidR3Dm+tzJAQXGSbciUiGOtsq8YBb7t/
8l2x099VKeEpdu5wrUrdmj4fKAVbGbVxPHZioiNnTLVSEYN0bW2uu09FvI3ugz4L
20gu+xwFZdLCqRLR51EiZnqPIUUyqucNEseo3da8btmRiiXXScUh/g38B2mwVGyE
U2pszezkcI8VuEFkOyeYtLd3mkEG+Z2UiQnE7jSgzg7bbJyf/bG1mrcWFIdiPemD
VKT6sTQHWwx1IEa8gbDwtVfkgk8NzjX9crkZwBbY+v1WP/LN+qp0b8UYNcJtTc2P
lzOYCU7SNqqUBpHO39qzX3ViU9pC5FZmBzqW9ObzUX2mVxkOdO8wRg84rdKX/dpO
63k6zk8ka3pRjTJR7ubtoQxjj230HcvNhEU2IwmiZW20VpjdaKIV9nKHTov4js27
YgCgO7IMPd287C4SaUtzmzeWXdBSfNfGBblpQidtffQY426lF5bgYExSr5fq4q9j
jLsI4yR9Q6/yimX4Q8RSS2ep4gn6FBMZ1PF1C1xSBLxWZH1MS4TN44xDT7Lkp1BV
bPgbzli1nvchqUm8FhbkpAl0SpwzCKFxT0/w9Qb4pjcE4f6pZEyCeU3wT+HZXqwN
nQZBPRwJ0fX43H0LGNo9xpeTXOYQwrYoxcqkfTzT2PXoWlc3qYrEWp45xmvkjdEe
t7khF7+9Q5Jv39QeJLr3D9SuBrx2HFNW8A7MK3iCM16zdLvBLn+FADo4MbPz0zh2
fTGn/EEIfvoYQfTiJayZC+A8Nxwrr5W/TDCLMRHYzAx/Z36oUgmh0EieRJkQJ0gj
I8msIc1CSByuvDY7eG66S8bZ2mCvaRNwQLu76ZWfosnyFdPyeIeYC+UPupbMf5Yd
Ad3ZEgKMDXsKDI1s3HQscfiINoHKcCNrnNoc4a+NQpm8hi90LX8uYhVjDkugiGcs
lVbh3MkamMw+e6hkaREpkhacdgtakSxproh3C7IXTZ1JHYxywMpNE9QHISFjRv/e
++20UVTrISb/H83DcB0wka+G9OB3U+E1gXb92VGfGD/RTidnRChWc1oSZVwV2ec3
cJF+Eijm62roXJMjafd56+tb5PGYYtMmAOQCLfx6apAMJAOfjPFkjOZ+wyYSdOE+
5WOhpVbBTNNg2J+woAScIqOir7cfCGubPs2eUhiDLV2UYuFUWsyBvAFmq/wU4c6q
Qsbyt7WXIxZNWOLhw1NVrAhE8WF0Voj1TnmnM647diUsd7lH6g+3a2xVmXQaErg/
2eBgFycDbssqcJyZelP4zvvu20WMvPvGzcsN8kzo1ffP7a9eeHAI46P4p0hSJT3u
PS8yKn8cd+zoarFeeT2/+IydBbTtreszqFUWUD/FnD2hg3RZOruwGzCt0HRgBxPz
WZPck23i4S1e0s9j177NUPtVxxsTv9bfmUvsVLAbGxFi9xHo8iqMTTBtkhErHVxM
dlAZPrMITjSV6KjUxEvnDOx3ZSD74/WHcEtHkMkW0onrjyeCfXCX9iuBIy6RtFvm
RbBElb16BZ0iTRQL0kWxAVG9Pmhmr8ylttG/uRG52+b4VGJjfB08KnnXJA0uY5x3
K1tWN1cc7hW8QCYVEDB/14VcYHN7+/6kaFYXUprI+QjhNuK2ZIJbRNGVvqmB8i8J
018oaLlB7C+3x58uxr/7VqkDn2imRz201sqckEFrmUARNj8SAEboewRMXmSVgQAy
+MOOqIOewSYw45Ouo6f2oDB8r4CnHbTsqeXPXvxLH9wprte84GYPLffMlE9ZPisD
Hx9XfyBwu7nDz7kgkoEMYw2+HsB4zuX7OjIxWrFAOliLFNIMJz1ypI62HGxuyV2c
R7Gqh7us7VL4MTuf4QYZJnGd+ZscGO28SALWIQfXGb/un8NxLKfPdSwlnI0Pitrz
vTxAiKBOqKCRiVtDGyO31sqeIdbiq4CrC2vt1VLZZDAoCu/r9ghE1RPICUrmI1N3
/2ajyGDxwxcuy0ZX1fGWABIn/HT8jA9+M/Qjmcn9WsqO+iiu1NNN6b7TLDwbG0yO
AqzqZcR205bsnPKJJeBgDgc9jrZIF8yG9q5VYAx83PYifBujiAIW3b+fNOrTGqnE
8bWpA5kgM7A0C2O1VjpIikJyegRDZtpMgYwqzni7Fi435ROvcLUZ+tz8rkwtK4bD
wWlNe5osHkzz1e3CTK/x8C2LfiFaflukVEF0SxwUv0wOtQbPJVavPh0TxnL06rQ6
aAUvCMleKLV3mFU1X21z17RwJsIGODNlrKaJYidpCnjTaHE3drw5m/7g/44S4R1d
DbPw9xbuKbi/YvNAUyA6nuh+wnrA+fV/4/ariaIur6NyeZhfNH5pCQ61v1pwxwWt
YI88v0m01WTuc28200W8l0wD1bGP0Ltr0/oSeM8W6M26Jdl5LurE5y+QFLUydlcO
FlwzCLoyQkPu7YPP5WELUDmmoMiMMPV/VWPyc811JnGmcbkvR/r/YRnNTJJqU28k
bgXnU7OgfokrbpDC8WcFZhZ6O6UHxOMDkqC7/afEYAcjpD/87IHYI/NMaRM9hvyF
skRgWamqht9UMkEGYuE1I2AHI/jIThmwQprtTVYqI74l/wTfEBiXYUIc7fsUPpfo
2HRbKEbiQThdJqfILtDwz/eMrqeXKH4pLBm3T36JmerRhA9a1PcGczZv15/qbYgp
Z1TT3CvFxl1KsY9oU7U2IlhJhfWd6YAEEAdHBZvTq4tGn6ibMN/9yuJ0VBYXSP5V
ErW2p1oiGRRIKgLZQphN9ik2HymhZ/jmZSMR/OVubvYB5Tu7czFtOu93DU9tfE+P
9+aTyNQCJYzyJV5mV4wwmiH8Mjlbhv410fqJcEVpL14DwlpXkzW8ArfwNovT/dvh
rRds8wicuqTAxmD+n69muyA+W0AjGZBnsbq+5b3FQLE2WLw5k7yorLdq30fGx/bM
PHGamZUi2LplC3ihl3gOsOxFounivVyUlYTiWnCTH+3ZFJJxmbqkaTew2cdZieS/
C/Kic+E8YhQsOA5mZeODH5S2yjheigM1WsDtnOMpjDta0j+/Hix8aPpF8H3PXbJX
G6U0QqpZsk6dHS8F5bQP/1DsLm/LbBrENOw8s9rf5anykxbndokKkU6mLx1A1Kd7
dzYZPFGECu7QwCNfEC0ypEe/NrFj5NSLmoeq4OKdeE23RsQ/TTf+vU5+DICeZNoZ
PVosibtismTqZkvFCOuvcq3JfmDz61lJcjQsdPggSllkESCP/4dlF/ghvq8OdgZL
sbEGOrHykMkDtd0mXc5aWFeOj/c8TFBZ53SmcQ4It6IKvV2AiTeJMkHNqFux71V9
4hIwIXkfI/q2Hk/ielPIrfL/rVqMD3VJJlpAOFfvbOWLjzOot3pr5mykprqQ0ScF
QjJKkSQgJfDbZH0Esp1g0wZs6hHg9WVaou5d/+esgWZ5UR4qD4/memgbHsc9vIow
ye+SZ2739oftp05geE/NbDMiISklPfyr0h3qIEe3Cun8ZDL6B4jI3isfeNr9o5JZ
RY/hA1iOy5tGdZ7GWmkodOZNvC4VGpXjOVB+8DQHe1bUiTFgi9yN2ksAhKWfGYTR
4q26GDk3JNlGfdfxjNaV/oQY+pz4p2sAk++neThKQqMltonuZSTd2PcDuP+kFhjs
900fV+gdDkpupli9ExABZ4wk2K4om+c0wKjJdGcsk68rHEH0Ej7xqkc+f0V0OCBi
vyDLb+H2RLuNvETObYs04xQHRMoBXsB4nzpLkNhYtr5TBxg2f/BJ1HaNyGNPpXgX
4LLDYV8rkbl3rh9kXUdZTUtvtyYro8n4byR6+5D/eaaQ9G3NDgld3FaSmarR7hit
pb0fJnEaBdQ7Wa+kDhtnqSTQ8xSD7yTF3OsbGt5SqMUdpc8YyQyDWwgP7QAqS5TC
6A9mcacKGi4c5pF029OIQnNG/HEuI2a3JaIbR/3El+IpUPWnVg+FHtT8DmqyoIi0
a6ZKcQ7tzXArMM8X/Ov0Lcw0+nEamquEVrs7XO4/D901WuPQ0oQ+pi1SIndeNGrw
Jy6yFq4RPcLYl1ggn9ffgofwbWxNcgBgPzJicnlF61/JJvo+8E7M4DkVFhiMN/Up
Bl7SEUuI7yizq2Nc8w3WYsBxrr+iGxzTRY0Suz3mlhr03UoF2lKZNa12G8OEZTY3
z/SKfOUc7WiO24MA0UaaNmyMcx0bgzt2E8pZEQo64GrY+NSjdGWkqZyE7Cd4iDM8
hhnJpKd0rWY6vzCDnu2ru1gsqFVENYrJGEYf/wlCpTBzrul6rGsiQxsfnSLU4G1Q
JmyJzTWBPNJEF80by2SW55pE35/SbPolYP0FXOQdfhg6yIlzom9+eEGoisvT0wqz
SyTlSRP2ri3rg3S/eubsSlrdJJoFDh3iD4PnzU8fWikbZTfTQBfuqDoofDTGG1WX
/pBBNAwjjwr6GuSnpgDX35EgtuxPYAwHAy3EHlb3kOD8YK8UNjV1ZUj4kTq7F5JN
WhptosXH3rxW8Zh2e552JLcVwKCzDsSjaNCwp29lxHogbOcneW5zrk4/q01YYt/c
aCbvmOHu4qi8S1X3kQK8ZBOAovpBtRnjI026Q74BA6Y+Gkt81I8z9e8tvDJ8EJbz
i+P5DlW/R/a/mTE/QK+UGXR2zSRT6cTxsMklv2cw3XP//yfDP98pHWChx1CfQAIT
luTyHV6tmu4CtyOgVsA0tVqhwLZ9/kUC1OpkR1/oBTAP4UmcL0NsW15b/EfW/USh
9NFyfX57BSBGg/toJtxn8FNrJJt7qIZgGVUfRLotQ+B7FfnS+eNSrE9+MrbVHT4M
OzC8CUtYp6lzvsW/2Xm9NWhze48AXmpUzvdByhx2CPH+xWSIRTYEkXpTDwPxNuAH
mx9umrYB06O5+NJsynRmOjaaPb7LgjfUsQwrVDcHUc/e7feBWlPHheV84Os8hRDc
UI8l+ZzgPvK62F1LOoPO8jYkR4n+oaH6HomWIWWOR3p8ggb7VWMiUzrSRtn8Kag4
jGg8moTnJJON+gg/cNQN8gnCMKirN0QsazJP2mmzVoUSP3ZCjA/kBAMwDehRykHl
T8+4onOAqLkILSp0BNKYP0mgRRI9VWuDau71Jbe+qffmYuuj09SZWxNH6BnsMeeX
Jb77gAM5Qioq13I+w+fFkrdcSb54rswdlaDRINbOs8ZE7j9NjZXYGz2rnnaS2O9t
j1qlz/proucwkRWwu4apgLBOS+jLLxUeDOZV6B1Am92DQkmAY/A71T0WlzQSiH+7
iRbgBKy4GoMyOXY0PxS8Lx/Pa29DgUr91QhiC7IK3x/HyuUgkX80Besc+U036L5X
gkDF4nnqsiqsS3gcAeAOjkSALfeWsMzUcLj0e1YAFiHXkH6v14FihM/Lhsgyl9rF
RGuXpkveCIEITm/M3NTC3ZT8dDtNae7ATZpfGQnO4oZB5OekMZUWmHIm+ptWypKX
iSx3tFTKkWIsuTXBLTloxDwRJtnN+lTGvg2ZJ3mIDwLeCZitIN35/dN2GlirB7Bb
J++yDJwyT13E5oDPeyFdN0KdKXyhIE9d+2bDctGSh7PKKsLd9p4+eva4mKRRLGyD
TKhlRfGMQwDA+dbaOWyZyYw3pCrmxEAiXW9TlSY1BP9gqv+zrFe2YYTfene61VoN
0KUwwwh9aqeU7W6r30FcLYUp4wECF6+8N+L8mijKSCeNt4v7yla5qjXCBn1tU/II
kuoKqwFxyrCfG03rz/4d0u4P6iTSz1YEkOY5JVKTc9shEGcNVb/gOvhp/ve3hnpq
xQ5V5pu8HNh5IfTxQYyOyNYh4Ip2n/K9a+NfjazPeWyoVCrjOuBSCunEYvjZeUkH
e4sQ4WHj6sxE9Q0pTd54fUl+c6ExEJqd7DI/iVFtFtc2FSLMpJH6YwOZ+VsyTuvk
qliDIPqZxZ545a6VA/UoRV6P8dhMXLfgYSt9hui2cQX68oKTKrsPCgNenpRYXkNQ
N69TRRH3e8KWZImhSfkziJzVhBtA1AoST6y1V1o8ooaZYvUhEEmSjCwDFgnbe1Wa
SeiPfQJZu+jIBPYQlrDZpLa+vtZiyA3TvwQORTSSZwB9Ffa+wjMY2Qm+3p6ocGca
wtjg0AwhzXFxRNzhfdIr6Y+qzjTT24DKLT17wWipBRLjTxCnDDu4/2m2EHchjARg
dOjflGT4btKOAtVMusnI58gOwUtzZuisaABjXiGQTxLiEdsRa3Oc+IUrOnik+5zU
61pVt3VyoJg8foiK2TWtxOkEf/oEOUn/1tsr+hF5VLvxXZXE/A6+LAKvh3PMf6ki
CR7OT6eswlGdzAwcTd8DIVDshoFvlewJzl2P5JpEEdXxTIYt0yMS68RBbqzwQNNl
NYjFJDdSaHEx8LkeoKVzkCiw9NO5q7CvTgO6Z7BVQug9u8/ffFU2fYDUk3q6JMvy
sb2nOi8/ADulnku8yx/Gsd5GF8hrb6pU81p4+LZbMcevmx4ocEadm9rTVegWooIG
4+rBLR6QQRARv6nBUvV2ogGBe03eYOixXq4sFKzJIEDRMhAy2VYcJDlO/LYy2c4O
ppEybMf4hdEbOrIfrs0tNO7bwid8K/LC5PPvZ8obrM0in4QRdgCMYq1hKSCBLzON
X1oLJA6mZTH9P0Rpq0IYb6b3e+EWFRIdq3xioRIpnh2Hdz13U4LX3AMjwXCFK9aA
8Qb+yAUFNhmNYb4eDHQGHEWQ7YaepufhfZBPBtHtld5ghcNVZSxEt+Ovt+TaM585
zMPgBz7r/KuRFazWhopOJ1HrtLfEgepxU/MvTtEaIxoUN06THyQrQ+E2IG69uBDA
zm59rOKsNdKuRQWYWwld2PyJHP/3e0+kU6/SLD6BxmVuSsahwPqCq8wF9En7v4sJ
fEWhn+/km5GzYSEcBJ93z0oaspB/hYPq15K0SKzE+NhTmKPr96jzNNr7AJSqDwfu
uOVovwIoJK2dSKcLJ7gDXD7ZAhOGyDCVgGz3w8Dv+OQHiBf8imwHvN+5Y78SHSY6
e7mABAbr8sCHuozaJV932F9RXK9NgN04hCKdIITqZ9wm4x7E2H123iuK/DBi4Qeu
ub1JzG8pIs+qYYZc9gGHQslT1v5vSlfq72V4x37K6HZUwb6OqCrgqI4s4tJ9o9jE
qRFEq9fqjQegDAw6GBWWVaq+k/K9lNXDV/3HzUSyPsYPWi+FFladmiAXB5fHhZR3
E8fELShpVZVjCYi0uO/+h0h0SCCLQ6HU5aphPQrwUHCee3vCaE8hrRTd1Kg4fWEp
2+oqKf1wdgpwUXwZk6DB965owgLDUQs7hwqrOoXOi5smCp07KN4CisS7M54dRCRi
VZOHWVxcm3sYZt4hjdHnC9h+BBg+VJWu2IpuwFvGh33bD/IeTVy5HV7KPheXjxfe
nz6GWKqHUZ5SuMfsxlANJVfjg1qyC25D2u7SAX2r0Ww+v3ZcU+tZ6JrhCdz+Zw7R
qb6qxKrYSjKreebJEXey52zDCVx/1hBdQB6PYx5Drsu4e+7f8Ok4/lWupL8jlBlD
E+1EyqSmLZxP93LbV4sWPm4OeZaNEzJmhL6v7p4Y3ZXLwePrDHHUXwel31gZima6
D58RMjZlzZrZVUsLHfhIa8mqAflgm+YxlBtB7m7yjcYzVdOJ0xD/4bqdyvUXHE0r
EWrqjjeodRCBVkcU7zjEOuRWrgq4dKjG2yUlDAMOossw64Fxaxk4yX4LGYfqBfz6
Fnx25X29JMIt89uPODUoc1LZfJPkBQWkWgOTzU/mCW9ElTELOmkgR8pU0saprizz
zLuqRT+aiWZJOhEnruALZcc3BaTwnUud4KnBSd7IPUBDpeYmskuvjbT4M1iKivXZ
36wk7XSG+pDTKZPl062MsB5efK/8RQmuBzgRqZj24ToKWTe6wNGsijOW6VS3CkNW
YpglZ0yB2Xy35euooQPQvxqX7QOajbrVH8fhq+I0wB56y7Tqnl3D5CsoviEfR0X3
C0l7iIM1FIxQ2IIakA8TIGNcl3U0J2v6Z8hjFIds5l97DwX6bnQnM4QnjFuAaPfi
xBy6cr+3P9gbVZyTWySS16OVmi4zBQvbxd2NTm04fGcXvJI8O5K5ZApJfVud8bVn
e45gUZir1W3shUt+JqslwYDk8gpmi4cvks5vG5OViU8fFHYTKq+Ao2/o7xph/2r1
LthXJqQdA2B4raU0QzJAwgH0j97b5ZGJN0iOhzTbFU8OKtYV/kTY7YasQ1HHxVr1
ppLP7zpO8Q2X6nG7YSKcS9J5CXU1Ct2gVZzdRdG8DINml4Z1iAenlUoLCZQ9XXm9
BnZFWJMUroKBRv05kkFbXKR+SP+eECuK3k0MPzbHJk3EIzW6PeuIWoUpZ7iEF7+x
zCLF0m62gDAzd+cAS02OVOz376h5/9iQEcnkl/g6JtPQhzqjELHcsU3VAK7xRRRf
DNLf+hvC1YAiQz6OGCMwlhqfZbCW5SQUXv14VN//CgcxJgA7jEWFt3yPYmk8c1Oy
HIL0Qd72yEI2Z7gE1n0u8bMuc0nSUgTS8rkaPKHqvu1MtYIIycK9JGITnv8GqwB0
pxJefXimzM3sscKU4lZEtyN9RsVyJJkXW7xpGRJjqi4J7bsW1S+eP5RCiIHo/rpB
AFUopzQQwLntIOA1WwvNImTbQBhsDRQUNLUV6X4IaA7OPwzRMGIuzVeBqJWaWJOv
WCOLKIRvR8U9OPcpZgkesxvwQKRPP+ClO+DhnbE9GyT/bsfaFkUdv3XrV8IGKS98
R9bOIvq4dtnb3z7z1Iuyzvd9dx2T6g04CwrPs4jJjceUx9betQjL6YOVCwEif5pn
wcFGCBYWsrrs3NU7WdBWZJC+eYcgIIbtXznvnGFrd0bu3M0ZVIO4Brq1zcD05raL
fcn4BdeXxoqyWmkFiVdEQLH33XqtT3PJJZXl282A/rqePJLaFlZ66w1x3pFO51Ev
KA6dE+5ZMHNAKnLH6LxnDBF8rS15lcsmn69yZtZle+5L/Ash6z+P14Ybz9VGzkl+
TacY1pxeQphW3PYvvD/9EyxyzSp3DDRgXKsw+aUpWlfaCPdK8OdbliBfNrpxFaUk
P21OMHImo2e9nwdK3iJ9JwWprI8pLePBIAWhD+XHPPuexRS1E/ILu7avyXvKrfUK
w9cFJdsoZpE3ShtYWua1b+nEW9NO+oQ9MgEf6HdMuKuhX6GQThszd4MDcrCxan6S
1Jh1rjY4LWszYFWEmsZD68fEkeuz+JNiTDiDn0ffCaxRaBQ73F+hdpwZ8mkYDT5i
43moyV2PZXQMddPEm62VpQgbVb8Sr8vJrdnHwVyevaqgvzh3hNX/jrp7QU6RtP5T
YxSdGC+SSfRSvBOPBt6+gZ7HB74SOhTTLSlPyW8bNrobSbE0E0WFWGQZkM5JP9dU
hDQjz0UK4rwZWEdj2sBFF965GEkQ44owi2YFOCuFCuWZzh8u05YM6blzRHiw5w3L
e/bd+y4S6Y6rOxWWd2NC6UkAKCH1L4MD0nDIIE8i6ZBKsLw9h+olhG97AYUsPCek
ZAKZOwnryQlJohveIyitsPTeO4+jIfrLMcZmdPxvrcRaK6XBZKaVjN5mkxvjPRpC
o4XuPhlNBmexfoEL3+CTEnHvxqAd3OTVixUWST9h/ZeVFw7B0nZF0wHNMqLlsKJ/
k4pmINaP3PGJ9QgUyb2u4GVGHceAJ7U5GODJ1pQ4na7bUyOUxg60wIkgn1bxl42A
IiBGXbismYI9ynnok6D6ONV/zPwJG4lrDCYIugnmP9ec7oKr0VCsx3AptY93kI1P
k78Py53RzWYT6Xr9sQQc+Q1o8NtCjQmwNLC2fg8UPyo7RkAYT00p4SysGaPRabj8
1G0Z9UJKKO7a9wbzKynIPsJ2feoSpUqfh6THMjFDwhT9XcUOZDd6QsXR/89CtGGZ
9gEVk7PyLN8YCyHe+t/mFdrK1CVSRwEaZdTs1O0T3+Ztxwcn6/6II8ktqx4KoSzN
XsZIg8eIBUU9TMgbx9mZReD9FQYxXyNYb7961MiIkN6rBNBLNA91xHP5qGbR0QsV
ejRqnIQt4HyYHIjzcxb+eA==
`pragma protect end_protected
