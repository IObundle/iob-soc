// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:15 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hZsxwvkeqfhM4QEaA0AJgJeDXcdbfAShc/dOEPH9X61v3jnYmuiv/sQ24rVQa1YU
nEP47LZfOfr4aSj70b0lqz6z9Caqv3PWIwOl0uM1zN7y2eRrb0ObBmYe33Q5xsBF
etRHp6sIqDlAdmFosFOwkOdgoalGOGL0IEBuI4aRhHI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5920)
oH6Kk/VAtXDzYrQPF1YfL++cj+t47dd6IzL1qPyqcTXGXNfSTTPgEfJPFUjNWVBw
7vs2Vhf7x8GMannR/wP5IL9q3LBwjyCVn9T+rhOMXOHC+Zpr/BXoh3zdDWRnvd98
RnbRqzgoULI4z0pOKTBY1B2nPzR7H4wMt/hOTPp//iYviHfXLLAaIl5UnN9lbCoH
P6Rzqb/2whjDo117dV5L2q5lTM3I7F3YIbInbPiPv/SFCF9c7uklP/LcI2PXhF6w
+IePd6/MhZij9tcIcSeAHEe93pNFQBXUeoLtuBY5nivHzW/O1Nvg7EgfywhTn+1e
Py2xzcTxYoIllStBD3Mcn3XU39uo2RFV5NbToEUn3qKxhw65CBl7A3XtfZ4I9QZp
JbMrXjsO/cqH89jIDIMPH/vKTAJcZ62EOsZWzHd292IkMtMAMXI6FN/G56xzda4O
jMIaXje5YDgbtaSrbEhwLVUEOAej6oVahaYy4ZYW1bJkabWVNm40GDxF1oiXuQPX
Sv25XpDS++YAUWwqcd0ZThV0eF4VBr/Q0zAQ9+aE9Pv01PnfM3adB7j5HVbXbrvc
0a/lJpnksnqhPC2DvEDw2fGSbl6WnvvEGOnMtzqSPrKmVFIiZkdUhWjtFRvVWqvI
/sKxe8NOKMzRdX7MgBwVGzFFTp7dVV5lWfklOVvEymTmDgF9dXBmfx1RrvykSlM6
1NkFOXmx2Id+UOcgOYj7hWh/EAsgMWTpyI0f2WWxkTC/ZCJ/v7GbLKfthRmaSVRp
vZ4FSHEhqc8rRFRo+5q55lr8pwLUAl9wDAlyfsY9OnUDj0Dk27V1ii5TR9og3/1a
3PCFGiDLvFNAszMtbjlwemGoBaMXotaWfq5pvEi/qCnb8Npu24ZLFL70uv5mSxaS
YP+J6hg6ZiVGAldkEbMG8T10AJQ08ICRahzwXduFGj6xBoRJ0+5knpxc6GlxF63l
eEWAeb+JbqUODKldtG7NRdv8aj52cY7DAHh+Fg8d6Cz0LHL6rD0a8korbGsCSts2
+DivL2Uwmdi2EK3WSDicFcRU0f6WtFdT8l3UmowbP0ZVSwJTAN0bR2+soa8B/93w
Xc5/4OmhXCI+YURmrXxDDwmVd59AlXPYb7Fd8swfvumruclRgITa1O0LTKJUciO3
p1hqTes41DGLtIIeYQyYrzjB5GKXRtbPGA/1vf/0ffSwRW+zaTMIiJwKDyndAlGG
1rCF/UeYy3XKudSM4em12Jrh7zz3l/162DnsqB/W6KegxZY+nQkVmIRRGerYdkiW
5YP0ghJYBfmvw/riYcmhhue2Eqdu1O9Ft35FEUd3Ny7MX97WHzabolrhWEusqthD
DAlk0f74aTFw6e6ojlUPs8LbrlNCdg0rLPIaaJ7uA4lKHPuZvyw0neim2GfoPrmb
kzNHz34bqFM6BXMh4+gnMw0qlvoMkGXCvXaRwfSsjziHnDT79GGlVhn4MhfE3quy
y2s8DKif5vzviD83hiz2scRTW0/5cqPcmtlVf3Q3L4npwfrhGxy8lpxrApP/0Rvx
/GbHT7xaVbxmv1RH5/JIhBVSTqMuI58TII2IvDPt3IEMvmYZuwflfQicz+wyWpHl
sEJ6IwggfOvY+vxSAvdWL77OIkP+XL4tTRPxN5kHqqZWnzR27Tqw916qVKxVxig8
9ZSAvbP3fbJ2O7zKRP2xecOKIx/FXYLgoPIDVn9Ny7NeAGn1qzUPGFex5AfZEfQv
i+QKcfs4F8+fxQOTbuXUwIiqW+ubTEL4Eaelr5+crXrn8RASGwGIH0Sd5zXvSGea
vY/xwcQ18zcEsAacKy7xt4y+6KTKue9M0uvJBc1jHXCxPBhbdgnuR5xh+iYTbckR
aIAxwaRbvxGvIp3TShvK9o6BzkZvQ3L+jkq77GmpdJXHbsj7lzcPt3wvqPxAO35e
YTDzK5zAAnxBXJkGka9O5zL7k5h74kNVnhxSnbXL7xhJne0NmkuN6vURBnUyNrZM
+w7+aEE44e9CcE9GqqtuSwbn6BAnF3OypAP3lVKXA2jmWSALXI+GahFBJkpB3+Tn
34Ob5DFJ5OjEBpZS6rJhEkZqr5T7kj11+BtFmbTck7AED6sd9oCV30GrFRAE++Kj
7iFeTiCiPqM+KuOr2Z72hAkQNWse9w50ug72tm6GXNh1RIgu1QLrC5szXg96edUp
4+ySxshrVGLb+ACo5JkaHZd9/Hmq4pwIhKhq3PhBbcwd9QUED8TNAJJnsIXxe571
O1h5tBmfTi37AXdh2SGMwOtZW1EDifmc5o5zBK3M5fSvLfd+METJmL1j1bgSHF3k
lLv3hF3uIixwIYVdbxpyJDpS2roGjaTa4O5MBsoWMLLF35LDZQNzT517r+XWxJuT
IloQds/8QWneAt1NQnn0R4Wb45sfDew0c4iwqcrdl5/zprAoMLwyffoE9dNqVpPF
VOpXxRj86SDnmABmoEhz2DK6d2xeklpn0qb1Oy3x2L7gGxOABN+B3ujtHrltP6JY
TtJL+MGZkWuiqyxTt740N/wzI7F8Gq3sFUXGMWVtfMFvmGxgjDR45W31ymYUyBH9
+dIpBLRK4/22guYmKbKa3IONGcBnF84ZVn+YPAHusKmCil2ZJS5tekQd4xcqshKS
g+DhTq+xrZPX8G5ebRbOXpn9CTY2qI3rvTXv+2vDrJ1r6q+zNsDerVq6Oxt2tXgZ
KIvaEdzCReUiINeap9GlytofXHOsLbw9t5cm/z3yPgA6NdgVdDJU/E8AVau9txGm
UBrdH6EuqtroSl8lGK8MzdHCShnmX4AgqOFSxSqbHsGtqcyFN1/r68UhMsvargpr
FplJZMBL3tt8f+hvZGSmvyVjKUv0+O3qXvYR2UnZ25Y6pF65Z51rG+8amRK8c7B8
VdVkwApwdju+yfxmeTuvDjmcSq/oniB7HAihboDY2pemY4Vi3IRHFF2STsceCDiV
e+AH18UwbjWJwkMjJPFUWuEsbCTpZ0ft7B3kYkZpCfuZyhC1Yi6iO5+1PoQxAX/9
BRd4UVT32j7Kxt9YhEBU/Dc0Lwol8DOoVYP0poQkVpatfvyKZNt3HbGmVKvIDPs5
+cxun10h7jtSPRA3xLSCYzA1cruSb02NzIWwIApQdA/S4sBGOVtMYwMX+W+S9cHc
OgfVu5AdQrPAQyNtKgaVm8QpIKywD+jSmvUSEwPTuznNBtlOoXtgXVo62wlk70rB
8PhdbgMKCIXVsIbkM1mc0pFnOYqz+/WzUPeF/n6g1yI5I6aEbFeezw/eBPl/sSrP
qax5+lQFuWQd8jYKCoYgrNTp3zX1SZrE6Hsa2o0PCVZWCGcFdeohBEVZkg4ntoY2
81as/R2jD7AUibiT9ROTDbRK1mndCrYvQ5uc7Y42pEwni9Rt80HQodrcUZbweMIK
aUEj6c8pPHNTJdmCci6xfdT9JXVegv2Y4Y3/b4TAGeB50vG3HicKpFad1s+k0Dm3
l3oBGjHO45HlYmW3doiuQNH0V2t1WhCXZheyxReSDOR8hp8YXuecMGRX5w4D/qtR
8C33t18E6YmNjZrCKJ6IO6ISxfaKMeSQK3cqoNfmEo0lPhOJs08TCnWKT3gDPcnY
LXDzH3xBEmNMXZVl1r7Yz8v9Myie0kECDf3e5QY4+2LnZm1vM76xrQ+UierWxMKx
+Co23ZFJYu9LQ4Nj/830YkZT7NIMdyROE39+T3MmFW9lSvMMmALXQgEbOBaKOBlC
ZDEl2/kJklncxRos/411wIUoZ9YITNkD69Dy/ADGOaRqYWEg+gUDO4HX+I5SBwdN
QM3yq7ZttdoN3ab/cwY4ufgyRi93N/7dZPq7Vs8bwYtgRPcl1QIEsluMZQWnlR+w
T7ijSXtGJ0yJJkUa6VYFVR3fpmueCcPfAVngUOoWiUDRoNpcTpTFc8AbvsELix/d
aaIm+19AbCLtFuEgr/hmN6b1kaQQVH8lJEnqgGj/pfHt1z0A/4PXaWTuaAGdtSi8
60sh74GyDfN4cg1ncuZbQGGMVR8SXuypEacxAYrBQIID2bi3IxDfWNgtVB1WRgjX
Ii+kMFRD3xMs74oDAIX13QPnXBgsua0mj9AZL9ZWX8kuwxpG67U/2Y35dap9t52v
4MNFi0TMDVuoF1vTYn7jsnWjcrUe7ZE9lopPY1TK7c44Q5qT9kflAIjLW9EMsu98
TngGiz3DNljhxL9BPUPUZi+G/u0m6YwBL49Cau6AEGJC+b8vsG6mKCtrKq6qfACT
fN79D6E5h/gqrIpKLGhG9E658xZ/ASwogG/jGqhBirSQKHAFun0QWfoFc/23dD2N
P2nWXZiL9Kou3qarHdoOe41USeTyhUvjXaXwgCGK8PuZzE+5haS71kMSIy1m2ZIB
XpmTKmTzy5DihYT04oVDf8x/ezTnuLsS9gWHxTNeZrt20bSlON2LOCflZP2I811G
nP5tb2NJT3MA6osEZnHKM3LdF7+Z5quzx5qCiRi+/JCdH73AuPnxzTJ3kKDh45/a
uBbKQe7IJISKSKWfrsSyEd5kSX7Ls0M/hAaQaEDgrdkzvINiXpXnp5xI9RTgdiRe
lFCx2HyGCmQX3eQUvK/G2GfOU3Wwa23NReBWmaFdmwFrOPDvUKiCASTUevNXF6NM
Yz/XgaIsWHW34l4r5oELrdI4g8g9qWers6P9jA8ceMLxxnhZgDQH3GuPohaN5+Tu
O9l+ZyzOj8qy8yfWifCeIKlA9IG6mSLCAw1cP8ifkv8QsF/rnOMiFxNf4qogyXxb
Xt2jK0HlvgONs2BF74tnpc4E94RJacp9mbVzYQx90JuIgqBbFJzYJ9zdkUvN51rZ
oKbiTMeaJJSUCJr80+eTx9nq8duQV5NPvsft+LXymgVCH0N0hL5rEZgemxVxXhQZ
/ZXHd99LvVKO3faI89MaBanqo0ZiWB9X+bcBgqqh14MfRnCYLbdTjY24h4Ycm8x1
bqQ8fSy7yo6wee3JjoQq2BBAbL4MXrRMNd113Ecba+26mXu+2O8EO0rig0Z+/p8E
G/jkiXy7MmNiJJrFtwQa8GXMV3E4M2bi8DcLKB+324K4knoISRkGkvYEa7hVZtQZ
2AkT4SnU5aBFKm9okEFaFOg/chYAqlI3qZahG+MRw4X5RYMgh+IeTFUJUzNqEv4R
c5/uo0zb9DSV6mXQXFEB/Q/OBPlqj2sajwaDCWTSAfUn//pPb8raiwxhba/FZyIu
tgmOWHBqbgqy/6syL1dvBr4ki7H2ORD9fLxVPrRp4Vqzalht9LK5+2D2O6rKmo9H
2bcN1GoM84N4tvNDO64w9WO+68+JkStcOQKaw7/iMl6968/hB7o2bOXFxDYEcqTH
C17uNi55iC61ORcMZlnr4R7qQZJfyi81F1+VjH+AxqdwrZV3rd6f+GtttlLsAfNQ
EzelJoJvHwNEtXKJr+YOiqih85t50iLmTiUIPg0GrucWzNVBd6OveUHpMpX/Bi9o
Dvi6TPsNTODf7pVaJxsBVyN46EG9A1gaHc0+LzhmOxCdTZIYzk/NhrnpEPAxP/IK
BReswE/dU2rbo4pIFCUDlNL2+d5Y2sGnFvXj65e1AvKmj0RDsYwJx8Pxw1g+9iMB
E0wi1cZVrWe0bMffpAvO/f8DUH9QWGYWWYBqFuUpvrF9smaUwAX9IIPRjZQYg/Kq
ylDh4a8aAhv1aoYZFjejpif3eR0w1D+2IwkVM6fxVFevQpjL06q5jmRihkMlTX3S
rJ/u+pg+/AyM4Ge3Q3AvyqpXqQTuy7WcfR8ju2gqByX208y1oqYgagHXr2uPxOSI
pST2g28mPHtexSJH2UR6lP4K6dv+YAC0rW7Iy8G/8fuqNF8Jkyz27PNgAQnJzrEp
ZMlwEGxJC0W9fN2cPdHghJozGV4CTvGlH4gcT80xdnvSQQ5zSI4I3EiO46iN1pzY
p5pAPrCJdHQePIBNDIXu4n+yJ67fQp75RUCExbhdY3hjrpbVLxvREhJNnN87u3+3
I9CgTLt+L+EBmEkqe/3U1vEys8vEqk+Q+NXAy4F/eF+UWhSeMsCn32ZHIvbWvQ2d
Zpybe/u3v0oaPiuZtEDe1fZwJZWua95b5IWHNdXDMWsg5/xfX58I9zMh884u5w+T
sg1Gb4NIlZGnUsy6C4a1iTYIVd44cKPvrqKiNps6xoTudA2ERrf6Apz2cmNMN2dP
/IE2NK+STyynShYb49H7hvsPtfP+GGZClbVpYLHQqwF+xLyBxy6G5491D86VpmHN
NyaJAqwVndH4a0PfROQk0oTC0bSt2X5w0/6jucuHazjIhHe6aXocookAPNhT7yv5
8nJyX19OZRRcYnjlqUsaE0XOr8zGjr+UqJKsioVD/KyW4iy9xrBdvx+czWF5RMlE
oOYuq6+/cU1FLxcr63bK/njfw5ElQelgPmtzErFx+pkaVShvI7I8RljCMyWfIywp
OYPaBKUJZQgga5tewH/Z1l3dOQczuAdc2SwY5zjuz9CN9h9GMCjK4Dc4t8HViY5K
NkO3AOg04jZTz/wYBZZbgGBRamvD6luMFbylT5du/RO2Vc6iiFxB14rGiTgOzgVJ
aPEUrK3iJHOqgplxu58646zv5wdVCopIy2UwIW5rhQzTk8Jid3bFbZsNI4S/pFVi
lLz+fN2BPRhPPWnPwPV2CEIn5b5GUluHHI8gbnw96ZMjvvhYG+0KmUVI+Qr1Svxw
yW06101ITGlV5djQh3QafHIRwxmMN6m67avNX3PHRdbAEhw2udK7qLbJ/tB+Tijp
y2S5DBcijFJt52EPQLpUAqpxgTCZ0+f5cSMTPvHeHSZvuCtNPFPSg6+ezfTTQCCt
O2T1voi5c+BdaYRBGLVdeisAfnou6K7pbYLSxcXJ9FdYZ64QmER3wOij/tj2yKYE
XoK0dEe00NNS41qlcNfl6OgHOHajQGQdq2dPwDf1X0pi4kKTC21JbmavEb2oWwt1
KRexDtVvIThHSCgdugSN0DpaQUDfdgHv7sEYodynVLzxfQSJ/W2Gott1Bh19bly6
p/R6lbXePMJfYOKB6GlkE/v2YQ6kG6MX0me6ccvlvneJcgF2s1WqrY5zqFTV1RXU
AxLpZfHlydFzFS76z/0Nc01t54a3uL3bvhaIR79IndlQMtMAapuhAfFAUrhC/1a9
Y/JOYxAA/KNrjGr1zZSD20MFfV0q0+v9QXEutDwbS6EWOOo4LvIJBYXmeQG7Bb1R
xPiluDmeS9svmm55xG8jElYY9E4erYwtXUZpzCFx9CNswBTU12yrPgzOOPwo4BSY
0ur/YznN0iPYqIRXoiei6oBNK+KVM5ZNQeJCH7hop93nk+BKrW3Ct1Y3xEVRo7WF
SeFJ2YU2t9X8tuhATaGRF1qXimwpHO6tfFOo2F/Te9crqU2Cyk7GMwKJUIVzK+MT
squ5wDXXvDXdahO31OgvyUm6xL3CdeYHKN/gAhUZvHfyZVROo5BJ+MM4MMviB6u9
mpsOIn1Tcav299ckOWY5h/bmCKTRDPKarakXdFr/Em9M4izaq9sLUBsFA3Idb+Sd
KzIzanCGncfTStHHUFskJNT5sSrPCGKPb+WcpRo+1TwpOeDUh7T27+S/3ChNUxJG
4FFIhmIrKbGlBPo/oigXAADnkuXMLCIOI4FxdDcdLMWv+M2sHIZGsvxyU1heCLFD
zWh2L+J/grX1Z8GCMLnjv3g1UtyWul/ZGdjTTy3GDIs1ZlSn4TVBGR9+LvH8r7Qg
SVpQ8UpXfSb/w3Qab9EmIwY7M7BnED8Hpbd14RpsYj5fA3m1OxI0zOfg1VaBpEOg
hbjqGQhrH9crW7kJwYQp4Xu+UeyuGTZZe0nULlON+nXJnkRRk1jm5Fs8y5AnOngg
Vc1nwk3v+m6lE1BcJoZFYjL4m1DtIAxV6g8i06UtlKaX/R7f17cvEyyUGSeEXPIV
Ui7wj8ad9QCwBMfbfaxMOQ==
`pragma protect end_protected
