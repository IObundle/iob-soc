// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jTQDv+3j4t3UdjBGRVTt97G9ZRkfsbW9SbvuL5UAIRb3DVYgGyyl6i9M5r8GCLof
1mxzDpmYqhZKV3Uoo2NSKX5tg8onSpQhLPJeD0IUOlUF/Ojk5atnjivFSQ8xL/ED
Ppbc4P/iq8PRcTbBA1OvpdidMkxxXtrHZl1wzxbGPjw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 178672)
G113zgThTSiJdXb73xZEKhlcUTAMiPSgFFSoQZ+4GTdRdHun9eo1wiFng9VVkbE3
/D8yEg+fxaPzb4LwF6YW1hAw9vxoESjxXrXfwooJpISPn+ADMXvza3mT1NewPjBv
sESU3+COJ5g58pBHYDw7GIlisGW609gLO8VaNE6g7efP/u44mf/zyezfyxvnuQhf
n34crMqE84mnOYCyTU+eCxEN1mPallT/QmaPf7/bg3mipLM3aNo9AufN6Gw2aL6T
n5z82I2rC9FkDFT8Rc8iSO7zR8Qes/gWkwo617pAF31ooZpTfAfhsP5Fweq7mVWw
OCOzmzwQca7fsUXTK9CDOVbcTuKMP5PuIMzrlgmQp8U8BoUce2YbJtGi7gUUmr/c
3COn5XgoQuQLfm5rgSCf103ZRbPoImXlxSDaG0jdV8WvZRidm7qSbGbmXQwAiWmM
sDbTUGqvKVG9OmvCpTYej9iDEBJ8eSdRaJzvewmWlS0fE5Cl9tr0jAfFgaRRNl4G
N8kLFP/VvT5/QL1H6Gda3hpq55TzisTjPU7GcVjM5lcj4YexD2Vth/G0DNNR4XJQ
ReTT4bnF45M77pAHY58wd0jfwCgTLLqHPjDi0LenLHHrZZxVYyCttpauNZUnbvQW
AYKk6gBbZSFHhPCCFRQlz2ieo6cQBDBs0wCPDjQ+FfnunENlzOKuDVYLI9nROauR
oGtcWBddS7esBd8Upp64ijB/OtsIVc5RQPTTG7m6SQXiKkULk32PiL1n5e5fku8b
URwCqzKv68JNZHURjFKhzwnuQraQL30yCIRdrbNTNvUGC0CTiDkt0iS3HqDQF4yN
zoB3HvSXonGyhlYIcUQNbQ1nCLG/pQoCh//nQSL+crYee/9snxBSS65UY+F1pF3p
zV5/+CkV855U0vtjWvmLfR09Vc46Pz+boqjXUNBeetdnd8qkc0IiOTVC1s1bW4gF
LHRFIH3ljVBu5pAaij8I3EEYpg2Wi7uluCuQWQXD8iweSVQ73GQphn6eTmm0LGBz
+NZA+Z+Rbl8oa6CgMRA2EJRxefGD3r2K/FD68Gh0gc47FDECPK/xD8lfVd1TaXA5
XvFxuN4Vug/Y//8k8FrO8uXodBRnxIPhxYd24p7f/8Cpkk+TedUxsz0jFgObcljc
exmOeZ5kMoJOceBYtDLqDguNjXRLZfRfcHBc8etlqro0TrVbg4fwi8TAaHmGKq3Q
T/hsT/CGwaNkIfU9EKdY+NgnuSEKJAI8K44MY2jTP/xuxf4wd9DGOFunfNipyUez
WsuvCAIIRvqdqChEO8xgQQW2/O/EUAC/RiBLXpA3Sd7PWOU+ytLdZ1ylzZa/14wA
YqlHfCksTcY2p2c2LAYURpTB/b6KLFyry+jE97DLoQAK0vQ25+wwrK9wzoeXO8bN
TtAR+L6XRciXsujs9vT2/SGqGYl0bYqUJwmyQSyk+bkC5RY7wXMwH9Be5C6tQsKX
SLUjsISUD1v6O+9XOU0aoDYxU8WhjIX42Ox/x8GW2GpGHEbZzqxwhXnuyK05iy/G
5Y58DhykEVRagGxEe7q60zJ7FDwwX3mT5HbERNOV0HLczZy1wIWYXkM0Llf8wk2u
ulJy1OpObvC+TUFHc7c1J+n5ryK2jPg0aVF2omo7g/uEf8cdIoRzCimDLXXtUFA0
0+nGY3sk9A0c01T/KGJsGJlMzKVp97cNCMYrq4ybGsYwQWzgdXt4KNHK86JmNNJB
wuPxC37naHKENcE5N50pDIvfgMFlSaxrdxHm8cZannrW1/cPU5YOFd48y8Tjy4SY
Tl0uhLPxy2YbAOyaXo161d4Lw5Q95p9lS9c7hOHJBM2dZQ8rWKw4a9m1ua/wAqaT
c+M3+gOYGOe/OBy+uNwLHiPAZYRrB7gLshzYTxNEHwhfPznn7CbTHfNQnzd7BirK
iejwRV13QIVm4OcIehrCyMQxduRqAmkcFKTrDY5uB6j3u8vRdBAe8MgMI+couJxb
lv9k1Vu//pdKZ1unUAnVl1iDJGPsOewGZlt7VRW5rLZLRF3h1EY3jLqI2e+5HE2v
emMyNJOfCfcDlqmqODOdcMkCBGf9uH5Efjiv0viJ+S0vJjEL7Sk7fihpZC1efgt4
TCToVWtTIZwJtmkI1z5aJSqNxvSUV++1fR9LO4PEdQmQBS34lAwOB3RxFXMlgOV4
2C7Pybn+gJgU4Unrx/6ne4+QX/ocV91wSU2QCEcGJ7hmTik4S+PfIbiHcnZxH6Fw
ltuWtc8mJmk8qZ9mtHJKqOdXYfijOZ54FX2YgezM7JZO8jFOXmxU/CvUzxauhqAx
TmGrt2OJiHQv5S+u7FJBK4dSBOpO9zo5nob9g4+yKuoCkTpAC/PTqRTwuLBnbNrq
7gMxGt2NbhEy3RBaAVb/An9UZVvTxgFCZcTeBxI4j0JhpFJJmd9YHqJlR+SAnjBE
uJoo4y3OzkC/o3WD5bLbVUMcFbJSC6B6Vj8Cf2EjsjZLaxKqq9L8e94apJG4mlQ3
mzZ7YgSqRUc8ukVPFH/m+reI+YqLUeeeWspYHa2KUqUIM3FxeHE6JM4ndRdMQB8R
XtyjCGLImDtE4zf5O7PUwYzAyAev1ykYWuAhGJeFV97lSdsFbz57fkbyS/Zexh8Z
jJcWXryhU/RY+a9+AoSSgaSxWrKhUSAOcEKh6z0tBLWDMa4yxmJ3Myx7/8kYzL5a
wqwTqZeZ5hXIQeGhxuMabMJfp35vi/Ou9qRtuG6+EY2UENfS6vufWfSrQ4M8QHaN
CujJlWf4QtsP1YMvAydopwW42Pu/4PfwPIf9tOcRwe1r6UAIBC7cUoTU1DDcUvsV
hkj88MvP720P7A4x/MsGZvN8gJSjzycFA9hg1Wnv91Jm71AJ8L8HS6iRaJ/WsWFb
9jju3z8fvVtV/wqKMM/+/i9UXvGL1BxaOzZhRH5vnyBD2SO2rixO8tXfrjuzGdX6
SGDlkbkSn0OBQoht5hABfwKQeAHrVILyQi8lEHsptMeXB7G9RRpXEXFax5Mro97o
MaXx86lTE10uAMbtVAGwkzHeCASk2u/P8xpMQezVfsLbU+3BjxIM244+KSbyHnwN
0KA/0l8DKll24irJ0VVxrH/WZEibimbsb6iJ/u8ThqF02TgCNwaWzmXjN+5ni2s/
dWrsmLG8w/Al0J5krf7VUuUeb+S+UwCs+eX8eagQ7Ra7LqN3CsaiW6IMEDMPvUsO
gb2zWD3LnRbTtB0T6WXwAK0qfD/9Mn7N09e+4jX5kFjNU0VnGq8vVtg4lchStVqW
VjI4RR06lOYYwFaTqDBbOQ9imO4wco3+CNzQ7cyxLyj5o92mtfhSvRg9p2d/27rh
kWcSjucSg9F0OnwAzdI05oswD0nPqk+eodYsMXAlHJuw9kpdmAA7LG/x+BIhBfa8
DB5quwB9gHNHVJ5vNqNx1sL9zbWiVJpbK/bmmznFhBytsFA7mPk8pjWvqcb8ndig
30LAb88v+cm4ITzUPPCYA382ctb8jYWBKHe24EUsPH0t8wAx0NvFw/LUXuGooEdB
c47SO04PtAx1Xxqy+5TSAvMBwHLHDCc7NiXm+GSg0mmjoyYyoK9DevTQTBUi/G5s
08KwJFKG4MTjdaFfq8XEeySFhH4PU3b+UP5bjD4xXmp40mhLvSq41ofPFwdl7xwd
l4Hdx9NvZF9yqgXrxSCeEmc3jDnXnSuFMPqOOqHjKWjhHUQqS1wX9zZ0Cc2e6qci
eJTA5MX6S/Fyx5bhnnidNk6lvD8nZ5TGxD8zdHJtIw4gb6hcRR1mkMW54jlVAYby
szNBzeE2FjPFkKmx+ci7jZDV6v5JUZAqYCtbxjdErajk5U2RoLeU5J0pg+W+/WKT
cUlJonT3k4x/DXon7WLfr7Rg/gpmFr92i94ZDFjg/qz6w9VUzOOHAmQOOUQzQ2ir
I9BfGZUuTuQs0RjmF0damT83m+Gpw3lYhgHO9TBcyw1Qju484D2PNBHKlblfgSeT
zqZEQE6gbRoh4SgSUdh5GwnnuXQLU6xR14b94BBNjcpNDEGWUuX4s4gefK2xNEDd
PPz6sF3qIZ+mmceIZEdc9pWRKMA5CoG3BtKOzJPxnwevtuL1A87Gkj3JoM6qGSAr
3RRBG0zJrmId/Pv3Q21jYl+D8PPOIMytGzcCCaGSt9c2lTv9hkAMM1pgdt58W/e5
i/uTqIGM6ql15QIzitDA1ZjRqHKkkmBGtZwOYno+XqT+U0kkJgUf2+5yXO+YsH9J
KmfKGASIOwXWo2Jvfih+WrxhoqNiaxZHA1BnPi28ES9reA/qxSoNF6lEPeYzHdY5
hc2xyVbZQJ2ZUsqC4733oTvTgpGK7whD12ggCS+hqz8HZXsjJK2O7xd2LycPzkxW
2CRnf23J+czWZyyRja2fTWfJUuetPiKseLZaTlm4yahMusx7A95gAhVMpUq1mf/o
LIOgJaa5MNuzWN5+l9ZSBCXzka8xtU5mPUaa+ilG74WxvY873jDkMw3+zR0Cyz7d
s+AWylqQQhYZ2RhH9q8msGOHwg0d9ORapNpmcHTsQYLOi/SSV2cbGplbR2pWwaIS
t/NaOPWvw/OX2wGPeedzNBgicmC8TsaebPS/GwAzrrGs7eIDUiAx53L16gomdB9A
6Rfilzwp4eSQ0AsCh7U6XzfV7AGDf/b0IgcA1XYN1PeP40+4mSIgnwAE7iBVxxZ9
3+sh1CjpatxBQb1TVYloF7KIUshmHwa433PDNuAFXvNn4KVi0GYHEpGwgjdGlmUm
cuY6HzIOLuvWHO4USWKoa7z9L1iUIPqmWqOFhjlGqQwOlGiFT2LXlZhmLye95gGR
/CWtJWscCLVh7nefTcJU/10QxFHU1g/qfj5pPmNtWXwNwVm0psM0pp2waxkQ/tYc
y6xN1f94JXVzi43aCxW/JkEXvjf1RHMzNDTh+xbO6GzL5aZFsqEdY0n6uwKVdwZ4
WJa0WhYGZ7dG6RYE7DvYVljLNpF1kHhesRaoZd49ewBeGkpjWROkWemsI8Jd3VFE
vNN5yYvd/HOlnCvxPiBMHNs/x3hOkbBQluWdJ19tp6IDIxeMbBDYKfM8vuy+MwlB
esINq1m3jrWuKsQ+Zq2DKlpzRmZyQw78HHYvPyUo5Qb2g2RN/lYr9/ad6b4nbyd6
tXd+dQn//Pec9C0Rw5SgvAxuaYae3fWC2hIhas1EQlPjLbqTJLAlvTYOMpFhLqUA
pQ8AISnrC2zxHsQfUVFqQTvhUeJLpHAC1QsZvg2UMbY/Shw3xk4cBD1rteBQFGsz
TqLC+5HtfWVnG3OQM87FcliVEeWoErIq13dgwFlqpt0q3dneJt42uo6CY/ihV1NH
epDwNhMBeO+uKqO+DvZRPxSTs+fuGZyWT7UChzKlWLLH/Nonsmdc16YJLWqwuBNi
IeMX3r5AUIBypM3WPp+38yBWlmR+itYcCps1oBDXeQnP9tGLNzTm/zCAPD7ENIpP
zn07utkYJNnnAPd+WxvbFQosTe7mwWRfmAHuo+tlO4zrYEtTT233A3k4z7G6l3/C
3kXobhbwotzSGAnRVnfQcyxEP6ro9ZsjFHQrwE0m7LVIJh4PvsEmGDbieSjOr7xr
97eEH9zhodxJve99HVad09AZL6cM5u70htusKG2t+a4o/MXTFACEjv/PtbBalrhs
dLMtFG33yJoCaHXgYFOx1+LHtrJyJ6hh4uNqS6/Q8w+PVCJcheMtazY+PM3fjK5F
NRZD5i8yhiYJjQ9Uyu00r9GENq9fnE16mPT6qz3c06Ek8O/pXksNB+atTUuzkjoJ
Z2kvaxhcG+AlwxxohtImpkmreeysbtj5wf2Crm49Kh2lk3lRFl2K4S8i3a+FyVUs
0yszGyYAo/XYV0rWBGxW/6FT6RTtVjcXfj8yEsmw58BktCz9k3eQHG4iHwgz+cob
NQhmt43RAO4AVPi9J6whclApPvN4i2trH5ak2d3/7gqzK0r87xx4E7wFWVu/7KeO
fmnZsNHfIgZdnGmtBIeySR7Eo7pYbd0wqBNi0M/c2hEsZhbQoeVrw2OiKkUoG/jq
Lv3YOL0FAByzGemsqQC6hvvCwduXyrzm8LypshMPlni8dcR6UIB3y0cIBoVKyDMZ
4l+BAeUyddh1ubO0M8GWsz5NYsjt/CEP072OavxXXEV7igG5StAnCHZmAuS716Fw
rQd2/FX2JIK7ydy2w8xAImMfDhhCqW0Zz1Fg+MmECUCtgvLQqjVFXWfoEc6us8Bl
ZIsZrODVuBQZ9cDMMZolDbnghJbUw7qrbC3CtufkGU928VVTKJJS4EcojMhMLE4m
VHVm/kkOABVD1DFJqOnlUEGSmSxMk82enPS4ZCy+hKFiWs+qgIIjWVV93X83Ksfp
3wwMwh0X/i0JWtkW5sCKj8uT8P1765b0qkWXcE0rRNWX7NAz+tkbK+jtFA/nEAYF
mI3Mrm2n0cJpfx4SZz8WLLILAmn7OdB+PecZ47GHaueYFLT8cgB/8LxieQQSpRFZ
KuK+CA7pH/D2k8FUUk/Y1rtQLyXqgglWrb8IqPeX1UETSAx97pt3NxJf2eoVIN/L
YoCFxJAPq0cNZSxz0J7Y6WoF0Cl/JGBvjJ5uqePBFEWn8t4SimGg0/2dj2hKKiLp
S7LqO1lFl6xnXPkqm9Kc7F59+2Z/dXYGXJ2rZi5nZltgB76VQYg9Yo4vXo/UbouN
XjZRPXtoAEkHwes372KevaFuG3z3Cav0ABAFMoMVDf6W+vCSZn34SydJC+sUgxZt
Ls9Q+GbcFSKhEYup2LLkQbiAWaFJHnc292iGisU7T0k2Bix2OHYQGZn9chA8KYfM
LbYHYiuKUc8jLKOkauGVvqa9cvO1p9S0+v+Hg/EfdcSA22744o+vIMXC0MFf9OvU
l9SQZWOLl02Kv6ojd+4JvqCaSHlWy4JG9g71gRWSpmMVzuO0tySrMcNjySW0370+
05k+GTgdn3v1NObm8myNMl1VGDrWjJzQNZ0RpfB9PCm7r7Zl7+ksdQ4ZpS28DXEe
uwkGaXC2NO8qD3dWaSIIHkDVnCmCO2QnKv9Z5Yf6fMOjbZWVDNYKARWm0J5wFHHG
Z0EpJMoIfccw9I98mhJZ9o73cAHMtzgy5HSeC5Ik0+sAwcnjtEVa2Eu9gIBVvB/J
IgfMpHpaTef+x6mdOl+gsu+uTmkbNRuhREBcTB6CgLeXGEyUaWwOgcuHONSHD2H8
75CzqmF0hy/b12rlVwDgR+dKhQIk/4rLK006/cHwhGo4Ns65cl1wyGLqjIAQUqGX
KC454a5zougYNfaokTvB6Oc8RxL24UMO7SqTIxf8B3UNfUTO4z4lhjLaBHALlwQF
L4qUUiN7JjALK8PW/mWq45950OV0qZsldUDA9naS5qzFSazI7Jzwe1Njq3vSZEU7
eMR69+eAZFzu4DdWVJ+y2ECtshV1QtV3ZFW7VnFbLk8Z9KD0lp4uiA3GZBXN+7AD
4A+WbymRsthDJDJ8f4N1yEE1Gux3EwoOZnhc2UrX5makZzOGDAOyppNB8hqDR6T+
MIuO8JW7a1LLNf4WmsWo5pBuci7yj12ZCWUe1+EKGtkQ9/TPxJBbJBLCgSbl8FkU
1DbRXly0r5NIghdfzfwzvzo8sFXqeQHerlzXnRH0oB5hgFvdeLHf6RIagvLZQGAE
JTHJxFkHnNHGEDPNpiSq7Ll/G7rl1+X/xwSxmkkOEQKDaxWNCM76iml1BOU5SaXh
dvGzonECmmwYNAfIdaLIScFZXBR7ALqhcI/nRwAWt+vxZtD2C0blq32AeChSlXwt
9apRpSFSK3dyvtXrm22aE+e82BYYIRX6ozGtId747xh2fBu1J08K8tkVH2S+hfOV
GtrAODuvWEhNz/uzs55yLiaz2ZaHTTJDFZ2URr+YfulVdE2K58sYIPYcGgmTVCe4
RgGh3ubc0D6DiUh/cQ4VCeHChePfE/VHTVzkouSK+DTmQffbJqgMMP+KC+nngrCD
yOP6pJvTNewQUrMmSFkRCiNH2rguOJiZai+cOCjKqKxhtvT5cFBif2OQ9VsE9Pel
uwNURvKBmNwzRQb3XeLqDMniD+pFIEtD+7NPILq5q8soWWlB6NZTsjMH9D1McQhe
VJFORZvDYEJo7dEX2ur4W8ePloAKA1+pO7uha2Yx5VFZ6oOsbCsv3ccp4/A3w0gP
n83H/Edtv1uKA39Gf6DvkOoLt+KENjaoZLHwfzxuRtSN+Y3sxkVvEb+gsQ32Flsb
CKugsUPiyTlDdhsMj4DaoZatwW3dw8XM61PTQoOYsu0oePeeenhj0UL1N1vYr/zA
lcP+Y16hXJmhDuryZk2Og5m0w/Ey9CECqcnWx9HyX4h1hs/xldYEiMav+UB56Asz
ofHizChpk+fy/+bgvdM72EhSpuOwX1h6Wi7qPOdqnFe67D4yQyu918/V4RSXxycH
g6dZkFpBnjEeY7NCWWYnaHuBLueFFXv+8OKJuXovb7O/vyzqD0WdI+tJodCBrdin
G2uofpBBZdADHiudRx/OSo6wPAsaLCyvEGH3YjxslBnwAy9L58IwBQD5khS5BBzb
rlwDdYV0KAhWYCOxWayZNg3zrGrNYIUC3jR5aqE6XmhDXPy3ANVTl5lk/17/Ti7M
IGVCn3hq0fEaQptagc8THIAaHN6mnjX10DloGfpBaIe/uuzkI2VahlIuH+gbWcvB
M8/eekGil8/LsPG3eIE2KmQiHrwGAEp+kGigBsKFXxbfnsN0W1PXqa95362VeG/J
ZJAiLn3eE6m0kkif0DHBPz8oByFT8hhCbpxtW5O7cBBw/pCzgfuUArXJlyu2PuAF
BnsUgZSdC4Qh9pf/HW6+wCIeYnDtXCbw3vSKqLEJhiEACMVFYDun1RgCDmPITHva
VnLBEwSorlndOs8v5cUBWyRZiL4d6tFtIIRCOVuglhUToHKs53msF3RzgKeK6ZZ5
whM/dIvmtSqWuefhANLp2qrAVzp9azsMIQEp8zEl2BMJguteBxJNpr6+SOPzEIUF
+GHgCtJ6FDGwzAf6pvc31K1x0p4SrwOFcRavsTbJxODcEem7GIfTzF6632YNTbUs
ung7/ZmkHQH86gjZZ0myQLlh1reUQsks4fg+j4HVOxfWXZQW5/45vJnUl8BUhZ1l
VFq6dcQdZWlSP9NmA7DCfqwdqxHOY0KHVzTocKVknGCFYQc5+7Raf3GBJOXDUEea
Ov3wnYSZfa5UJZ4Y9PKDbJCMLAUIEDHAsn/pr0kdQ80hJdC4c0IHx5BGIXueDDKz
Wb2oA801d3O9aiBJcTLwf/I43Zbp5fgBaOjOwk18awP7N0sKDRH1KeXl4nQdLefF
2KYh87aMzSvP5KQ+HdCiLG7H6BJdA5oASHYiWNdqNCsUihbAj2RvPATVie2hPYIn
HwIpThxuFYaoL+M7Ym7r9wbc8WM3Q/ifWYD6hESH/d6ZaiGCswXkz/xyBe5d7mTK
iRcbWJ887xhlmkitlFBbTfZDVubjgpC20TKU5//Y9WpQUDvNVV13PeK29WGRDkbi
53Om4rYemYlflmveHHCe1VIY5uGGrKFXvtoKzoX2ddAgKl5ModDnbc4HgT727jCp
iqZQKylBd4qa55XKG/2gmAAWgpHnaJbsoxs9w6UZWwrPn/CEPiVTafEX07qkAuqG
W4OKbn9elSyY0DGSJMcU3Smpf1ropQmq8lHhJaZdpoxRlhwQS0exOvPRy18XPt4t
fmXz8QrxKoRAd4MTdCr+WRQhxnqkbTDmFZpVBRugXtRigAAgseNiDCqWxHx3UAY6
j5HqBBeNLXoESy+HHGGPENFlxBH1XYmGejthacgN5kkdQUDnjbbt/lugVhQ2kA93
9EJ1LF+Z1mAHAUoybF5w92XKFbboegH4rdxQiORekFhcfb2Kfa1ZP5h4+cvXrUDA
CdRNvOBO21r1fzrx1jUCGtyZQ+Z+muQ2+YZQ4EbemmBhDdw3WUtvR7KdxyhlUjoT
UMlon5C+71nezJoa1oBrQFwkrO1KshE2P2OJjQstpkoYEZjynvlIUL6cX2EIPrJ8
Y85zQUwVYo+s8V2Gp0f2Gi7hB/PHXxy48CeebZvbeZepW8lsyjmptsokl88vraHj
AFZB6epjo7LoaG3Ur2HB8A8PaeSi4Rqf59dUFtFDtZ9i3xOHbPz1RSAw3FNckbjf
c/5sLFceQHsf3jrhWKE2F8g/CdcPhl08kt5w/iQGxufBlZXpLUCfMKO0YIl23wG9
laHsV/soswGRfWmzxAUwO+xpA7KSaB7jSVAxgFor4XMGsAOZt1x+AnrqFQ7Z7Sdc
XYN2RFJBN+tZp5lcZ7S+uF5oWyHPCETlNKTi8KMdnYehYwKO3QRBzAMmwcWw0ry6
5jw5EUPplsSQQj3LRK20uyV8r+e+8hkEH3bxbJLMll405dxRMpYxhp/XqTU5NArX
EsaHuZJUL4Hjv9QYU4YhPe7yIaqBPMlT2X925y7ccXwWKrx28Qofj0PmxZRJThwN
ovpwtTg5WM63k0zxak5HtC25ZUyp9W8OGBxzhUK0/GfHpTVxF6KBoBE2sPg8+Lh9
D4Eiv0SG4lzEIwLI5A4wqytXvBwzBNhgW7FY0B+906vJuqZWe7agyF1vu5PsKij7
udTiUNXaBsSR2sxvluVALAjy6JqefuqtpzE+hy2vehCU5RpoWmu0jeF3focnn3f+
apHrckaL/F1H30yxfT5/Vz6v+s+CIk1j3j8jAhN1V7UZGIRLyoCbRYMO4Ge33a/j
6C6GViFH8/Bn7W04eI0EcsP4bJww5jAOgPt7WXC5jwiHJbHBbLQ5mYF8kZ9Fh0nH
31HE0Dgasbz9ctKAwcfVix87tuw/BHhHpimvPy2mVVhhmHJGthItQJytjpSgOUMy
eIXgotHOjSPk5koqxfQ64MWfp5Ulpohnu3IhCqEKTF8Izq6oD/VwZTqdivysMbqJ
1FHlfXLFNX1O3LKuvhHH0b2ar9dMlemnkcc0/3VA6EWChZMGNviud+D62HhY5P3s
KChvdISK90HCJ5uECwpcJ9Pqq/q+nlSrWM+zYCc2oMCy2+s0O2ywJe1VTx0l7MGu
/u9tGCljHtg5qYQ8fXV8uCnfjUftroHaCWAMNDuDBP1hAi6ICAXKI2c/+vV4bVWM
km4YBIgQn7Opt4bn5sAw93IgZ72QT6EwHsvqVb4Ew75o0Jcd8LNbZ2D7HnKjz0dC
LNX5gSofxyB65841/IGovCF87xV+7+wUf9CElfDKB3WNMhJR8Zg7ZF0Qa4iJNtiT
7EuMJ85Ea+FPs8Ojf6GLOh32Z4bxNQOsKnhXd/OKiU2p6GKBhyrNv8td2QaI+ggW
9Ka8GkKV+HjfCgHXAvyiiu+IWbCABLpanagRXReXwFiSe0/nrPzir+I0f+KOIeL9
alAngnukZ505QJ7nzGwJrzQP8o5hGR+tsll9o0QlECQMebK0ewIG+5ab/JDiAapp
9vV3cL9BB1Uk4MNAD4w3or38cTFZcX8bV98f98gBmQq9rG7fSeuFCfK9P81ZG0vl
zJ76Y59Q6eHn90XeHI5ZIp/b7y1XXcXq69XE7I2JEhRt4/wJFS+mQQM3ZhcyZddW
ioAsd1XQ37J1j5NBtVKeQd9ZtqFRXjZLF70WlPi1mEz1yMezbvrZeVIw6Hk67dhL
hIreOge7nM6P4w84/BLSDH14VYchc7s6hnLwSrYdazCJQh5spjwLNNLkXnIZa9PB
90bA+Wb84z7soRY1dG4zVsSXYaByPdZK8l3hWe7CxQ2d3eZtsQXFDace89hRw2eW
1w4NwOhrb3ml9oRUmSO2tSFR66CXqHgcslU6VkJOTkxGCWKLXwot3Ozql6IH/GjA
dfIR8n9zwikRa4JOyDNBoEItwP3sQC131DvvpRTTPkLV1Q8HbfetaW/57Q0VV3cO
b5+lyQvVXBJJwLlaSxUiCkSv7PggdcNpiBgctps+qxdZ0IzVkkBuMoIYpJN4HYgg
7sc18gRCoeuVezM8Nzk1unLBv68DbK2+yR75XfUK8XCC8+CMAMkarC7bfLNr6Y47
nun38bvvxaEGFu6QxvWEWIMdYxImzWs/kU6OCYgNjOA8tdV8Nb9tup60TClErBig
HUrB7Hh/IlM5KkDMWwld0L9bkbDfLdtFp6O/jjREojECeYnAIJ0lK6KV4EEiC7n4
MpWLbBTUDpad9yH/qi3mAxLrmwgi39OddcQU5cTEIY439/T2NveCNOHfD+IrSUWY
Efnc/gAhpBHHd6WoaJ9eenpWtBeFP37CIWJISrQh30aKBZX0I3Opfg4zBtk76YtT
+VwFttL9IooTS7UgzXHWT57bBO6maZLNc87V6mmp5TjRogvleNl49A7TYUC2bMhG
LId5aedWBuQ7mEJE2t2QuZPa0kPrZ3cEz06UXbwExTRe9p8lDbzQFhRLNnGGiR4t
vt1fXngbnLdtpnM6DKf9dzqnxHp/g+6Vxb0S9xwI+mdwP/t6LeJs7J+x7MFDdMhC
mPHbumvLzOSzZpQTZ09skQUiufhRwhTyIMAHQQWfWgh+wklGVT45tgrKa6txBe+T
rMw7bKfuN1NgfNWNslfUHVyBluOWwUELRh15WoruUYUVP95pTQ5Q0tcKLrp43/r/
iP6L6lYHqo0GDPVuqsDVTknuOyA4APrl9rGavtLXsM6QfTwraKjDKfct2f0yODEQ
L1IeL3ihOdF/8uIkaW1o1c/GHhTe88wznnJsi6gWaxZP2t6WYohiV4bUpsZAS8Pl
9rORk4CsTODiI7XfFatPTNKqnMctO1NEs4esms5t9ARt198LKCPV/zDAVaFg7vqU
f6QGQ7zPdvh53nKtViVGvZ5BcV9B5CQ0b4nCS8csksEyAJg4KNdkwaeJcvbuuBDm
tt0l3OM+l8qxes4BDpsIBVfVVFDZ8dNb1l4UTLkO5CgETEz8MnC9NEFSdLsFQEm5
345j/lDC6EIP6BclXBTLd5GEqM7SXe76cpPWspa5DE3HoXnmwWySauYjy7rF4aXP
fd+EvH1dBYvJZYOVojA9+dhsa/j3bCpz2lnMm+O8lBHjHGLwiUhdcIEUSBBIYlI2
KbHkibw0tLBkfMJTGuhmzuviZX1Smz3fABo1j50u3dMInDWwXcn8NA1lQooJvTlF
GplXyTZz69aaGFkXVk2w01UyePIrxjNDleDiJpsqn6vO9+S/qNPKBGDzN6kcoRwv
Ab+OytABrC3m2tkHrhjj74Rj9jTRLq5P4gokFrfXy/EBzXtPNCj/40BWAaumMVsq
RXF2XdsbJehOih7NQrNPLsqNisZAV7Upt7fkn/fRfIQHNacWs+7M1viM5ZHwimJq
HG9lVTbSIpKxEt9IPd7F+iG1jXMlnmxPpdqY91zKKV3IeD8UIh4Y8OLRIasyJ8js
s2PNQxJoW05iIfptytJljFMIsxNlyxtPtVNJH7hpfeWJXW9k5xKxwVeNqhekkdSn
D9BZLpKkJsQXYBmhXSK2aBHCPypnK63BEKyNqV7mV6VVUGUaqzc5yYQg2deqHqTk
chVoi7zWAZEquBHSgvNObfCRM7KAS+q81rQDDKfB71pFe+OEOvObf1po0sc5cuP2
Bm2ZoHfL4JGwN+2K2x+P158WRZ+J5tgN9QUAg5Ca1P/P4RWOfw8sUwNTCZPN4Vqa
h/ijLADSobTwcT0byFQj32MRIBscyl4d/EWqdw+iSRKx066gmK5ov088crOzC87F
Xij1+nG4DXsxYfNely3P9ie5jLu6mJUP3j14SMeDuC40lUdcwEibjP+ejtmHcIen
O5TNXLmyf3U5LWvNTB7aLI5kTOmWG0KPqax3xGzNU7mbGlsnTT8QR9z2gpQrlbjS
5j/AI3AY+fLAIROuEuN6Y7UuSH+6IyzkGeh/4FtyYT+5tT/LdtC4PGM3sxGtFyFL
STmWi9jeFDTx1ZW/1IfHJRsi1OJottiqLaG6UN8FHqCvetl9ArZzjHL5/uYJMIGB
K76cJ3211g+hC716yP8ezXvwvW3Tl8eTCsb0kEHQRBx27O/9qAy/4cghUZYY+dCA
Gkcu7ZCGrUECOtCC1HemZilu6mvRbPS/QbwUQIvs2XwUvcII+ID0QHvMG3HddUFC
0dOCGXlnj2M5pr67FlUiaxi0wjsgBgNS41/o3r0ki8BoZ47wSMzoZArHS5tajJqw
EdiyU7fLJSvneeIbr8ZeqDWfQq6sV0+ZU5iL7o2MqCU7WF9WIsvf94Ty56Q5TU1q
TyJ5tSsTkFM6bzf/Rbt89+zESW+bDSWOkn+/H4xPp3h1F5tjshDg+Lmk2tZoZsUH
PY/Hjip9+cV6AiYAB+E1R0Lp7+dI1ZaQjiPJY0ub9OCJgINsbhcLfvpeotBn+XBX
9CXeYwRskp5z2RqN/TtYQmZoP12z+Suop3y9b5c8b/HsWL6oSzPtcTyoSOlLZ4mI
oezD+UAK6DLqmZtWnkzoBFG4r4DsDE+U40AcCiyMhw8hAxAK6b7QqRbYFvjl7mlq
ija1/JwdhZ8R7VNcT/LYs+pX5TUXCgaa7/C6bH+RTBlxoCFXB9SMIvbabf6gSlyp
quq8dWIXTFpbtLqrg9RqjD3ST/x0Ghk0zDe8N67Qa9mDSiGaxdGWQ33h79C1BKQ5
ePhfAqEJLsPuD4e8lBlnn6v+p4DhWbG1N+wAhyVsoTAn5/pK/UQRqWwPv3RoyWC3
p71h3E87wekjlmRxT+wTQAac5PU/QRmU+2uQByNY0cZoyKtlxWWWrKrg+y9XGiuj
iFNhkOYtpQoP2h6Hk/jYUTamwUM7X+6TnF2BZfhtmYHEe8ljEdQXng903yKADb90
1P6u8PK5nhYVYnedxCm8d1OZRKE5YQmHU+b/NMvbKrd0bB/Jn/9gawWlppKi9qRR
H53aJIIYHOCgf4tApqbEoztKX6GS5PB6EiWgIcy/BY8+yUkOppwlRHhjchbbsreX
GPfZMwZzLrc0H2pH4X17iOj99R7YmS7wE0stSu//TQdsO4zRJmH02EC2jjwyuVOw
rLWuIAqVizBezG/WwUScRxnqf0FJunN++c7K+AMTLQ64KhuJ4Axtsc6XqTmT1rrh
kz2nmCea1qxMMDxSdCPbZuotqZ1J9+XWzxuYbZ+I7gVodiPfDvlKXtzorKikVvmN
nAdn7Kcmdgqvg3BbymuW+5RmkvxQEPkYwVNdkfUSLH2Btlnjzbc3lhF9NZgP7Mee
1ufXFw8XdxreQOVeomqGoTilmQqdZaX3HeVDXpcHY9Rl4NE3cJJrks7rvL+J4RXk
e/UvfUM7KKwaCQoVW/VfwKISariF68XHK2q1qNicmMyPeFeEnavAocx2urrRHvcP
DKBoLLx+BkyUweqsl/46nwRfjE1Dj9XRfFF32XgBZpbKE4i6TMje0TPD8syquROV
8kAXique34/uS/JOm5WcPt/ctyHjEQwnsIK5OEILRI6aaSbo4gvxmPylRwlLQy8D
CpWwTv/bUnlbUAO5NVbNcl0zBpctHAYY9XlEWTYcaO6VzHf/9D3ErWow/Yck8RLe
siTdcTe06DYpHbTdmxpccrJ7uFCfc/RRr5DluBDddkOD3migVS3uuPJUneOit3TF
mAX7Di8x/PTSTN78zdinj8ywOltppQ/olrNuNruzQUOSmmMIus6JL2tuHtIDluhc
rpUUoIigOKQBe3lJovNGUcu9VM5t9QuW1lteNyDquP6b+dRGE2COtHb41kcZANw0
6+nYrMuVX2dp8m8JR8Zp/oPkw52SBh0fnzdZSSr6i4vxITT4l1Qn9uWreUORrxcn
obGxrQxPVJgjJBp08w2A2vDbrK+zAO1NJHSyttm7Lun5tyFopTMTVt5BrAwEh4HP
OPia1VVpp+axVd1RU3fp35urjDk2K5ww7vwm1kGO5wwBnAfKiP2rPNG5qT0SLlRR
cfSIcZBNudH47gzwBhDOtQtUePlCtBUDI7tuBQPxKtPK8a3r4uffN8ldwlVI7G0Q
i+0Q/fy6PV+ZEV3bWzhS+hiyXE2l1wrDbXI2KfLW9d8O9qabJ8uWc9NqpLp9qSOP
/7ikhtBNDy1CEK4xmwDyTrVOUYolvsJvMcsa3BZT4YLh/ZmqssurTj/zEtwabwKr
01D8/To/PFxgjIGdiGoA2JdgfLHA/yknTk8fLTXmNc3KJWtfgMwZURSBD0/RxTxu
vc33W8weg9oyYpIx++Yv22grSSSm6QKz+gcQStUhBHivkKuInNpnYSbBfA9TpaXz
gYb4ScjDKm+Q6abxgqXS1T+vVSpHD8smQHGaMKoz/b1wfBZ/5LPSVT5xYgUha3RE
xIEPRnCJsBti0n8dVUktn3pXtnGjONi8G6rx4lbo/fqESkcetE+ZziUpVWY1Sopy
+21mkv2QKFyEk5qBGHb10KIISUPvm9AcThGB8sfguOfbHQ1G2O0YoqL+CfYizlXI
RXKenplhxRQRWkwao5lmxJPsL5wEqDYHZJ795O3T5cLEguGI9UUCtZYnLDBqu8Gx
bi1M02ntvxsT8QubCZh8x3CY/Ak9gPaUI4qcYfx5UUQAo7PHy2StBm/wMnpQt43r
yfasRxKykReL544qaBos/LRWeR2y8W1cC2P4LKF5WFswX67NYEwicw0bdcdGF2U/
M7GBPqZcauHIH4RnsyT9NvruORjcpxeUKp0+32j81OleuewAb7x1ssksJIYb0bKr
MCfEz2Vp20mO+7SCroOTfdC7sPDDTKpHe9BOG6H3uIce1WrT8q2FtDjK9XxNWWsP
Bu/L4v2eQbsFVzlD/cnT5xqXxU945SwimQXBLdqeyUwDgv5aKG5nlAJk8SM4UP+T
riZYgxuiJGssQBcNaeuVjCUWXRhjlf8Kwr4B0kSodHVwvXwVxGiQrJKRfc1DdNEF
QtiqP7aQ9T4cJPk1Y4DZ6+K0Q22c6ECnz7RgsKZ+Z+LbUof/T6niHuNqfDAIYeI5
mu1tHL+Q2pNUn2APYrYa32EaUjMxCn8KbKH4ZKb5RGsN7DoAD+hkcS1UaM/Cu480
tTQVRBrLW8MokyLKI7rUFmKhiCTaMwpufzIZgWuKOAeaf/VqlF3q1diUr1f7VeYN
gGW7QFhA0tz+JBvWk+rI7AKItgdYzdHEEeVLjksXCxArNCmFcrSz5TXQiiY63mNJ
Ql8LjFtNJploEJLHGdFsiIFBvTTftP5n6QIl5rgGsl4hWWw+Q5z83XlxiUs8+qz1
fopFycA3BxMRLIWit1x/BcttHHaWWiNU/bb8VXf1nW7Az+e11BQaUrJxs/z7eD6P
lMDnZgSJg/zUqoEOyae5TvO5+GY1iOQ4ri6vLArg0YN0JWIrubOGU6/MsS5kvX9D
s4KX2D2XIPw8eereRHI5kRCZdvvTaUwwQzHo2eQi7OJh8vwYsg62+JtPXrej2Q6Z
SpskwN7SGifNWYFgSt/B5Cqp15R5GPkzt8Wva2kPU8E1rpljUT8b64zS3lcnNz8g
8e7AzOugi2kTLCIO3NRAJHUyJ3O7jznT8l/ZYoJGRowsWmAedr6pOjI/imhFp4cj
zSJws+cI1mWFYpho0EYMzol+3LCRCJKgpHdQ3fN+eK9dHG60bW52etEtWxQI4lfP
kKSojtDj7shxtjhaaC75PRiGFS/0XValyGmNNwvpNSLy1wS95yy/0GJGjJV+cSji
m4MSA6fHrvTDtAccK9/jd5uLP+1ug3bOWXH2EFWyjaSZAQ4yj6EamcEYRwixU0X/
ZZpU1o/1HWEVYmAJGiixoQGX709NHBc++Gg300+i/BQU14i3CIP4LfP2tQR9EY6n
zaFziaVoZOvNOOAeoh/8pT1dvZiY2hXA0uQ5/SLo1QzcHXmMe9EJYgKEK63n0XGl
+02WxJL1CeaKHf0eeZTZ4CaVOOrtkdVMWE9Qm9blgTZSZ5n1DIEXsvR0aX8306PX
ncSXyYlwr8EKzxflWPya5qDs9sbBzGa8x3wEn+oEQ8jUOfkcDyKGJ7hQNw5ozpS4
VpFhM9Kp8cQcjF6Jgsjad8DxlWiJjmrAQiOfFYUagUBFL3Hsq2DtSvZgsrmHpR1O
P7EQR1GVG9a+jPZo3rDZFDLEcBszgwp2Fwuah/A/RIXd2JcwQ6sI+Ax2pJkei2Yv
r55+EcpjZdXaDE/HZ4wmRFjrdM4BtB8FvBZdOxHtPJ0nhhA8dnOiqH83c64R/LkF
EOQPcad1X053jNGCDEBipkXvQYvIXuzhy6oCA+7wPTZdaYA8ye66jlM6xq9YRUGK
3oyeGmFAManQL2fStZlDIwL+G2zKSBFpn866KzR95tkkRW7xNoepvzBd6kKfLJjg
+GBwuKiKWO7wLX6yKTCLsUriN+ALSdlSanZGR9KwnwbmesixwQ9lpn6CxUcmd7rC
C0DDMFzrh8c8GgD9MkPUy0it+d38wAt1mT+bzMpdtD9jdw7/IPBvCZ8UO9fsQfw6
iWn2PkDl9Wj1X6kojW8/0yRYfkdjbzNUTq0Elcbww4I3gsazmX9o2KTCWkSG0gLN
Th15JCTtLMEmFdK9rKilhIWja2xaEM88GkQgE3/jIG2t8qEdjKH89sGIKbPKIm//
S8vv6dncCXQgjvJLtgdisPaofBUlRkGafIuW1fVvjvWTIcqsRV96nMNbbc/nPMIT
sMTKKuzL5hjH/k7T/m9/MTeTjFVffv334lXGXrpC5J6wYABa8TZZetDAEpS+eVrn
hQIMQ9tI0s6/pL52XHi/o3Um1chL+ApUfDRZ0UbKxqVqU5pRjS/bWB44+EoVO83r
SPaQbLrIxTaPPWtJPCG4RuBgof7LbqhXYP2e6u3CxtXcgT1J9AQwIbwsbOqRzilX
G/uPQNEKRZKRdvemrNK207Z861YPO3whcp7FA3EfhwV6+fqZzrHEfP89YX8p0BY3
vaPH+xTfudFa8BmUbK3R2zN9iJWOW1oOSRPpdJ+0+DtvydiM4DKTTNFeHpB/paK4
jad7Br5JaoXMOxyBPJpAjvGStugS/ujyB+ow86vXtvzq5SyGHaSYeR47sF9TyIYp
spV8StIliuyS/YyaHxtSYGE8LYGVS2IGYxutDhH9ytOQx2dvYU/YnZk7+fOO0l2I
ojCqfqqaah9vR89sjgWIUcDCdS9/Sf95V3aznhYmpzwc3l+vR7g0qC7r4xwZqQAM
HdZbuWF6/SbUgZ76ubvsm8JXnewdZr5V+LDTisePEG2qPRY1wZTGdefzqFaeRCWF
LMnAl4Jz5peQ7Wh8P2pfLrQLcwmCF6wxqQ7c1S2hWiE8nkP7wVQGhGAduls4kaE+
wMCL3yqzH+E+AUnqnst2fXo5mwPs0Je0/ZD70VM5O/LkUjnZwX92OMbRGXlIkLi6
Z/KgaDbrV9mHcEE48e4VA6QiEpMtEGC68WgSStq9suObtfjMx6PfLCUHOrWl3aYr
qR3G2x6Lo/AgVycFrslW2SfUev94aL2PNypdYG61b0ATOReVbgK7lid7TxxE6xV8
RIgprA0U+Tq7/aNdSGRnV8kL+tmVRQy4qMr4Smgw/j6AavvKr5MjODHvzd6+VM3G
OVAZCNT0MwMLKLl3+eLnAtP0Ncxrv3TH6xmoh9xGT21t1mJ+uwERcJVoYVQ8ERvx
ZIyUmDZEkFareo5dPsCI07EzYNgMPWaGVCN2lndmq9ZmUMOoLoqECNzTsNrpz4Al
OzkwWOfOYb1U9N3AJ2e0tdYNlSiwG1s4JS2l9gYz37AkpxZEq3VdDndXFhq8hFQk
Dfnmc3Lhh9KN95OF2Btf31ubKBmKg3Y9rGGh0FJOEVvtgHEEmflZoW//ivfCCItw
V4Xo+Y2tEI1xJzTgyczSTquN4zcFHQuktmrzzA9gsq9mYtn9A7f6E7J93yBxHKC/
kXyA//TtVCKaTsCPyYZaAruPVDIHyfzTie9z1pxz0mKhFxipUuYaRvPztJNyk2yF
iPuXWGnR4oP6a9Q6TfvdAh7TlkfrUdbeLUqorB5GxD0TsYSRYPRDu2mXJOpFjWiq
8/85/Rx5fmbzDWdEEF7C4hQKQsTodPHOcjprxr4CXUGgfuA4mYZaoLgktjTCqTjb
H2TaV4FzDNfqHxyq4JsEpq6ohjEmCKwSgUOxQwS0jcubPPo9WYibrp6MfcjaCqoz
KtLf1iDCk2dCevImJDasqspDei3nWDq7KsGXee34JLbU+zmDuJmqpK42YB/LTG2x
yRiiHSKXocO/IFSLkc+s8AHo31Jb176yZINPDuY/j24zOnStkycsv0NEMMWmywz7
c93dFhIz3/qTHBBf7p7NtSzo0k+hcjviRP+9KXXIRTe3jpbrvMMREr/HXxae+Xt1
kxSCMKd9NgyMIuGtLKoc0CUmAOUb+IuKawsCmY2w7TiAMaYnglCgiZX1E6KFpc1Y
VHzo+eXD4fgJycDFMLVlXC3MXTsN7/brf6zvJ3+ztDVUgJP2bsoYavH14IT/UziS
vD8ffZd9AqZFzvf1iNGXXxx41rjXHcRFkBBPynoprW3inEXI3fNk6t63NooD5IAM
xnBzVv5YRbRXh3+pxfF/Wg8+TuyJ/WkvEio/k/xG/2EUZTr4ymVXRgG4oXcWSxqH
WY68NaCjJbpUnTBt2W8NC2q+CUcWqFuyf3Dg+2WQa1Pq9NGlsv/nz+ykfjmRWTzT
gQ+W0gaWIyQCvfjotiVsYoHe/qqAAfqRyLpG2r/+TQhcQunqVqh4Jvx/56/Cuy6l
QI2kswr3WLuCtIwTBeHOoaybdZMNfNiKE0FbMh27gYVGtgtR0sGPY10bRRaQW/aU
cO2BhXZjxfd4STP12t8+MD/jZ7rHE/VHtPK7g1JziNHiM18NR0TVyBZBvVvuSVgY
b9ofzXcvp1CjoGwbJlu3wl/Dg7tsXd/45Yi1bp7ZpjPuxsoHuhMrnquidn71pzPN
MZGRgTAiGRqK8g2Ah9ESpBVYmOrHAWTNNcE0EnU0gzcOeft8zXtVBmb2crxE8OZq
y/EmjRqYquzidjRPW+XLZZ6J4eflofK/Ah4pvpFaIpA8O2l+jlFLevuLtRUA8hGv
Ml7E0MaAWT1YdSYdAV6v/XPOD7HtCoDGVBnfjjU/ASbdL7tOLOje8kmOjnoA9T0F
3FLOiKXZufxfovodLEp0+C8V6owh1STDkK5KPoik3WMwivjWZFo7tweCJIQgQzN7
57LBoBsC0RJMEWTsWZ/pcHot5MlPfl68jyc2Zp7ZC8ZGJuGqv7Jl6/NE9AlwwXjf
WUhJ0f5zqF9HsG7/eNCAygRhSqBHHjXcfM+2FdL21nYEDBtxgODFV64bHReXWSSR
qHWfYcxYBXqdEj07t8A4m9soHAsQmg0LljGLhhCDk+hzYKOM3TtIjBgXufGIlsTq
yP2qXqcy9fLoREE8JqotDO07o8u0ipPXR5GM5wmbKQ1eCbSkz5/wmVWup9cJNWC3
cSFyV5XjJtpHyYuHWgL/lAgcBdSCgaQibzfBQYMi4HM2xeu+Gy1VbIcHtFDppFYp
nlzIYpt+Oq5NO1SWnchXOssfYZn4lABFYjen3xuiV9Z91SHjLmtLMWP27ZvO2MUF
mn1XnPoHBx/1k81Tl2pITPQN3aYZ9ZGSbjtS2rvXQNwvXduBt1T9SWRmG2QHXB4i
9rrxlRKZJhyLrsNH5AmLaXVmfF4QCWCF9tTRRBbNcbU3n53Pvx+tFmDcUnTLloGm
J4l/dvFkk1+CXNHjHOi5XFN4/SEAz4AcuTIRsFIyYc0x+MUeLN5ySuP7u+VDshiW
putrXqWo+SDUi/8jsvQJDbTSF0o8UmHwu40jpOlAaOWruVUoP5jKqUHyDa3uZQon
MAEcGYT8LL8Nf/m5oh4HjnZGmBlYFXt7T2nnbBYjk5s8cRVa55WI5d3+QGJ9buLZ
EkpTwT/bd6dhKt8BJ8/H7Owb/GT94lYK1aFCqUF7rFCKkfyUp0N2omr0is7ViC4Q
DIg0YODtd7CkKxXmOTMiVK40ttfCxBiaRgz9kyuL84nHGEVZqUAxS+eDf76dn4vS
12aTAvCHb8uQykaFyVCAoJVCzzUYK6u5qf3EXtLZEaK0aK56vvaC2DXpn2hb7V6H
rthZ+xp2Hsl1yedR5zb+pQkxbnbkKbXq4KaYbrKdl8IakRuH1h9GMaNmgPwXFdJ4
Z9tYEJ/6cKXZcGigZMq2JO8kGQUbcZsVPHgRjJBCkIM3oROYMWZtsTOiWHGdGMpn
N8aQH/jEmbAxcZsoR2z0zUtYHMW1TWHMXoALYZt29EuPbwGouuNdNvMcK5M+T4vv
GFrNz3GKLR6/4A8eoyNNJOEbk2FCAowNRTsa8EW2WMKB9ucdvHH9t2KLpUXcg/3H
zFHUST/iyIDmZRQL35rKyHwVvcTz/LOKVVu+PvpEmi6etFk3MA+r+GE3iT6AKEr/
8yBihfybRie6inlBlS5MQzvGF+cHsbpqek84ujcF/XQavdTBXRaj2oVyRTAYvPXE
wi5QnmfBq8pnkxiIaBnWtN6eobPAPeOzu9+P9MGSSlrqJmKtdjdGwyzdi0aHKIbR
ZEJvocv05zvyDgkV+vOTDgS2fjQEgwXaOQ/4K9MkZHq1Jqvg7N64JB0i05HOBozq
IZLffNcwu65M18CXDTIV/Uj7ny7iCIZcS6/dDdKlKAM49kkuAuzI9UrDCuuGKKuu
Kr1PsST8O4l/1vCDB7yoTKXHOdN12kBKEl6PApCuLuIwnc9zEKyEYB5mLJe8xK6o
72DQFGdkvSB8YK65CnLy6lylS98RgAxzJDjF87QUVdFfX6qqQW4uA/9ArK5fpMSO
+52pBtDQBHl+J8e3B3zd9V/D2rmMRJnRHerGrSJaIL9ZDyaSSwugZ+6oVNZt62GS
/gQ+U+kaqOeaw98rmrgYE/2m+WfwgeHGmVgexx3/SGIqSOffFkRGJNXw70pihwE6
tI3TolH6iyzuU387/CkgtUZPzY114YYNQh0jYD33uVSdOwm/hwddsuEurE2n+K3o
1X7eJSVARsmZmnaWspP+zxLF6+KxPpjAqfY3E3yHfbndCGvGU+viW07LH0AAq5BA
wD/eDr1/aVdR5qjM0ngp9Dk6dSDkXU/SgNTBx/c5TAQytBTydxNFyBbQGvdcpryx
MZTvytvaO1Q/mqs+1Owc89P+7/+ClGeV0SIC93QcZ0w2Ym8tM4/tCYdHjJ/Tlagf
wcL8/AIAd8cs1vJHa6YrQGzmWKg5xD3J813EbSsZpjGrFXEq3BBGEbjHKY7Tyyzk
sGsrw2MBAaJQh8G7rHErUi3NAfUUSpP4dGZdZ8hG/AP0U5ERTur0YOqC3TUdS+ri
F37XabY97xjOENU1OTSJ4FQ1BMC9BMH4brhqVzX6VXaH5hqOzr+5i1l+55kU7eG3
BpVr0BUxMLYgqcSWbbXAtsYBsovyYN6BmpJlNZFaS6zgjeUIAObczuSoKLY+74VT
E8/UsFvIXqDXvwsw5VkQaksaa9nHWYm7J3OVyvku+OTPL6A8kV7UazBzYV3G/uVQ
/zW2++9Nm/SO7fyejfJ93EnU14RZebexZMPU7C6HTdgV7fVaoQVRm0HpdWc/Ft04
iI3/8y1oH20iQQoUFEfj5xpTrcvZtA0kkOGaTIP8nPwMwpakN8tWIaQFkpp1DiGP
Y6rQlovFQNVVfIgk/1jI5sDbG1rSe/zNxQ1N1nD8VcY1/V5k96/BRXtQ5pCU9S7e
CiJVjdnOwShjpuVKcO/5WeIYkLx+zCCKeJ6LhlH+cdQ0C0BaMNTGUVuoZMvLzYej
PbWtmY0pN8NcwW4VePpoiI0oPjvdDpsdXdwTb0y6ftyozY8nOt1DAatIwXAJg424
noxd0AC5KMxT0F46WJnBF5eUkneYqfsIeSsu/BrShK8OEE5zKNC5jtAeqAeGd2j6
vcatNd3s/zBSEidNs70+dgRZSqj00eIiGSRQ9IbfdB1dpm5ION/ODrIULgPGTtxi
ebMy31JzynMxGYuVijbtKM+N1Ri6hViEEV49fLoL9lf9xXhEpudUhI0htuuGgi3R
1qO5TElNgtwXjYM+uoLcauXOVVaA05GNXtu1kJKlONMzegx8/1uQc12gQsYRxham
oR0CYTImhcfo5p+UTJQkeiwCpldJTqowOTGJ1zcOFkgDw+qE73EKCWfTyfIEhl4y
eGj7I+LxqKotPWUN95Y8h3rJ7Pk+QWVdZ/TaehOS+nCZlQy3YGWsDDQ7SHJY1baD
hWQBhPKX++ExkR+qwjoYngIcLm44zlxdVTMzo87NeRBOj26CnmO5Gex/+XzgplzO
AkjtnsokDYO0nqU9eOaeWGh+7Prfw74ut+sln4PdI2b0CaHUmHzWQzg6i+45fa9T
CjwWLy0ZqIzfVdVyaT6WyL3XpvajwiIjOsyCaz0r3Nu6hIo9/ZvNsbk2HQfHXaEj
RweoEbXgTZ+f+5ZsXFxil5VBV1d2TI8KpKoXOozZ+IhHHeCmMYWTzrhq8evHunIK
IOvnd01u+lvSjJ/AnIFoON2xtQQd11m4wqa1N2SDUyjWIs7ibrCvQC+frHXWY+UC
lsW+nmipi9jNrrvxQrSq3uYZ+x5si73Kye+FqKDk5bkrIEugy2wzFd8KWF3pJfJn
wHbXp7pqkLoBlbcF0XVfG00kOwW57A6g5tmg3FtGGr9t2+94/4R7sNdZO3UKj5ov
fV6cKTWXIDMjNTalXwCwrmqByYrQEeEHOxMA4SFmNL/qK9nmaWvRptmF/zpoKBg6
2T9nP8H6LnKDpR9N0aOgO8NCOLFbKkny5izyGB/jjQ6bXn9xQ6p6NqhlzZjW9YqB
eiXLeSKg8zpNPkZRgHfgtYzfuaNva1GsWyUWrKXSaqSmMwlOVE3pI7QWSflcW/lg
ec+MzvQlWcRqUX38shR7T5yinDXFFH7xLUhdVpM6WLwuGGWqhACP5lJ+jsY411SQ
qGKDfrpvxLl6hFDjKQJ4YUn6GIfZduYoosm1GvKXvHSQOm6GNV3+AN5XKpJnJ79d
/UG+oKHmU9IRd2CLym7iYdagOxp7EJwIS4aGmx3z9ek2GKndX5noQEkQGT2RX/a7
zDXFH9tRSleIjbfrncnCWAVRUTlFRM39ahYhZwLQzf5xuD/Cx7bXi5dRf/YqFT2C
DegU5hWlAiDtPY9nUnZkuUyF2LuJkguVgp6VE7Qnk4Sz66tPnx5qxWAKWyng9lAd
qMsM7TPZKTGsV9isuy3oJ5BxDOiWYYYwaDGjTGv4mP3cMXBEqkWGwhPTefgHgB7L
Ue/4iXGXPWDTS1DZQxeXJgLS42L//o+3v7iDRJt1om/I2yCLvs9VjGFy7xbCDCuE
/m5pwAoJL5cIpogjJS3NQNqlgOoUh4dJsg+FtWLGfMWsPJDsZfBF33Q6a/CePKQX
a9A9NZVsQ1bCXK8pYVsp1BpnkW+f/H6IJOKGghl2yVwoDM4nbIE0QTcxLkcKhtNL
bTaWHC/ZAmlc90ZaoBD6Nv2n1pyUAsAJXSnTiLLSxUXAr46Vbk31J2SB81iirIiI
gH90wWLOw3fuEfs3VFyoZsgF9+bplk4L26pzEJYH37PYujuhU+4jM1YvYq8XhmF/
G9Zuu0FI+jZM1+R4V0tP/JDME7P80UzmE2O/JBe1w0aA633NL/PO3IRz8xuEAK2R
LlBuLKHfpgtbt5Xwsd1VDegzlNO34OprLiaZBG7ctIrjuJBVa/xVzNDiaTgwni4K
b4PCyS+tkOOyqsSDr91rqK8KQenO6D7CtpnBcR5iuFAiEusPESxPxI9wpNyRisdL
L/HrMkDvlquHdcdgnYOJA9D+XbYHFMO+q7bZv981BccYlB/7B832T9mIXN3/nF3x
bVykaOgubqtlxpahxD03ykZcnaQLCpYJ7Mx2aqfr4KV0ubvFlRCXM2bFHxMDVpUE
adxwMZ2Hdu8X7ACXJ5eF9O/+4U9WDDAZt351IWBw7T7IhDsTLokcZjT43NTl5CBT
zVH8kgLJPzVrzGGcaufBDlaraFXun0J4KK209PAsJQUi0Zozcbf/PfVfFbHPE0GX
+wDId/WfJ8nSbVi4zMLmuOIiI/D7EdtHOZxbBsJGpzlqq244ddIFaJfgBYluKPjc
cAuGAQoE+kvwS0rcJAyKCExnk5rVIpa2iVKH9DN5h8607s76At3TjmdLw0BwTDP+
lc766W69f65oeYONbFVxoZOuVDqx/sUASW7Cp+VOURd6w0DnANTEoJqWSd71b6zu
p0AMYW4OPDDcffFdVIM+EeGP3ZSmj3X7JjCWUMETKfgJkqBiuL0vb3jVrLw1ImlU
wtoxD5+I5l+vgojMOoodEnrHqZf/yIwD9grPB+/U9Qek5F3BUdV63H9qwsf2GbX5
NV2GDkYRHDZhS3ww3vU+ZxNbrRD3F5N1stOLZMZNDE9DZZ6fv/GiLceAQR2/j2FU
k6DbQqd+lWGU/OgJS3tdGWaWxJc1wF2CHi4wlO0PtaRZY/P01FO284XR8+z8Snkk
OQ9qsgzAX6Yg/vSJ69JyHxbN7g+Ban0WEL1fw7CDyNSHCqjdU4wKjAi8cCFymTrC
GB62jnrh3Z5T3x17WHq5wePsgpBTHOSrYyXdTieY++gJ9daaEf83MrJxmw5HadJv
M10aIBhqBJJVu57wLUrri9FIh1ZsvF/f70Gbo6b7DeKKcLOHcnbyVJOhrt6mcwuP
3MjXDZlTH/NkTFCtZebJWsReCoXOVQ0R70+rlMvUW3uzVo6WK89uLIPp0WOYfav5
g/SH7pn5zIIdT9K20/Cnj8itRUaMMWx/bbBeID8aE88ZWd3nSklgnXt0DSOAtHNq
RJMxIVapDY/ywQwcOj6qchIQ2+2So3VVnugIpLc+FZ4/umhf0o70piIachm/8tWE
xuMYsFtfo0+gHnMbpBW9118GHWNHgLqImdgeMMGwNKGeQNRFbWs8CHDsbh5YfdLv
GBFsqxMuS/2Ic60NoBtUaDn4VNb3N2tZxRQikAhWadGJ2FA1baok71dnJMmB7aH+
YM1vxs9h9jymQpb/tczYxXiXMxTL0oAZHcB5kZWvriWRpVSOK8tvFMkHasMTmk/4
yaHzFEgidROL5Tqtj3//ExvfExi15txT+3XhmZ3L/eYblTS5sYcaItvkWN9Iemvj
Q9bIjDdeFPNUmkz92LpJ1tF6dpe8Kx8cJgPqMmRwgSiYftnbkkutPuEJo2OI6pkV
OCB0rJEeepafxEzXFJnDgIBuDJR+jt4Y+FL+FChhj4Wbudzt8Elg1a+kR6wh/kfL
CZ7SoEO8ghxMuRJkvSAUjesWt2OtX+h4JY50rkPf+1q7BfZYrNNbqySlfPtu8id5
294K665ti/+7hHfyUMmz1M1bMJVgOT8i4fPn+FbuVKGCY5UJYqX0pANSsh+bCoNF
vqa97MCYyPhdUh4ipHxFfvTPA9nIK8zEusgKlOjP6JG1HEUebNcgEq2Qzz5JQWP6
jDxLCYwwRowWjEhdpDLxuwQkUZEJjwrE3hDVKwnOGe5Lc7rK9DgpIRoI3yG+E9r/
kSfOFq6UtjInoW2WrmNfEtjWPSLgwFhMSWGMuJcAqVKXqMp2jDgmf7PEpAVut6Lt
6o1x8qvytM9GXN4zMCiSi95FgIt5XmlqgX+CMeNIKpysiq4tHjrdlp48i3lOmmSv
OGd5UEBnoEtbb+9gS9x+lC3Nf6u69Lb8/dxRci1fbKYU03je3JC7SQJWL0BITs6V
mNIj6n3IaOPr0+ToFQVDcbiYYJByKtet6KMvoek8/840ecYszXB5WWF/im1pS9KE
C+1FbtYbROt0NmP5A6erFlNwMMJoBW8mTU8WhgvWzUKA0+mR8fgHkYEmlU5K3cTZ
Xh4epi4bMvNsvrVFQ++8x0wLtn/LeHOWWOKXzgt/56VaefnufYMqGFJkJJvdT0kv
2O1/CPe74kGZUajriKTfI8EmP3vnVVKgnjPcVX4sSvPRRA1W4/lBzkouEAs4JA5e
34hMxse3WMoVrC2AR0mqgRIPK5DKohgmraAoeD5g+Zp7mZs0tSo5pPUI7PLFIgeg
FGrEK3nE5v0ryFkNlOWiiiCZbn6tzUrgWxtzAYox8t78SBR8CxvZXIPMzrL8xMiG
YuYO2Y9HkrvqIfN4xbkjf1+Jl/UL4tNibhzJltFGbq/O8qJu1UhINhPPftyLxgzc
d07Ac8EZlmVJWjJZjre6IpCsVJqcOAreUPBKq+yUPet1VSZhC4WZyI1tkyVC//Oz
NhRYZgicw+7aA2Dgeya+sQmL2pzoiWHnqbcyySOP1j533r2GiUvpSRNIeMUtYOOe
XwIB+HTomrH4TZQJGSl8/j7vMJJQfUBH7ijejEp1tzWLY1wgZ9au30DIHeWAp/Kw
rwYlh4wtuVKZ9vzxkCtiX01w5EO4BUSJgsdVqnTsLOX45k6UosIFffYSdmCH+GKk
ePSxmsMhH7Bj8XLLTy3rcVOjLPbWBMflAGlwhylEI7G88hToOHaoB3N0mCHR1khg
9nhIPAVrmQxqrslW+RQQc+SzL50R3hHhgRX5HnvtyEe1pcDdrX3aAXd2vit18zTx
Vr+CjfexHMAzizTwlZ/ln5yP7X/gDsfOXjewP+GyRwwYNlE+vOclrIjJjbNJrBqj
QFIJ11SIzP2HY2N0J/E/ya0dy0hajPovApHfA9jizCGr+zp6Ma96VRXJ1Wqn7IWA
wblCIjNLOqn1GCfIdGXmSYeJfGyyFKvAxKp3xzNkZVguIcL96IUJ86Su3t8lW2DA
hQWFvmOoVZhr0zc1X0G/AjeeaTkUXjk8HhYih9hsn/HlCZPfua1gIyNk0GUxezNS
vYCST+Nsa1ORThIJdWhkwePVnsq5TmQHqwFCuSUbJ7/09wAnttJgpAkx1SOiiqd7
BYtbkyA0ZP/dpzLkaU+Njb2PrI7aReSpm/1UzsI7xZJWfsdr/p6QIpx5k8mTMoAI
FnyWGWTMijSSRo3axWUt2octkc0P1On/uA4B3eiCcRBdJAHr2s47q4ZAIZYZFOL7
iKFEEIrbI3Og2IwXSXyYlkoyiqN2F5uNF/R/2SRCQLz+6bIeUDW/yAVDpmbGtcjH
7hkUEbzst95rtP6RdezUwJhHDT8hpBLGEl4Pvz9hvWU7PE19CwvS4y16MTkdlRdc
XqSKGQgcbhm4n5GkhGw3Eo1ZWcfusjUPUI1Y3aDfXhnYJUos05qVaml35acuiADR
1Z2dtfBRtDADA2OZtyW1rmhfLr0PS5bmwIU675+waD5XzzJfKOey8DVRtwk7ozor
i5CRKq/cw6z7nYmuXikIpRx5t03tO6HqkJxXhp37NEQBaHbJjsIRYfA6UXa4MWmT
ZgMOUjFqWsVAhI9QPeF2WzS5weTiTb+bEhPCOoXfwus2BJgOPcjyMKYr4wY7vchb
bfUTwZeJl/Dr30WhMs79Hc1+ItHhYt+wXTRTE5DcXQqLq5bfQSnXa1PTH3+ETd4b
Wxa/evWYkf0AZdioj1uIVD1XrAK0a3Ki1/jkeWI84kTT7czZu6F7UIsVTE1kHOxQ
3kFsSRyumY3hSdDCowpZhbLvHzaS+V0U+KwHml0SUdT/vGxVC6mKc3yCl7SkY2ki
k6QjfsAU2Pu+QSWdwr3/zmbA3JUZECcRQBNF0cgh6C9brqJYAxHLisuTgumk41qS
DsD5UVtzuTIcVmG8lWVFQzbUSp5PsAIYey6FNmxbyd20fpxDDnox6cGFplIRMR4d
XqUp/wyNJITaFQF8lJfsad6bl4rulcVMTujB9hczh2CpdgLpOW8rJfTcO+laBfTF
OoOEqajPodZ6uhpEzqrl+31T/dRxqg0yF/4wozrb2QSKawsZBukEGRjt0Gm09NF+
2WBxgHmQc40+s5UR0aPmv7pggUUY2v0no1c0WfxY/icSGSQATMZ8ZS9x0hRwJQHa
q9boMYgvMX3G0gJzJ9q8T+ugwTpEo+DWa8Okvr0lIZskx+1LWdapA4GPxf18YgyJ
y3mjz2IEmv4UTzh2oBm5rbFvPTh8Eh7LnXazbGCINwMCO2kLeIsp6jGStg9afxEC
IQ5KLglpe3ZheYs/y+coMAj8ce2eeCdmTLK61QA4qZdHwuZ2Gz6C3y4BW7nsYAej
R5MmXspsSkHfb2d9HFb1P7UVzzdq4LK2eJrXfOlFTbfyl5N4eRSYgHkw7tsmsAO9
98gm1GlJbqPm4iTqMP+I7iSFt4GWZ/J9MIX9D3AjiG3DeorWCaMeU/79CSQhf9kJ
hCMHDeFbZD+gzUpnBm7os0SL5bi35iAYNl9t6KVA0z+2fEc0NgnfxvlnJA86hWZY
KbluEFscmrfk/6KawMMG+PLYE40W+gtMrEVQxxCJmPjTIkUdbawSTPDV1JLYdhwk
VR9wOaO7g/9nv3dd3+3hRGahVk1aKHABZMCjsVSLHZOtIfmsi9YaiWSMB6BAYN8m
QCJ66f0sUDNmWJvsI6KNf3aNwuznESpk+WWyKm2ZNx1OEde6tvYlGx4+/8iSg5kB
EysNKwFzTOzGsjvw+yis59fy3Dm8rXgvmxHDPaGoQUvEiPVo+LDFdgIcTkGvWeAs
0PUxB37HgxRQ4bq46L7otzgwCqBXdGfJG3FjriQTtnhlbnYsMVoXtzS1Ylkr6JgW
jVxvJfkXwVDuqwX5biaEMViujB2/zDb5GAWytIG1W2OcCOgTrrLKLbREDs4+BQg8
Z98cc3m1gByXWwunNUrLaCKomQ75Glsh4cfbbGhTTJPTVeUWfS9CX6xxtUfCfH8c
oK+ne0f72T9CS2lSghr5n34BVe+9pFtavxq7TObFTQRvVG+ulE8ksgcgOxY0JlQr
hMxPE1RXA4quL3rZD8YBIzgJuQUEmy5R6HaUN6vgMkJnss5h0y13c/5Mn9SOk9Fc
ZPwU1MuGfAekqW9wq+ESsBpKhAMaeCZmFNRk4dTYKyHbsYbV+NoNsbVmOQmUlqSG
+dKWQxzX38QgSJt+APiw2887UENCk1nrHdmHdueSmxFc3OBmTAMHBuf9n5AxRTvs
rw18bxkhEIMaZzxAjyvCVqeekmwmy5GbCoATlGyDt5UFC27k3Ezpnk9YYXoPscib
08yTICZgBhNO4CwRxQj8nW0Q0uQoyWdd0Mss/X4EzLyT68aj14Qf1y63p1+aZ5m8
pjXVa+ie+qUiH3p5cLeKv1I1XrEpcnHMrMJQsnOBlsnjyMxi05eP7MsE9huAiWup
cWsFLJEb5yCWC//5nU4WnH+imTlSzQLh/oPxjbkV+LpaEOXzdJeNMrmFJVFvouKX
VsNchMcXpOERsG2LIKy3ViH91k/2toMmMQjo9IxsAxJvA3dsc6iHkDG7UNKiKc5O
/HFySjklgYZ04dpZAnjNOQ9YJ0tDGiBxc2pw2W0XbN9i5cfwDHzyQ7Rr+104igAm
yDA/Vdo7WghIOpr367Fs0ee0p0DBrlQfCNnfEmZsYZqGSZrABvRygiJe/stuTpE0
E1FPMn8uV32UpCUOUJidju6ZBZuefAMTyzgeIIxdDtAi/JKG+rcq9WOerdqLxL7y
h8PNEvutzcNXZ/CfcHWXFLtFpvLPG7uURxuclE7XYpVG8xE7OwHKcAXaqp40MPZ3
Cs++Q/xIX6UVCWDSioMjXKSG/mSTmDzXdDMTqs7r9UFHOEuQBJwP/p0ANZW2wexn
lMQg+FunfOQUQFLi1FK6o1WfrmmS1v0Bx6VOP1KVoVIyGOPPR4lqLN7q1CTF0Gd9
FeP+29tPHQPiyWW55MxxDHLGA19FBiCTnSX8S7CebR6VqHwyGGkAm5I/tBqjg9gk
JCv75gMch2yqJWxlL/03jpsRF2upHIX029f3e8Kj2MoqLP7ikqi+mJMn0UE8igVE
6RQDqFtospeeHQvTz1pAgqiyNwcmGOZGFjzYDX85gQqb39DhOEjHtwx90jnhLFKp
MwP592tZaqxMapUG7ZXXSYo3iRVYMaEUPTc9JueE8/I/qMN0FItyMzzqmKzER84L
oun+IEMg8TVpat79KU0d2fnwK4is8ZmcF2eRF3dyfwrghbVS+vrj8jEKktH+Rwdz
/db1bDpFT131J3UHtrNy1qyTBV/KwrUxh345456YzpJRYJPsTxXQjqfNqAeIveZC
WlH/Dy1b0Lx86w+LiuBq+jzOgvymvnwweAJMjnarhu606f0/OduLN11U0bRWct4I
lJQKfnwKtyJzyyzvtGguRXvbSGd2qUGYvMeN8/l1UPvqSF4vFXRJEQtuoAyaM4Tj
lA3kPxl0kuttR2iVvvAVQ2d2Mbitq7vnPSXG6QFTNxRsNseGngt8n/cUbXoH6YN8
DBTMl8n8BWg9cBAAY/8IkOWUUxp5XHJXEE0QSTcXcenAMLkrn78kmoLEq5+aIgdg
tz8nEaFeWaWEbVXsPYfAptOWLtR/CPxu4+T1AhqXhSTB7vwRlTQ5mSRMKn9grDtl
lFXnzWgTwfPEtL3Nyb5BApbaXT3fjJ8YS1D1XUyUL0oZ7ZRGG3RvHFcxN4uvYYtu
wUOgr2CyJgRhDB60TsIw411cE0Mn5h8PguHXMpnlGR67Gf/35RDiMqTfXLB2AIbM
LVmxfqRb+khYniDd5/To+Lq6LogcyEXGKxP+3PRCjcKpPHAvPKjBE1LdJccT11EM
WMXNk8c0A/oqFwZmMQDcVCuHBLGMCJ9z0Zlji/mVQ8avgWGxzxWnyZeLRTTFEApR
1QlyXl04ARL1fkF1XrxzFF+4UvMwkUrpEgQHbvO1Rr7+h18ddb6YqKxD20UPBZxr
NkJRa+xcRgEDk/tN5iAmZK3GC3595T/untmUC0Dqpf8YaFmQ6MhVsUL8ITrFxA/i
PDziqYNnb+MQvFgv7RUqK1PrkFlIbxErhhB3NYqhgJ1ZuoriL9EMyZ+qpHutAME2
R8/abD+I/Kng8eBrqRHgyKxlipMzw73/Mr4tj18hT9oKbk5RyPA+1vRV+0C6JlNx
w5aRQAzi5K10Hfm4Fjc5gu03+VgDKnVYatJKVFsvr2CLFo1hVYWCpG4sXB83VWmn
Q7rMhGYP/wEtRVviYuMGis8gVU4tPDWhClTFfBCN49f3wlqqgKVhxLYi9RF+LqWS
DSLtbRbv/5JyBAzG5HcDnUOOngyrWVqgSSIwo6+/I76myx1ZpDBZFCKSNX+/qBor
kSTcANSecOw0LwxQ9mfHhUZ7/CAdoaIYysgpGVwG4OlY0lf08ya6ZAL6oqSeu09+
VE2K0hjpRGSDeVtx2l0gDnnm5XsHX+6EBUKSpnX59+JgAr0336vh0gwwkdV2+K41
f1uHJ4wkFKdLcPSH9vj1F52G9qW5XPC/+fM5ALsdSeAos/GgWj+AFSYOJtwCeawW
yWUmwiXG1YfnKZoF5sfGYngx7cMcDLnQIJ8SsPq383T93TKyajAj+wgV7KKx/8Jl
tWADiDfqnEJhgXVWRKyzyQ9acgWYGY/DHVDfELh3cyga42L44fw9b0CvcQEIv53p
pBMWc2fSg0lZXegh+d739580AM8C+VHKT/pcAJ+fpxndrKFYk6hAEb66JPUL5pQs
iTCDlic285yg9b2maS6sJh1YvFUtthRk5u8MAKdt9yv/8sciL101gq9q8fp1WYH5
dlRVjmmiDo+gZJtP5DPCbGICgew2M/iVEUdkzOiqpgUnut+puJRLKKxlO3irAxu8
zU+hC8OVo+Zt6jUMF5p65nsuoKL/oGQNemU7bxIliAXE2mlzWzknsZMMStZwj1Dg
m3rrWuGG3YPczMfuU7YqYEwmo5S9FTSamUWVDGXLs8a+HGf+2vfZkxt4b+Gbxra8
2hLJ2zpeotn/+jMmxS/K+CDxLwYr7RcvIV08zwP2PvgkqSRAKa57k4fwQQhHEXjs
PNNuqqVQ8oqpVNpuhLFvS1a/Rlh6Qmle+TfbiSIXz8aal4mZBH6oe1JrbZZv9Qon
ngVLoeUBWS99bWkq1O28KZOnOZ0ZjyAHRNt9SfT1sPYmcVQ+/WHK5fWgFEaZ5h4n
1sqj6gR1KnQA35Cl0CVHgt/ag2PqsTHvkB8vvKZteANjIsfsOIbwdSAf3tiTKoo5
drNARIJABmnK6HSi48CSef2UjN4V8vODa3pi/QbNg2Dlp/dXVQ59BpHDKkybamYk
3G2zwKb88e+vK/rtts1caFYvNCx+PZOpum4S0xYCnMzoqCKlDTIlcNB9aV183Qf9
O94sSbBZBe9mkPspT79lQLoMv70go6Za9WAtB08m/+55AonNYZIXL9y7WFydI9Lk
jlMjjKIMIR2VtZU33rPo0x6zmWag5CzvnZKYKkw+6L/stcxWvmy+KFVjk/n8SpgL
eZSET0pBqn8YI7MwuRNjR60KUz4sX/Sa1tAG/O0tj5N3KjuUPanNxdzUMLZL78UN
DjIM8P+bPljv1iFTLyj+n7cP+N1XXI9BKXca3UwjA/sNsV0ec3DqpZPduOBJ3Ipr
Xmu410nbVmAGlDntsXkVgUXPlWd2FxrJyEHpE+OvRcizF+X2GwwCZcQN/mDuuFfY
rSmJD//yS0yHf4GShmGbHult30B8dvkeW0vfK5xFTjnPtYqXCpJRycEfYX+tGSsX
X/jg3jZ1HFwbA0Cb+LxuzV4JKAUO+Nyx1ikQM9dPE81axQ1haj68CdV3k5o2V932
skWzNULF1yl2SnNMW6cA8Wo+Gn7Che/3DAsoEawkHaMvxLzZwzmmNraqZUnQVurI
TRgzlt/4GQE0LHjuOvD3jwU04Raow9qgQb3m03LkWr+jJ0KKF6cwKa2zZja/ePee
X4l58uEIODZwRUk8orfWPRcvbo+PLIj+Q3Oh3e0Xc5OxpO85JLuYt0JRFRaTG4Me
cAMRN2ru0bUksDFW4B5VIRL/K9fVQntcOxt+bjwBRVIUwgC8ujMezwsuKH6pvlhj
6xPGPPaDAvy+/ohoN2USh3AFlkm8XZ5vcPizQX6fzrSjiHmXPtW96M++70+mMSvu
aeZIjA8ypyMFD3k1H7UO3n+K+/mTkpAtLpftoQnby5QKtNQmjydEJakq36jz5002
wTHwDAu4tZbNXJMrqIpQG26VMxX1L/0nZlYl5XtkMNBV0n1IgU63EZunWPdnQFmE
NJYztXw0WYkJPfnZL6pWGpfYkiA5ritIVpD1fIkRNETDlkxJOtm1y4JWN84dIBJF
alEsf0dK7hUYSCBxfJTx8QhRGcS5+xC9nBCbefKGNDUWrEXMn77SXPnA1+SoMkVZ
cGVriUFXxmZ4ny080AUejnsc3wAXa8KTampfWUDxK2hZxagQNFykzJlRuzYPbiXq
hdg9Lbqbe3PkZfxiW6JwRKQMQCCe2db5yKhYA6EQ5ba12lqrSCN4OffNgQ7ZDIsn
gKGW0Wqth/NhPu7Fj9hvQXr84/BdvQuKtjyXoiYG9pYhlRBQLLdziLqwZozW/yFt
8dkTvxPMVDohAuQWeXeriL8eyi3DF/kiHq7s6V3ESYWVtG5cKAUKhyVUqkvrpSsY
+gYE9dOnYc8oGwesw4O0+RdWaLq2BuSmZeaLEuY9IX8R+YSm5KagK8GJ6sIav0bn
amiY2Mg66c5SQFziWLs/vYpJyvX5bdE6w+OYaSoRlLervt429Tzhlxjs9uEuG6ky
uyLf6mA1DRAWyuT30EhPijfCeISc9M8QmAKBdq4r+vuox8PepZenpTCsC3jdYHLK
E3z3MaRk5lhYxKnl13vM9yxcsJ06RxzHYUImx/bUJpOPXLeDSlydmXMl0RNhD4bX
ZHiYNFFD7UwYp9FqiOhCWxU3PNqcmlnHupMlMcSY/iz0uzhxb+9C0Ez44DAizWee
7PvPOVCGVPhZTM5CrmhRkay/1gTyrAYsF71hsvIEePvD3d6ycvzV7pbCPkypl4CU
dlatonRHJQi/CVC+HMk17uhxrP9S1I3suOuqnGg5wYTaK8aRWFEVpd+jhRN5zqUn
xB5ia5urj2JfkrcwIDbEZv/STvnIHM63pivWHZnee/ed43NONWnf74EBwAlKjZim
XW2FwhFqx8PvM1nxvWAOVKby1EposIwrvUFMYyPECavxAbmgA1jG7aVRVCVMsvUd
9FgMwqKUIkgGTIXB1pRI24jpKIrtofVZx1AfbVwitQs6YhiE76XRI8UiGjqcBfeR
r70vt9nXmoMC5VZnCIiHMb7VZ2cX7QrDtGiFGak71sdSjDmgcC5Q/ItFB0IfdChF
ze/dA8rOWA7Cao2xOKYUrdmtbWcq3wLHSyQO/vBwehVpH9xvfjh9VgDxVKiEK6JR
jAru9od9hVmZJe9lWi+6Jbdjhn3JCv9xecFhCUaiMH/Oy8YP2GSX5X178w6opWAU
m5DBZUkf80A5X/9SzRZvXGy0fl6DdVD1wo/wdj6lyvWhCYqP8yT0yLEHlbkK4iLz
3Rr4nJpFc0v46VlefSiEhjaCyew/VTqf8pd+gMQZsC8OQ06OyrMKtDW7zfzZjuiu
+CJpNqE0XJ5IeRSCJrRJ/HUcuYG8MMbvsKvjYNEK/kAxJw1RNkSKHDF7YFW6Wsug
2RT3X9A+/jQKY0s11mz3MkFKg3iAeFKnkZZsRnCgner0ffH0qbfOmwlqJuqXLhje
GQNsKE9DZmuaVn8iF2NH2iCZaXaYp2LJIx35PxCfvHnXGUaV2nBCGYS/K1txkLDC
ti+g3yCdhP0a9lnkF8cDCHzGBnkdkbwY4ftqPw2ddr6cftCq+d3AqxxsVhk5Rmsk
nalCHBwQF2ttqOObP9vJ5LY3QXfOxW/qSCIlOr8rAIym4KIXQT60ZGGq7BOzbb7k
T++Ctf8Hua06r6vuXquQD4LMwmrPp6jLINcMMtLnikps0dfV5mTBjxytITLQ/f+F
dOcoTsPVESmTS5Q1EBxE0+JLJdhT0L9CH/JuEJy/dpPWX3oy6EsjT3FRmcW5H7Yr
9CxhJnodpfFCnnRc7lOQSudHnewVXe8PSmBQmeKlAeTHUSzOIv8DPNMBkipWlmvP
CB5ezPwrR/dDiSC4rqyIc8c3zdl7jGsHBSR9/DyK27vtD2a3pZ+7Y1IiqtIze58I
APN9kzf8POPY01iSzpHuGfkCbotJ1+Zx9REHmbVGhLezEUdTNWqFlQkAnO7XI8U1
eRpm12IZupR2dMptN7r8gqxc25CvBBrNCW2yC6BjJofjVufLA6YLlrPfDBUxNcyE
i6H+EwIpExhFax4A0jRq6MG9KWyQOp+CYNH383A0jlTwQLQI5LvlmQG1A8kBEa7O
J6UNNLRhl/3XW6uW5NYZIHrFQcA4QosvzLw8pK6etR85wI4Q7ahiOEkoU5F4jeXt
LsFbh4duapQ9rEr5Z3IeNEz2+43rLFC9i8kTVK5hYES4TrVgBUphjTQPAGfFLrM3
DjbAR2qur9ufdRvXi7SQI7jzYjUGgAUgaVEyttHO/e8izDsEEqwQ3OUDuUlQQgs7
GGbTfh6jZ4YZJQJDHwPPb7bNz/6i2uBkwg20xwL2WSvXPZ2MQhnYHMwDN9gw0xKz
hW+JmOLXunEYQakFVgyNFZ9gId0j/fEre/wH266Q/kRyvgs0DQ1K0Cb+9NZ92ApQ
XG73K0Nm3qEKckfm+VwhEOHNYDBvyen4iSCi2d3iEI6+nBBkVVB0yO9vNBXFc+cw
ICPvaWNUrfpJ5948qlrhIg2wrNgBu7ghnYXeqM6EfKG2etua6LlORp2eVb62YpY6
SHgVN1wb4Q3fNV83lz7iduvBWKRb+1eY2jn/yu8v17bgRiOhWALJrUVt4MQNZTF0
j/YGzoG0iv1NuSJ/2WoZwoAU1z5AeLNmbc9NIKDLE3kx5aB+LlxiM4Yejzyw5uJN
GUIfHTHVf7PA0ZLdR3tXka9YJjk6zfaoAPvKkQM2LYY4wc1S80gkwMSrVonlZd+E
Mpt0i0+DD9xN+q7WuEmohNxOOkxAyErfpDCANMwPKWsvemEkustfuCFPVrNxJoXU
7uLA3FJn+oZxw2k731vXRUS7rNz6eHkjY0WxGUIhAqlLlUlVbkFcMX9itjVw4iQI
1WBg13lzEhwS2ulKe4K9N50cbBn3xY0GduYO8oCiV5Z26Dwjui0d/5b1zKiQnChY
0bUOfppwGJcL4EDXWLcTrwWmCtUfyfFWpZI0Wx9wLat3feCjzNZ1WAl8gVzBuPPs
qucU7Y/GzWmFM5mYFscfNL3MvRpdg5bhUCbD2g4Rldm6DqL+jrLGNshbDdf2rtwZ
YZ+R/F+EOdePLw50mRZbnotiDK4NhSa/oYo3eSOYPRRsJGPEKJb+Ihk2hH/7prav
TEhnA7gGa4JQXtPmJhywV77jCZtrracFoYwqkaUoENbR6zaJKCGEXFQUiBomKkVP
B7rNt8N0o7ZSACB8e6QHAdP1j21l5/LxoaaZbGVQ5mGLnDq8z+1PDE/jk/wFOojF
kK6alHorLTNvCV5BRr1/Iry1dadWWLYZmVlsSmCutE7orPwEPpL51ft5Hb7x4awc
LDpPYzrEXretVFWv2hLqwkHjmU2l/rwd+daS9QC06tjumgWPcxIvbPZoxxzCxj+N
vqtErR/zcoHZyoePictBY0AHNUFqDJjHRxNR6L4+K6B0unjRdfCPU4e97qrUSy8r
eCA8kjZxgjI54WO8dy7XOrud9E6IBJsUZUlw5DVC8vXp2cQveZKotA+cng2XNOxa
z0zK79lxW8v19jCTO34pF9yYM3ZMXfkdJuxtnfbQ/BkSk8vaZUUC/VEXdg4YvHiz
DVUJ97YCntDUZD9jmtpgKXOkUu9kXE9sSZUWRVXVMbHHmPOZJ+KS6GpXAMYH9tKt
VXe+ScKaRt3jQ+Zj1/NqvqVjJRKm5V69zI0V9hQA3KzQnRR/88ZDEK7qJ/2xXmLP
wp1uitmUrYKFgM3J1hMb4/I0DA0J+5VLlMmHQmXJFuVqeskoTBAiBuBNlYp5qR4V
XwYw1xeE38bI0hy0VJxSxonaXQRzxI5CgGWkfJTHQv393nn2QlYH02vDxu0qctk3
SOWVG9uxqJPH4zS3s2/3zcGD6O5C8HjiM19wForfn37PxbJn5fchIuw45GPsdjXM
E/8y/EJHwf83/2TUt6CeBY/eSVtW8JYFOCxG7GnX/72G6gshK13MCJSiKUJcXJAb
mHSgeNVMrhEsNaQexJxL67BynMRuGLQ4IO5WxZ4gD4R8f03Q5CBCosUnXKSmvGlb
b/DLia4xUYhdRU3tsc1j+jkJeUj6dYd/AdSyMDheILDEiI3qlZl30tKzTVyugdJC
KzTW751AQU3GtplUAiahfjhxB9oV/eELTT+P9zNnKSbSIHCb4r1Dh9wEkohsZi5/
AjPNAmDsb1iBfqmj0THgUvemtUinTQyJKlANhNAeJbtR7loJWYdcXCoHzZzRtvv5
1Nfhd3aH241e+leGvwrxV2oHyrSRAuuu78GNlmV2Fv+GT9raOSqhv9Ky/Xn9L0GG
nKjhOteb0/kUnOYg+Dhc7NK3QTUQ/xVqkozhgA2SidFhC9CeXv1GNLOYHB17sDrK
fUT+JxS01uW9Bk1doXGa9f+NhqYgOQIf3DSgtcGctLORHzBTn8VzljzaqSfBKUKV
rdJcMqJAIwEXAZoIsU/BAkyZWECZiE8rvLd52h9xWnmdwWgRuvcaHZILp8CzPQLF
zxdcbNPk8kucvIO01xIbk6H+U0lC5LWvxgjr3i/St3KjSs8CAEBdvlrqo3/oXig/
CfYnfG0Q6JXlLm8bXUBTCl+QZN5bsZ9uySJye7bo+6PWhQ8U0+9XZiRhHJ+Gk8LB
iI1aRkg4JZWts3dBolA4zLbEjpN0Zc+tWvSiG0AUhzxswa2uXzEok5a/f2rtN39U
FtKx04tCz9WVD29EGolbG1GVmrx3+N4shAguoI8919O9IDJj2VwIS8oBI0LQT7DR
d/JqBKX9wsXvS28bEECsyiiOid5TDwQF+icSmiPo+/lD5rurr5/4FCWBColL+FBd
uuXMjzxZyvJsK1jGSePoK1NaEjo0cJ4eiFakx98+EWt9bj+kgm2c0nW8AM+r68Ps
H+GeMC9175Z+N6s8FRsgRjtKLKRe+PuyPWy3KMdOlX8f0Pd9uZWrTtDmcKSZ7d+6
+bQzUwt2DGE9OXk0S6ZAkBkp1S6iU2/24I6KzbT01ogW07nt9cLYu7HlrXOUucKp
HWQQWZLO/0h2nOyCOpIBnqjjGmMmpS4noiqyD+wQxqGm7NxIIvkUbNcpYCyFTt9d
EgCRJGSsbNpSo11M84gadYbJ3CT+r7qesbppjNpfsVjSVRSgvhj2iV3bBnSzswZ6
N7ZIkRw9fXUH1j2vDQcra1OoMsmcCPQ5JX3eSsfMO3oBjYPQtvMkU9aLNmmSPrD+
0hlDgHWV2AIJmo6ciYXGpuKkzMyWVAOd8hTlFt/pPnnS9PFITL4z+VxSxB6Axi7d
zLl1RkofQtYf4WnrhY4iUrq0iH8TVCK7uVLZYqeQRsdg7nxI1+gYxOdTOBlqbHjB
tgYearOi2iFRFf5BIxsFnnoRojGcYaK2b1QJIZjeyDnHFSf4gpwUOdp8YokBicMB
irl5Hhm3Q74xk4x2xSpofQEiz6r+WHVRSCw892T1ab0qVU9dy4jdhAe3dUg/0sws
DK+BJ2KvTCl0uthxYhI4NBwCLCKgUBgBkwqk2oXoDAQkrvke+OppI4GyAWsuBE7D
EWghILsDG7rKYiLp2FZE/X0NXxlEipIZKWU83HRtyHDQEptaNPUDHDb1mdIEwz4v
1G2wb6xM/IXRqB1/5l8vMh5VbMEH6RNDMZ2dMTrlVyo81AN2tflO/ERg/S92H0o4
tL3wreYEqgxgH/89W8QCB6Sl1WgaLiv9UB4ImYYHcWpVuybKTo8okyjPO+mWy5Y6
Z1+mjT7kAfnih5lcJ7LprLKbX1ykCjkPctnaCA5bYQ0CsZuFp7U7HIRjoF+K/Mlz
DiI7qUC+Ix+uZbX+b87R5QhmkgGKlHQeIbSvFFlPnsklpkD3w1txKLYKg+ow0MxX
hRDs9dV1ioirJoTOxz7Zp/c/aJT3dzLEpFP5HUkscBoDyptbJJQNXr2Lwmvh9xuX
KbFYL0MOwVKt9NBWWKclh/WOXzlc/EhvWu8YCw9sWimncgJ2vCxSHP9H+/Vf6XBN
0u8dNaj8ynnF/jI/m5eINTEAD/EKUrBtRMtZb04p/zdKXksLoCMD5zA63n37jLp9
odxl7Mo4RMJLD75TOkqQpWUlXYJxeONvCPIBJC2IvgysJR9fgS1xw+Oip/jt+pg7
vV966LC6kcJbXLdUfNItCR0X5kXJJsO+TrO7EDE81LdsCsepOF8c0VvlBS6mYYWv
pUnSaTNaWD1P7l9YYywdVkDQdeAuMJyhiZmcEv+nfg/PXo9cM/lDMOdYOl3S2O1a
mCld2JxQ0/coQX5VroWy97tluyiCeCQ95+9aOmhjPwHQWk8SA44z0BgOIiwMIsIO
MUNw5t9VtCdHHligmfRLPo952R0pzKC5ZUgwfRqNoylQL+8Mg+qHn0oM2kLEqGEc
UdiE0bgqXNWak3SkHD7MCTHWgd9kIQA10lW2XKz4mfCjc/HgVZ/LWqMzSklAoPes
gyaHpLh7l4TLsPElQWOOlvtzLZeSlPn+0CP5dFZD63MRqkL0y7uDPZ/ikixPXhgY
zFXP6uLw36rnoCNprD7BDNCkZvxSfp0amHCkSgb1G25v9NKoPc50TRE3+fJd+bAO
Hd3JRw+ntZ/inH3w/sN+LTneauPP3Xu6vIZPZUhJjPrBbmThynp1ApYbGsFpNh2X
3oiu1AQAQb+/+lAb9SbDXJoIOo0VPcTXKWB1kwPlMufLeSwreCB0QZ8Gw7OD9Kms
w8H38KUVrR19XSRqEQkO5a5Kz3TKMCLy+vlLwcLkxIkmfrsokSoiXUvcR7EpcuBT
8UUFOQ7E8PFreYq9WBEbz8R3zJsdzfMg6ErghkkCmIAgRlJuvZf7GJIy6AYvDXqh
Fy3FJPvXuqKf5nLeoaysZQmPlf3pPc2PPcgWk79q+QLHa3U9gyUVJ5/fcuqku7Nj
SxqmPb10L/Dnt4UQxBaRWFL3/YElWylwncad6QDWSM0RoZyuBO0KIWPUfDjASizw
qwoqs+e5L/b06DSFtYTmwXo1G5cAJTNn6hDFDmnkEjfHTCirRkGPkchVNE29jPBo
LdunFO/GT0oh9NOdNjKYK1gCvyR9+v9fy4GL0TFhx30D0a6qZ8+DjOjFD0/28m47
HPzH54j51gmxhPT/LI2sdRZ+8vgowSRg/2w9WRZ9Rx+qm+qsAidOM0Gvahf5NQ3n
Iwpa10o1WMWxWYJrTQYxxqsybyBO6NX3cLGpBQp7a34aiEouypkpJqQ/g2wkYw9p
PsShxw9NlRvrBPd2DYfU5N2K+CeCsiMtlYFHlb7fHQcBu6hQt06+exeLfVCpYru3
LP9CGorSrF/T8xrzBNcct9P5e//4yIGrw9VGMoTev3VSwAv4+UWuDTYWUlSYSiDJ
Kaarh3N6gwoaXa3W2cuI/+KDC2TNo62dMYmmdFvVlQ8j4D0kK+G2NojSfQKf2Gkr
6ShozxavlbsZYG8nDg+bmqVI9DkPloIJaTw/bauEFBnVwK6R88HX3G0tCFvNLqL6
BryDjYTi1swRG9qOCN0DAn2zJb6fzWrYxowuOvXaKQcx6PRzqFrrYQaBpcAWxrny
bERdGZv7y84RG3ACCK5PVNOTWG7z8QeioWeWTrecBhGomBQfB0ne1QCyfQvk2U1I
LM71Mbvzgbj5rA+DO2HW786zkFzPeYaW0aeY4Mb70hjux5EY8D/nQvhLjFZA/EZV
aHiMZXveMpQXh5AK9iSIIKKFaNZMvndlIFZpxbh6eaUlbx2B8ramy0x8QZZgsc79
VCJMPc994P9vBUh10TFlWDkO7OGraA7gdkjOU4oK6p4ad0EYsaNy6EYdjR5DHSYO
oydqPxd/ZRvMCnJjDXtaxMgPDPaUdU3vq3hzOz6jgQHx9+drrDd127pBN2FJ2JCp
nKr+55yvnS3XyGk8AwfZegIEbFFxgKUMiimlnz2ARxIalFP1ZbpupeEYx0fSAQ9H
P2qA5npsUsmKz4GuPNF92QhVrUu/nu13+AMRl6AU4ogyrgM/kc3LV/9eCmah8F0l
jlS0wJ8k68kKtoM7hA68XQsTMRp7Wy80/dYRAcdI807maNsnGYI8xmoBS8udd772
8tVM75ZZDDMzQu4mb+6v3SNfmVMatcN7j6TGwWLZV6Fb4icKbcXOJndsmR7c1qE/
DZigIZegxK5S8OdFbbGKvtAQD4z+PDoPVCC0R506vpITngW9AEJcGjas6L0ZK3oZ
Nn16VJ/j8cfQG08ZGAl8AfZug54MVpDcLXYiYclWcZcg81lMpW+kgo8u7Xq6uRV7
N+S23JKVdJPwrfJGl/VKNkmfZ1uNYQpTVjf4IhJ9l7CZJVHjLaE9uC5XpVtpel2a
UhXjcbR+nr7S/Jg7x4hgONF7Q8nO2iQPNbBpkLqB1NoZcYcNHjKTw8ZWft2H/vaB
O/uik48+R2xfqf0rdTi6mm8BnaRUtZVFL0MQshl1FlXjZBmegCygyGy40D3NCHdw
Ltnytxz7DnZWk5/Q1+t6/5fhlEeMYKwLC0uqJd9YRRuROdPnBk390RnIFTT6eek3
Mfl/5F88ax4hzYSo4Zt5LXMJW5eOgiB96lKy/u9gPnjSgmzWAm1md0wGRUCoCu2p
ZEGqsl0lIqUF0EtHow08oz37qVeie04E4mVM2/hbyZAkcU/3XSAf53ghmmoar6pR
h85KsEsjqR/kzIqMdFX47+I/2LJ8pnCbMOzgcDTprSmloTTtJvxWTg8wzsqt336r
B2yeEwCQi8lBQrYuXCA0rHy4FGoS9x3hQIGfy9XR6tJ02bDjhMj891iEssi9Zxhq
Oq80exffeV6hSM3T7GmZDvaFJY+VUu5x27cvvQZYurO4lM4waYGT/Fth4k5fLZ3C
9dLv2v30DZA2rHj5+b+t7NBC+N3bIkgOPgSMMA5BTUjp+U4CNgn+64ac9m5biSlP
KsdndE2oGyoFomfH+/UBf7KMBTVluZany1sxfJeZU6dVxdwZleTUTjg7FktPG+B5
tycJ5izIqYzmbOe9qMgP7lfTaGkTuGHcy6KC56+F7QWrGgEH5Phw+/wXPCBNtqa/
rEWnow3/YwIKZhLL21q53B83Z6LquAlZbhM7JvrKOFYTHklGHxoGFLwQFtlLdtTZ
lMmhANWLvv3CneOsbvIY/Zk9OsDDlfPJCsq6A/wuwf505VaBRDxtqtdsnkMMLTD6
lJGQuz7Czi/ZepiRTKzoSN6zsGqj60K3anr622Q8Tt/7cO8LYgEFSZ8voCog9uKV
vYmKQSzxMOEQYoAA3pIwkuX3Wo53HdA2IAuytY87BfJa7Dm6+H5MJeHLNM68N53i
Hhs0HIlFjCcL+rMdWpzIblAWQmU+L3i/Yh+vD8FwktBWqXNUKPaPAEoojP61tgHb
/S8ZzzU2ey5+SwPkvFZVUeRao2QDtlpZwFQvPupa6dZKPjqb7/GPm4Z+OqT4GfLX
B3Cdlb5QSktp7SXhBwR6gL5rhMv47cSFISws2hQi2GnTr402jxpQBgdJtgPZJOoy
TpUZl5OU2mlOUOTHzbdkSAL8sSxg4NIyet+oG58aDmtSSFoRVRPy1qlQpNQu0Owu
vP7znkv44BKY1TJsfoFr0Ov9wV0To5emlx06+9/1/3e/SGesztiPEc7qdJORXOBO
DecCu1Mz1DPCNYmY1WZRtJfZUFPPh6ZBjHfrtUKiDl5+kFnD1owXmpOwnKHgos9F
OXS7fzYEG+FlZQdrRzr8BWyRVL3AwTOn7WShOzjoBO84zlLNXxbVKZ1+twU0WTe9
XIrDTkppCrwq2Ak70hsyFx/hfu3cYWhkv2fXaVZe0M+bhDdhpr38FiwY9V7R7SlI
Gm5MKetEX8cI4AIClUlgo+CqeE7k8oNtmaIwya/ICyrEauWDaZK2M/j3qGtOjqJ7
07l7wDRcYvIx95r9uvR7x8DdsdcA9isKBFXo5c4nfObYplXIuocGu5a/JTUBE4X/
GMaPH4SthLjCwlzruoksLxon19gx4EElxDeCK39v7YeZw/+qNG4GAbO65y6eA8bg
kfYCh7yalOgGN3ZnJhEmvj2JGfhSFZyw21C4gPSh9QfktySvcquiMaTdHYnb2vGG
FZi93mM244i2Yw4wVqjQW0VByt9QvCXF+Tg+rBaoFZpFCIdlv7LVH6eP1pPzRYA4
Z3yA8vQSmO76fM4ug+YxFSrCy287LJF3F4rh+HxFBrDtmtdW/u5hbBvNw/1sq05v
CfbffhDRUuskXAHS7ZaBburzkAqN+uheKKFe3HkNZ8QH5OwHFwqQZ364nfBEDxeT
iQqBP1VB65hzw0/7Q9IETvwnBCkYzYI/WsBlhwTIBAw12uO1spnkUQ61zHT0PRg1
uIyfdcTauDJhy/wffp3zswt9jmDhUYMid8hMeQapqBcWaEgS7KhAKkYBTJjAqVaC
aknJZvvBvjtjNLUgk85SR4EBXOGDdHn5F5B5/2wPcy4Ox7wqp5Aqc3EvQfD5XOIf
+jNANtAHcwoTdE6XdpmnX2BLbPfj+iTWyh69e7sesxsUdC8u29qIaGE5s8brKurq
Lr/pt+uht7innsNuUno/LaKHsa+QMJea0YEeXpji/SkB/D4kvPOOLjY/JNX3RsM9
XgO6gMw5ySRyRGnFIcERqzU9AzIpdonUu7kumbQQbPTRme3aotOsowbcP8alYZ2n
z0UWJgDUmaAje1W7jQIx74yZkSaLPE+uCbgekJfJj4P7CcrH/bM7JX+9P/0QrGEJ
u1Jm7igX0YAt24DQrpvzlLfsoGzJeq4xxn2GpXBLE7L+yE3oJBU+EfniUzTXOjJm
b1DVP4eec0GDBjUnAxNhfdZr20as9VqcppD70qUc0LhOHYOVrTIx+Wby0clOo/Ce
2XChn8jp7JfLyAGzIdS+uZ0zOd8Vbxq+7aFRmABKEtEth+rfYjfUhL4Jd58V03Ww
jfJaOTAtt23FWd+M4VqNfmp+aTC/D8Ncscg6y/wyW2RHLvBLBlKmUTDjINhZy0se
xzl2tAACdREPWYdrYgcAZQVuKMITyEM13fvGhqgjOno+sAWP/l/6uIqZI2kOslSQ
RfZzV5cFAAJtTnsN7GFxaYW4NuBnJbJjzcwNSkUrRJ1HHXE7fjxCMxgZmRUtFhtR
lSG2ZmLGv1h9zstgSyMjKmYSbz+FuOhb8xAjHp/37lbVThv+76bqOaf0bZAvbVxh
wTx9sb3hCN0N91ahczj36WzHPDlzRxs8mAFIupsLN3mk1R/EhuJQPaNxy3tl0X0z
c+Sw1hSjfMUYkxqu6pq9Xs43SzTk6wf8V9fxJTEL4JKeBq4qxIhCXhFstkk/yRSO
iuZ4Jt2nQXUP3TPml2CGFCojF663m/JZgUYW3dbbfVkx02d5BtIK1ZP5PxPW0i8t
CyhdIkXTSEeP7EM1pzbv5SV4VyXv9t+g12LjGiyvfQFg4CSRsg5IDoX6hr+OIhd1
1yzXPufMwNmJkItzj+inB/khKkCyfzhMXqN5V70k+A8GC9+Vjq5J77hnVzjCqxuU
oH4B7ZIpYcQLaUx0pzQIh0BXHWWey7S4uOixQQb1eEi5MO0QlYSwtBAPH2Ys5X2F
Qpg/uHUbbBQYgZq671/KWj39AQQGA06zo3lzk6lrIZfruDvhFx2Bk0fuIz3pC8sH
OAH1IIn7IVtHurngqBhIlHEWzoKfZZfJDCUJk4H6P6MZ8IGh3BgURnIVaRbfRZ5A
KWkswNG3c3xF/IbDWSW5hagAIRhGcowKsfWlSvlgjeQmIzFIVTVl1hh1Nydy5CHr
LJstgBX/k0QKeA1D31fQNv6dhzkes91WXmS7Hm4aO19fX9zKF5K4zoSz8fkoMVpB
JbrS0Qmx9HmXk2ZjNHqOziDjLxOw7h1BcsB2B3OrGGPukG8Zh53qyDgU7D3rnSHT
HHzHDaUifPXcoWDRXAcGkUmDISjYSYvyyQAky+OFCQQunG1pyyaeXDpEuDmY5v6g
AckpnDpC/CQggOjTeb0ouyj3O0vg13tbefJaeRW5Vak5rLKethkiEEKUP2mSDOSr
1RecvOlRpzzyOylqyywHiIu4Ky/Tzq96aMM8Kc3TyC6vB9ymcYqkiyRs83jstqbS
d0KJ/IevdAwqDSKsCjEv3e0WqORQ95iZ0Fe7ktNj7rkOb7Bvipo7BBnY+Hh3LAuU
XunXbORfMDYd2MHRdSzoQ8Om+TPGrjF3goShba2qvMevtrRPnIUlgFmWh1pneH+S
ajaRYIgewLJWGS7/hKYPahq6K2Zm6mhFroQ3NX1tP17WRxadKebNKNWyRzAJUM3c
dIIR8FWk3ynmYfZzcTF2GiiBc1CTJU3+KyjmY5JrTYlyptlDRP3Cv539IVqBYrXg
fBMkQKqkMlNQpfiXGVA43kYpVF2Sv8jzUEimftXPJZFOoX3fuq7eF7nYUijDC4sL
eDu+796Ep1LpgYpSRF+xrupXOWIrZbReVtWTURdzzT08HdXfle8wCj5yrmQXU+sB
/dD3fHHYjl1dFnwBl7c8szYsB53/SVm96a+x/NA21887+zdRsen+Iz0v++hY386X
AHPmtY+wd1Zj/L37aHhxwyQzly2LvvQ3t50ovGYqwihCfSj+6r0T5NNxcdj1ATZr
6Sbjl2Kv99Y0Wyqo2g9427eACO1ksKFp47f+LaEvZT+Q9XtTTi5RYYrzcJaTvXtA
ErZ+Z6twPG1X9jOmYlvzzPD98rdW517POAkhlOHWVbE6aVxoKupyLrm6kAHhcGhR
0vMqQ/WB95kUEgGkYxZ2GR1ymK89i4RoaXwmWZoYjlaZqAbpNL3QVVFup3vNVwBq
BCvzuRHn5zeqflhfT261FBQvGTFTmHndZGbJnzyEjpDoSQfF6b6meEMah2AsqOEa
PNrSmF+9fxZ9iqyHogenUkTW5UQX0OFPhLzsrf2pusFzUCG8IFwiReNL9/Kue18F
KPuouM1tDnD7kIB8lGK+3g1vJyxi0tfQ5TRQLDReb5FUkPJLYEbEPLEB5tAXujwz
hF0bGzjR9x0T4bfy3NtoEfSGc6G3GIzFvPqmHm+II7l9gy3ih5F6L3a5kWRtZ0zk
g9fYzCNXikbfVJpWf6i0Amh8g2JFPwo6KnLJYHyPwnJYinOKFM8Q3ZUnm/B02Ove
jVeE2w3ogVwu4bpjXEvPdSdLESXZi/SIFXkohWJbmPk2z1eZAdnG3TQGww28EWh4
I6nZwhrDKT0kkRi3fVaxKWnO/F26yzZc9Qg93rOItHQ7cFAq1zsfkWLs6Lm5ItjG
y6xOr86O3cuVTnRG9aTw3xXGVZ3N04YrKhVAst664hjB1rF7tYmNKhxr2PV45I+W
2ku5PHG8kKBS3QDRFnpAHy4exkggnDzOmJ6xaM4zQsFhj4Ye0z5+tDnS9zPS5UFT
PRWF+zYezoHHLqnVND7Zsbl9tKxMcEKa4o680LfcIXFn//1u2y6bBsiee1SIqUKX
Hs/mLp9dukYSyqaPTZY2vuMOpvY2lxDE+HuBrobp51T2qkgUwBGlB+hiN+TApe2Z
kNa6SuaRXxFx0+AVPvK6XWsE2ccd0OcdGlVK8OF/E7R1+dtBkE6ZzHMAxeZ9HY6o
9EIzBp7b+UnsALwmOwiFMs21IxWPAjjSFl93sPHnXrw6csPJYR3e+UTtoUuz0FIj
deF03FiLeAIt505qlxfZOnRcmH2pDrGtujAZFRGf0ZUr8JYpPf2T3fKCtDwMiHkr
m5uYDMZoTyxxNtoFKwgdR8Mwj2UD0ynECJZM/JxweXNInJvr/lHeqpkrQNUIdqZr
roX1+GNXVuW3Zsu/UFTEOOvCNWpPOxVKQWbC5XuvJxdQWGggX9K6lS5u3Ie4jsRJ
Dyw57XdPmhWodQav1wc5f8gtNUyA8HlreFIp92AbbGlEekgh6lJx4uiJee+hp9QQ
xar6QuJ+3u5E50MsW+5im5ea3ofz/unUhlZUu4EiJMOBSifb862vDps1BCl2b0D0
wuCtJYuCE6gzwfrCw3RZhmGeIND4nIO4W38zNe3ULUkI1BJPzGdIsmYuLwDpjQCN
93cq69TGBzCtaVRF1ZqCgwFa55NaPXA31Cd83GDgC3DCnrC3ji157kJiLGudx/Wn
F6XMFnKofam756srayag0QaZbhVE77JCMjsGYOe5vMQbUcBfrE/b8mOeruIoAGrK
P7qnXC8wgkmAnbBMGINuY6JVRB9SZMJ16D2iaF48GURD1cRDICwodiNdU3zf1PBl
wOsXbBSq47PLWByEt+VwmXxHHD8rp3or9DnqIrGxPk89vrkOB0VbHwEJTbk1vvGF
Dj01Q0hi5de0vX3thlYLf3HdbEljWZuX8pxLYl0tGyrmzi9KBLttOoEpHMh1aBzQ
WS4f202Bbp8ZVX+dS1W/0uQNY7UY0LMgMAV0WB6SmdLc40ORHIVLKzod0JOZZGhe
s5sjUq6zl6rNgxbpOuxMUOcXK9rJ/qUGPqv9YwzVfuERykNxU5B/jMAeNLnfNZdK
UpAJoUx1I/sfbEfB6K841WRNe537PuxKkOLI2Oq5zLZnI5DF8nPQDKLiEUbPAJzg
81yU0RlfVr2DOuOfHI9TPgOGDi+Z65EFYRXQ8knGRSsPeqzHtx43nugt9FzVTFnG
o4yGxe0DKTNn15Dec9mLP7gabgJEjyta4F4xZMS1A/5zxYisAKC0oP64LccVDnQR
FBWeBKKqHY6mAP4ApYyIB1dV8gij2LARw1eFefGZBR4DSm9DOeJ5tWSMpm49CabW
x7CuMsZpZ8gLpw7PCoeoxVXdnBASpoNzRdJepv6YUYlV+/fv6eB9xFCniQpoAtmR
uk1YlPJIDBww2S4eus+8wmh5ockEVhHnZvI5OIUiWFNRaR8ND9kK5ZPp75lDRtZb
e1RJHfLqcaZHPeYQ2z3bTKz5yY/WnMsAr9S/UP4efW3CzVnnTsqzT7agSX8IGXP2
JLYK0MxwoeXXTn4lTo0FqTKjobY/J1VJLibDNuGih4AWjgx8PtMeBQ3zkSwbStcO
8mRG8Ic3lPgWBNBZtN2sSAMKQLGzbotoaMpA7I1mIe61L2kscRZ2+UahmSDLN3In
rifHvWdgh+sTGoQTMkYD0b5La3tCjUOXnVHzZK0L7nUgNtIqJ0AzJ9zBfUSHAFsi
q+wZDSx9a+/X37Cezn/MwCB/v7L0/8nHVuwIBtl63ckKzlLP5cDTAV3lzQwVlmsG
Vdmst+vSd852EArsAx6JwJpS3aBu9qezvzEADGQ9WDmWqGlezuQkSvniaP6UTc3b
oYqg2gjBGo+3RQqdu1iAOLHwPo/SE9QazMca+hPY04YaQrE2aTIDcP2EH55vbvaJ
HTYxdRImG+zbwyoM8soxUrx652L2gM1M/F7joqprFH3ljaQ89zcTXJ3q7fbAEt35
a9CAQNpzqAEw/sn5mulIVtwroOHeW11fmMg03CSjaSmT00aaX2etjtAUzLWEPQc3
1XsbzkpAcD6VfnxP2IJKszDGejtslvgImPCg2XSGUn9GwiBoWq7EpWSdyhtS33Hr
4mnb+2apIFyhRvN094AbfsPyyOqvhOTSHtbEYxFV6rq/6HDldEIT2eA1ksRG1QOx
5ctapRKJkxKitnnx1KoJuQuWUockzM0lciFJjs8/bD6AEvPsoccIoJKkns2WYpH7
cexJENOmGmENokY0VdFkXX5wjBKLdM74y2eVVFZM/7nlmu0qm+Nc6zKf969+8zsc
IJAaBw7zk5dCtjo8TDSHHIWYqsaiYZ1tISoALT2lxDcYMCG0Obrwy7oveSCIpDnb
uEaLDiD2NQXtFkMDurpqQd57+d2/sD4kOPHpjCEDUD659UZ9ojhWCrzFZH8TTgu7
o05E29Ij1lDK59hgmkwajtuo/DbJO4qJz2v30Mo0UWjNhQD9bI0/Rhl4X3JVw/XK
NE6ilM031okxNK/QYLFJpdi8oBrC44O/ADOYgyI+Pi5A0tnCyhCPfuWwqyfBUYcc
GzMQNUme8wuBynkU+e+57K53d8fjxCOzoCbbzQHrnk1Nly9qUOb0wL5s5c8Mr/HO
yA2P5AHlvprSLNMUYKNk0dj3T40cDBlbLClknsR1e0TMegkq80WaGMcqKhqI0XWk
jxOM/qsGbjHGLiDRzVHVb9zQ31YvnoCbnsuducw40hK2KO2l8y/5ki0Ug1TSiIHH
jKu3IF131TjMYiR7V+A8lYXEnFUNa1Bc5EngV4auE6XiidCZj1Xsrv12rwu1ZTlj
HWY98JzgmADX/0JxPWF3kviBK2sVMNAVmbwCpnHPrRkNsLuydo2Iq78rbsQQfrUc
eVtZiHINQsV1ZbNMYXv2krjKBDkA+NeZ59aNb2y48eJpwVNyknm4226HvsIqvj0N
UeEWcvv5EkwT+YgW/wYM9AahTT7JUCZriFgAG6S9l5RzNSaoffvmGY+N4YrWZWeT
yFHJtVKKLaSSpjZy9dQY/VnPJ58oLbM3DSCiAQUm12or6icwJEDD/zjFq8tN3HKk
3QVF39D7ePb49ep805VwaUX4+t8SiocGkXrt65qF7Is6Rypxk8fwhvfRuI6Ay1VI
HsjGYhDwBpceW3avHBCzAUXHOinaftRp542Ny0+ex7qBN+OXhD0nSLnBSbCabZjv
5EGiOVhJFHLGXIr9Uf58PwLx+i572exDo7XjDhi+h/9afJonTCosDmDrPXBo+vuc
Mb6z8ROU7zy7APl+nVpuC6tA+0s7/C+FYA1WDnz59EVmF4ok9AlFIDTlQx2c+c35
MEdxElCSq8LXTmp67EH/1glSM7VRZSi8ourOHfknyWzw/NfLM+AjJH/b0bLaZ5DL
2wPE5Q/GVgmO5gTP+qdAQYkgMFzh7T+3hBeE3fC4pl4eXc9XDhXfrFGrwoPhrWLv
t1AK3GPLR1q730Jl92uu946M7hWq8Iof7W/VvMb58Lpr2Dmv6tf+TNfyZn2wgpIY
rKItZfXE9zD+JzxrkThTFbYmvOsbpOm/6e+xzDLjxbdWBZTvTPYalfqh95bAd0cF
a8IHXL6AMij25cAg9SNC4sgWLensPtnpVibHGHPF61pLOd/lTAUG3t6a7cd9ixqb
xL6czlimq0Nx5giMfCUErvOdW2NsY4PTyteftSCllD1igzgaYJlJpA4TbxuqY+cB
KXIhmxKRBM7sN+JQtoEBX9Sdhk89yTzbnqCXWlSH0bz4SHtLlzoLiF8QSbD4sUB4
1WhS4mjnktv6poP6Fgh+rmdVcQiA82M7MnasVKiXLsIMkyzO9KUPXrR/H2O+HVBW
SJd1YEYPr2Pwn0OUcMALsIU7ta5yRbyOmvGPEaEPwvzJeV4GqJwcIPi3quGOXtBS
Svtl9kSjGlgVQkiNr3GoYxr/XIL11GFgwZ7d4q0i1xTUMEPxQJXEM9/m5jK2bEEN
Umm1Qjf3UqF2h59R/TWU16z6NoIuCuWhjNIQgBg8gwEQ3Q4Kmjd3rQY1+aywgPTd
RyNQfis6eHoaVQf/iE+Jmuj9+S4XOt4+xWPwssMQDDkz1jHYWLvIgkBqG7y0qOoq
QRBh8fYh4Am2TxueHoS9wvN4tyRt5vVYNEHeIU5z3/bgyc7KhpNM68k3f6Cztviy
Pi+M0e2HH0TxITTVdL/+VrrgPX3CysYt/glLCGS46wAL7s8dWfvRh1nCaUMMhnrJ
Kx54mAwM+6GN31zrLGoWA10mmpfHeATl4ZCtDsTHeMaQ7yJDCuFykpavEdumn5Ix
NH003zNhOV+YU8dzIg+8wyoNm5gxjAGU+7JtnPJAQ3NztV9M6GbUQDkcIU8dHl1L
gU2RQyTUs/9lYdk38gOSMepNkmi5jFIzW7nqLfWlODqQyR7xlwFdo/bjtwdnoxSX
LIWS9P+k+X35zeDY4pgN+hqAWbPSIM3E/wlGq4GT7fbazIHImNVQy3nTexNZfKgE
pgS6DBe85IC+TufeFsPFNtvUTpmEC3Hm81lSQh+XD8HG5XVb+wDYwdmppDq5fLz4
KREfJTEsmzAWx5ZUIwSD35QqQc5vsxh0+gbkcufxjHGrIJm04eYfWgcIPAg53Fl6
8QRJtuh5328Uahlpn4zw0klZUeKG6GalWINNLld+n5fc3QFoBflr1zeiVeD7T/75
5ZIC4YvkrjK2USJTL6Mh2Z3a7L9wS2fMN+9aeBmzgMQUA4YoWpCxvlN1rdpGw88Z
iRcsWqWJ60lVUMKKxCrU2+/ZGAFAudqyZlqV3K3yzRBM+3+DeL2klMFh1iiqvaum
EuTnqio8BBG8P6oij3tLP31/FkCvqD3IFQe9tuYtw3cD1ymx39q+UnRCmkNJFRbs
yqMLoAs0PRrkygdjoH6KdDv8SXe8FEKuEsrgwRaTWV8QDb498LiPgg4Fm8zmlGDk
1rmKoKB3tka5UjIjMtDn4fshjp0J2j6yoULTagMsRi/mqsY0GDAoD0nfzlLRlQ9G
paxLoqlGrlfIz48a57wL0YMyL6QSnPqZxrbT0/LrREByLMBwqIXudJrhcMF/KT2J
zCb0Ihp8oNaFKNMypIezQay6Sr//9B2gtIvo+aAFcoEalrFZJasBe9zyr60TMwMe
P7XSEfMKgWN8cRAZA3Z+7kQX//noUuTa7/FzqRL9Zd/9KJLDwZWStVvFeYR1/ANH
OqU9+FVpnTRpBymNo+bwEd4wJ+zWvSd+jbQCWJhudOxaHhUKKb2CMM+Co8H9otbR
LhvaxU9y7OINJdRHyf/nvj8I8KT3ewnKAErjrUBrYcT7BknQO8PGOpZ99yTjqY2d
X6w2ddk9230Jr5gnClTi4/Paa77XkkPiDI993+Q7Njq1BSPYOtIqHmWmXkM+AF0d
0LxfxuKUL3mEAmXv8blfmdq4dWleqDc9fDS16IrZVc4q10SJEBCVPrjJYqEFx6PC
bYDS0/UrVg6scES9fV116uoCxefLw+56X+3+VAbp+L4cfdyKQrSgmXhEdpXpVoZK
tUF9O2ffW1KI0dYYtFlNQ8imjDkmPelGLxQOaDHa6XDKuVwuvDJAkV5SSmkabSJ3
M2JLLJjM8VgXZyavTU5uA5Vn9JmOYIvygl1lUgk3yJzoapOkJVF7T3t6FQFGBkbD
q/8wVyxKcNMdRfWJPltY2bWqErfltBlylS2PKaXDNhjZNCLsoMW/TvivQjDXaBsb
lRwM5POe2f5xkpVJaIB89cOWaqtwybiTWln3qCKez/kXx97ND23p4Nyz7d9aLlCK
XqlQhE9xUFoWXcfNiHZWEGiEeCyb3arWE6SG/3JG/Mhgjh2RpAW7tlOUB11lrk2A
IeLJk3oxGOjdXm41t5TJ/XX06NEKxUZzFUTSkwnQ3lDXs4UaUb1XLX8Jdhy6mew4
S/j0km/MdDZ+ewIKRr5emJhuJe46B21qFfUYqX+oPTMowQme4w36+ZAMNOvcA2j5
/g4tmwL8X9DIkZIiYk0mfz6WGOgTtto1S6Ryh8KTg0ZxLTEi2swkEvn+XBZQfiaH
BOf33DL6c3jWBJ3IssY6NcYReNMTMDnOJJbgiUQZh9v0i0ZvhNt9zx6ydLzjjsmh
CdMVWuZ79oF4lyPRGYXGG7pNwcHc16OO5UpslR6fzLAGO0IEXk35J79yKDls9oIR
F2za+ejJu3Uk7S3lfC40EncigYi3x40XE968H1soolbk/sep3B2arCOOBzIHFnyU
Rb/mu0fY8ZT1bcJCMdZLQbyl7+6HPeTcYskolBsJSBIvmjJZ9A17MaVTUDXioYM8
++7B0TZgCeCC6Z9Fi0L3iTHxPf7XkVGJhCfPpJ0emH/olpgGxxHyxwtOXxdAatpe
5XSLmn7Qz0W6PeRLUO7WJJAmNakowRiQOmTIMCb1JyuYAA2b84y1PK8HkspalWYV
5O5Iphnix2HsMCbYsn6pSabhxCVpa3X0ErvM7tX/1Uw3fFcaZJabENPZdoiUYNSt
x5atMhgp8k/ED2tKjKnIbLEpuLjBKpAu6BYlf9IZWW8kHjqLYUu0lsVmQtEZMJJs
vCEkV/pK8Np//jJObDSdUZzEjeapqJca0/VfxtAOtdLD9JXww+AtnZBL9RyqP4vX
8zn9I8m9iJgt78Wyge7o8WqT0RWyf1zL9UQoYe23BCHfoY6OxXQ0eGqz2ph+i+qn
gQr0yd6KqAtLBSI7iqBBWfCuR7bkgDIUPybWdclrS+9rlPKDpvieauPT0cSQ0QQD
+5JDAK8zO1X/Jc8Fh4gEYECY7f4LVR2km3xX8a1I1b120JoW0m/0cJrN6xLPEJny
j8FhFnKy5hMK824f2Pg0auUxRJzEydJgLQfB8wcoe66Lo6TmKdDisTLh1eHvyQli
/v5jsnswv8Uh3miL1w6M0qmsH0fzIUQQzaZeSQR/03GhRXbp3w3bGRnNMrwZbbyX
1blxzhvRJXrygBKLri6YBrnk4gjuAz1Lz85hpk38C4rklnGLwmIRx3aLqJcnxCrK
YLmY0S3kEKcR7AXTDTYPn1fkdRDFATGUZgoAzQsA87s/BGl0CVJS12m3+/KpF7DW
WPebSyNeYKXnEVLVlLzqAWFVVNIT3D+Qxgd7iEZPM1JDOU1lLMfPxME3w9wPAYdp
99bkDQEiFmNqS8kCoER9ZCuHk2oM2+4PmOqY+ub6DdjntFFsYqc9xgDnxmDxitVy
JFlDSUFxACpPjQ54BWyhGbllqN+cCtMGFN3htqccHxNFiYuul3Y3c9MDdj/CdkMi
vOtHDQpYxvJweMcvAgo+h34AtD5oPNhTchJIMfUlZS6xdsY06vruoxh6zh0GrC0n
0YBSLh+7Q1QFHYvmAH7lzPAIA/d4QXvIh46FYvXSZhUtPuMnF01xrYDQoqBOeEX7
1CcClkpIEN6fZ4vRSIixBF2zX8FLRzJiuHPL2hiC10dmI9deNfJOpw6C7PV6Bq/B
TghJkpjHFbC05ByAKKZm4j25Uv+6ibc16cNCBDtIh2blOZM3RAKXU1Ckg+bise7L
kgdiuhwdDMU1Nqn/Wrp0ShJBlibPd075PkKdaUDsYbW4zW65XnyfBVpeelaO5+nz
Mz8PHZrpZb10LEvptTt6isWTRvCQ6dNaYmSvQFY6uHVSDkE7sRZjA27eQmuhtiA2
PgKEj8Zqk39gE7Z3MfIQFmY/q3enZ+5fjUeEkfJFWVPg643GSEuEf5IgtF7XSWuJ
Ow/Se+QudvEWtNfedgqlo0N/wxllMIoaBLpHQD5Do0GWUNuykGGh5EsZI4gGCE+x
xF0St/0vsxUxpuHKZdXc6LzJ53IaNVgqaUmsJ+DHN3Nd5Ho/pCzjFBGD5HUbbijM
8GaN/6Pmw5x9BMLoSY1+OGXonw67xoc1QIUrjL/9mhQwqLTYYZQB2yD62phKO9r1
ZRrVM38BBGSSRIObkYHrVGLm+Fm1BUPlz3IKWj+U7szAjTBUdTvbKTHTeNwLTxnC
qOgV/XewU3P1xoJXdEOdHYcBaE+f9OzeFWez2sfAZJb7ib0JTPvUBAqAO8GEnZJL
lVtdm+HCUTzGrhoBwlestbvld+HnhYnJEI3tAZg13J10abpECuX5SH0GY8qmRy1j
1BZtwjYvpQm/TDsjjgVQplHovChKHjuYVwq3ua4E7RZd/QtFGXOD++9p3bHY1pvj
8VstbiniOWRAYJUmuj6G+oAavjcpzdz+gBE6wGzSlC0tpLsC3zv4IlGx+NXyPGm2
klbX9UThio3czOTsyJG7KzUkWsiWbwYW5hJamBoCjglbuSJ0gBulEvh6P88yEnYq
dA0mo/myZ8Z+FESC0RiHOdb1840JhFRxceAbkz4LwS64D66NJ0LyRUO+sHKzqfOs
/H966l0mSre38JeVFwBBlj982tZsBCgQMo5CJ34xkDb66rjX22Q6q7Ckf1UcSB96
qL5IjTjGLN8zlIlT3o0xyNPL9WVF/YASSoWCC4HJJH2ncoEOZVT7xulzsr6gDxUG
73seJ++YsjOyInGYzuDMa40EgSAyMTmRuHDzJG390JUQms0c4X9kaMpi8FolAhX6
4xbrV9+68NHshakqUBhZVfTOME2V7G3byJaIuEmEUPAzNR9pAGpqv5yhcbyJCnCG
+eLRpj+boFhszVFKtCdctdQfr3I7Ay9+Kj927pGQ3e9D8MmtKXs8E8Z/WbYpYqTe
H637H3mAcw8mhJkSJPPf15Q784iCuJuuQ58HgYBtNEfFxv3ze+YcWrpQSVada5yv
tjEe62/a7OnTrGVd3ZC7y5PVsgy5VhdSbygbLo3HtfZnf7cjxIlKAGLxy5equdSu
E7DF4PSTuopQ3UK/KoFKvUzlOFWaiVPGNXppDotYbBdO/G1lP2N2WG8jEcA8bafk
/pI5KvThrDjXIMW54tEYi5WCHBa5ejrb6F8YX6To4ka2ECqExmdoMmw2iBbMVi8n
i3k6fb8kIiM52e9VwcF3eE2JvmdKXcODaHP4IGiGurFWLMnSq9MrLowsAEaBfFAg
engfWp/BlG0bJPc9cNfkd5HPRgItuDvX2b6Z4tpqXvoCTAJH6kPb82q+3eEgiKAk
t6WJsNRNaXtWb9x3eiIbRmdx5Ud5E6Q4x7+xW3ssfQJpjhd3CDDJ8SyFj+TwSHeq
ltO6BDl+tTPiwMi5T79G/k8f47bAuHRs4fvD4HRahzKTQsIlHtXIjII+o0yIY9Jw
C2QRZcy/ZDhRMFomGPoVW76b9au2xVC6R4BEHtt4W4PKjUx2Hcn+6+rmc8uPz2QP
cYSZOkXJMMEEpwF+Y11f+n83JwxgO8qejrU4Qq42ZFLk0ZfE/mTGZyI3n9qt/YoI
1cLveMt2mWoJpsvMqqoPHpTVxTItAapg9loIDoe2cYjqYg8TZ9jiTOPWAe1w4BO2
66EFfvk1LSbprQuR0FizX/ZiOC183K0OxHeBHn2KDL90h44/ZDu2B96EThh/75Bd
1WfPjAmyV1iJSgkFMvsowgLi4RN72kBCVT7B6oLwJR3T2OB5LABmtgtZmeyEgTGg
HQQH5YhO07JigrzrdkmvpngzKlwnG3nKHK5+wfmZ6xXEgeBkjyQuIQ2Tbo8yMbnt
q0JKu7Oe5YS063GUnIRN6gje97QpRV8B4ab5Btpgwn2NaXQ9g13jGHHKxIHF66ee
daFBWILec7ef0tjhd8wFLBzSSWR7ez+MaK/kFafAYevCh5IGYCiJ/m2OoMg/A0Cz
ELZFUTipyXlorRt7RrvbKW5wCq5xRxfGfFsMxB/BUP03VE1XvDHP+UjMbqGeC6bj
5pn1hepbeO46roSYpUS+pCGGgr6DlKaFX7zLiv1YQY6RRTVPSQbZlXdsg3l/ximQ
kPE3d4I2O6osjDV/ZL5vxa0/wJMaXNfA84CZAbzt8x5C37CsjvUaaixfAjeKcogX
0B9pINQKDupWdYXX6Pm+oM3xWA18zOrM/hBYF7P6mQMNZB3BMsekQamdASYZHjB8
HTKLolMJchjTWBzRcNgKON0/InxhPaefSuXCiQDfhE3aP5F2+q9qxBDVpzwzd1yS
cm5kQV1Tq46SATN0s0AHkL4jhkIKcu8Os3Y9aPkynjjCeVKBoAPkV5ZybFv2uWwh
n+n3aRGKvbZU2zRd0dYkIiWPZFjThIg/QZvBKrfaHsFKRcmiWc0oEace0e7z69DU
Wt8/JRNHTF28+yxRs+DiIiVnPjpjxjCgF/G84Vh6D9yFlvizT3yRU+xjQm8MFykS
9HPAIJQVBFDx0ZSh/FIzExpkB9UEJQeDbKfq/N08z6abTWfGj4q53eTjujLr9oK0
AMPZDC131kYOcKscmGTGCghL5C8tn7gt2hsfJvxBeRAbUbVmkc6qJ6HmTKsjPNWU
4xlwYGZUULhoJ0rqRNUQ9xJHaJ+zDNGZboFIhSYXgl8gVZ4sOfsuSzajpaqXQWlt
uID6mXhdiLt+LhRIbU7XM5/OAohqbDDO7gWDGIsKLPZLzXZSXFq3WJQwyKk1c0uC
fKOM3LRJuCc9bObrxnX6PhmXWr67srGOrsQwIBISkiRozWPSrmEeeEGM4dL+ITf0
VVTtVcxArLl10J98WYfzuHhj8iyvyRIihj+W2HskvXslDyfybwQ6/Wfcd5udd4cI
W/KdHR0TRlGtW+gU0l07Un1gMA5dD9uFkWjMWDRJ42oqmkLsVVP5JiWnCMyVO9rd
r2OuIT0RbvdVOjgqYKFSvMg5EDeEFhekgAxlUxF7YnVnYkiwrvVPdEJr3iDLnVNc
gIUseLCHB0XThDpb7FS5INDE4Hr90RRgViYhLdelUdjkbnZA6ladeiv5Go4bWENG
3wWXixzsSWOPgo/51x9+O9VzNTLRqTYK/UIBeruAcPreh3FuxGMmeBhJADSuN4kz
wIhMUbeNN2uaEw8suMFkCNvqrS0upT5/0yeBOUmf54ATcRHI+Sl4NU3Sg+5P2QYA
DYZbSBqF5Bu05d8kZzC44xg7gfskhZDhdSXM/C+2Ipq7umqbD2rSCjCVy0DrULkl
hWaQupuIEoHbJJ804vpjnsm24V5FmXyMeNwdPuSWggiyE46S15dPSlp/y0xgF2ql
G/Y7U3oXRsd1mJqto4vwF1r7oaEj+41j++cvQged65Mm/FcLVnGyB9ViaEgyRs+E
SH7ZT0ArQPKP0Ja3mtiYIrIubyylh96TqDZH0R9ot59o6psjuv5xfQ6PwnekuWqh
BZ99CkP4KnvxwLBl2WnozQHFvPWBYxgOcE47mpcGs4mxkmogeXXd0s2ZD8iCiZIJ
Q4zn8bRk6sRm3n3henzKBm2ll3a2qEkeMDkczXGNAKaZ2fxTAmjyN0WgbHLzMqcR
9vb9ggPLuoOUa+JWtwZo0x3oT3ySCYfT5sjS0/DV4EwA1dT4fS375WcR9ctpxJi6
BufL4a5W9UzWClJvfWMh2rnqQbOcHXyXpz0LK+e5AYqImgC/tsFSp7J2ZBZ84YPY
7+p75w4lw1+KDgMW1IQKVjhnV0bXCFYxxWdNkielXjFrYFgJGdrqNxZRRs97hMPq
K/6bXjgSz0TDTtV6MhsK9EOyeRI4Ss7L8nAlLveUsrT1U3G8UrwlyXU6ba6Fwm9a
KRu44V+Bjsc/Hmm+68hKo4pR9Ck2kRAMq5emeeBVMaDGFOpdULgDMF8RUryZ5xHN
j9KnETPTdZKVIvjhDFpqw4kUAfGIqIEdHYxMmPtrP3OjanzR1sLTsFHkLGqQBsc2
115ANBeGGeZT1g8LnBn6ONXsIKyDv9IDZyXGAnCvjMfIGpH/p+CMGWxFVO/cc+8c
5Up40eGGxgMqDayX/V+ct6vMUIs2kM+jmKzvj/bFmGMNm0KLW7JzcC6Qd9Jahiof
FmPZuAtyUsNSShTTRJCYjGRDJ3L91MDjgTDnSybiYY/5vwbtUQ0jpKpWUtOej/I7
BfoHN9Rbk0xw6TDLrR+HhPAEO0weADc3yFXe24QVXdjMTK6+vqka03UQRN5+5Bsp
PY3KbPvakzlht04nFjUh4MFOilOJvxydrtYtFkS7AnNntkcTPYEz67XmIrXUSSXL
3E0JO9pbygiFhM/8bvQtqSzRs6xt3VoerlYFA991FZrUVl/8ylr0ykND949NeUhR
QB0SQaV7lrMSyOs+qaPk1WQyzPT2F6mPsOGcdrFcfRkk2T0SVSIbcJe3gaR206DP
vNc6lz6vQ8CAhhtrGraQZ/Q8OahptwK4UUSluLO9EhhMT7po/0Qx1hyP+T3p/0eH
Y+qVjkBjrbwFJ+pxDjVuqazBzE1rkf4eXnkhQJtKFxM+RmLVJw/3qzzaAWR+FlyA
XTogC0lTLUlQi+HDYZUmsKasqj1uRE3pchH94mHvIbiApF6BkA1SyZISQJL7qVE5
deZ2XAi4vZBykHQWkQbNffewYpbcknd6T14TTuVTp+RlHQxOZanx6QpI+pAiW/Wy
npbPMwvOmZiDi15wY3FHhzbIVH4s8IQQLF8KfCjWYgX/kMLLW1L47dbvZSpO+9mg
VvVeHgYb4Pt9jNFL0dRTQVN65mehKZH4k8cmxoSYD3NY8N0KU4bIBhHHoTt6vxJf
aLMNkkwOKc4wSn4RqVxQvwxl/3Xc3w9FYWJrsYeeH3lGvuz/+mtJOC1e7Yxwx/Uu
SZ9QufJa7cCD6lt4RcTukGmzHLH1KQoVhQyheES7gKu+Tcq51qSKKPj/UdHr17gm
yk6Fuw8o3OQF+nKQTPSf2CzOHUELOsZniuc4pk133UNdrBE1rUeqaqQaNQegxvtZ
DbU5k5nuAN+bA7bANmSWO06vmXSIbxFmN9CsXcsOGOLPwQUoRp+8exTWggt+Hh71
bIBRsOH4Hm5PEuKTCxDMhF0s7swmm7fW1kcd1e1iQCbsIcHcLhVf06cF8uWEbJnb
fKUNgJCujCMCgZ3QToMppK3uMCJxgZsCaVIMz/QK0Dtpg5CmfLb/6bB3WTZcoMT9
LE/aMlP8jP4zgZUq3U7ntvbejgdyD2x3bLTL++2fAZsl7SfPCr+60MpMk/CJ5cZP
JWPeqq5OAB7YulTk4O47Oe65TJi6ZlxfRDzlo9SS0qQzyB6Hel4QDcmz9SlknFkX
Oll1RB7nrjyGuL3nhgwE7T+ex7AOYPAwNbaVR4SM+cjGf2YEzLG9QShujmyHUUNQ
0Cs9zHgkALWggDsYMp4a4zrOOPYDat7Kid4RjZCkve88lCVtFjgdRIU1exSTc39N
oa/4/iDYNBeoiQbDRjnk1jy3WEZ8W+GaM5hdecxbG43QXgg5CKklKe4MBpwlGalX
TzrDsT5lciVeGHTtlKqdnMNSEsrvchnfMI1FwEe7pLluRZJeYMGxx/loUIYmxdzE
uLsVvVsmcCWs4w9FeMcDv7Hm8I2KgmILVNr4hKckWU5I0KkyLiio6Z07UsBTY301
V3tp4jz2ZtI9Q+wDDYALo1IgWsBnQODnQvAm5yDWEv5kaj6r/mvjbr81BW6+LWuS
LdjLRNGeuDfIDdwJuso0u28Q7uUrGfyGFP9yEhOn1g60TwTNLMk0EkzY8ffO4jLh
8KeGOGpIEkPsruQ5b+B6DrZZRLeDybN3rLEWYZNyeYCjHDursxyXPNN3oY/Pzn2M
5a919zxK/6TuWlEn+U7xgQ4fuSfwhmjQWafY+dz15+v9kMgA8rGOmF26BobnKnQt
JqZaH98VsUYPeJxahPFgo9Q5gA0fgqBupGjviH+zWsn1PWuN9sHbzo3JRr/oD/k/
6EE+iIbOTfqx7eNiv9IbxMB/A9ZN4wbDHU/LM8NnIn3teOMGXOYu8SPBy3XCt8yH
rgQEqDxAbp67o3JXt1t/7MXHQnv8VyT0aAA5nnyhaMe91nRdzQrV7gBIDTffkfbk
eNNocuIBT/0ZbHV+cHntY8ilrdAD3/DiHMsHPb3jEQxQQZXk3oBrPUExPT94d2ZV
eRuc3isT4vCC7nR6W+j7tZkRab3YA8GyoFAsdsREq/t2q0E592URu9OZJG6WnaLi
Wh+7AzDo5cmoRiNHVZwphxDrTgGOwnNsugQDFiPfF6qiA71qUvuY9tU6viKyoRJY
wR9T0ZBY5Bm8Gl5kHdfU8y0Po5bZj8vhrB6q5YIyR87YZxFJ6hUny/uk7qQxvVU/
bbVk92eWDEKfpE17p0UC46MxByrz9chGpwHbcSwaACejzZ5o2FKO+lf7qffdriJ2
OyrRxBiF1mKzNufJF8tyFJLJW2zNRa43rxI6uUZIW3rwYHJCJicRzUKVwidtPPaN
W3cLyw8OOHpeydTGSBLH9lAPP5Izv5r08F3uvN6ofPp8zEsF0R7Iwq58LtFFkEre
dCryq6JIhV/jPhEvrWAP3uOlHPlrZRE+l2u212JzyRNMR9cNxit//OEzFqY7x5L1
I+4KB+bWERJcTEmyeeQUR6phs+/Cd6JORWf9OP+nqQaO04L5XuSiLmcUsDiNpf2Y
QlICGAzH6ewecbgHwyC+gr2BQiqDgQmYuITrZnwt9QX55kjvE5m2DYBkuiR7c3Vk
+6Ms8ND1/uYiCCnpzgKN/Cyu25luqEFfU99aRPTRZIFviV/KwWyyTAPA3efiQbnp
SQ/i+yEto/EMt3uyRY2TdF8IFERMpuTpNvhbHj20AKF5oqBhJJfvZGuW6tQPhA8v
uYyb/28u9Kar3tJP5+DWwE4/SrTOcP/OK1XzEM5J7EFZrHBPpbPMnpkCh4zrk6fu
7lYALY9D9N11/4Wsh7DIUgJt8dB3Gy4PyDpzOnGrubhFCZk7VSjVG8lAWVW6iKaN
aiN1MOUVsEyKEGau1UCgHd1i45tjWg3Qbuq6P6DfPl+Nr7S/s/8LsXjQt0OpRMg4
zc9SeUKv7WbYsEQ1m4GV/tuOhfG8gLT8El/WymqlTzZVeqzZKF0KjO+CeVO89I+n
k3ghMuy6MNSUCbMJSvWplckC0Bwg7RkKL3tD2E7UHCGjT81ocshiR+KXwT59BIPC
xJ+UqcNfuQonWK6u3mTBJIDdCvA8Zs+Xl8kx9kwMdcojO9UKJ6sHHaPmM+rCerR2
LUqgVZ0LHeR5CiUZ4IkROyGfuOYjzpXFm854b6OE4KEsghfK8yTz5T1kOYBMNbyw
4uR+dIFdGijjUpjz6GZnvgeOqpn6sfC9XK+epcXGv/7yh58u5jjfdfGSxfM0GKa0
fGlkSi+/OpyNPg8hmAWPEMvO/+rMVnNq3bm03J2rFBMnr50MRG68KcLRrYutcJnR
CqRITdFIGBoRSfj08ikQ7ilHTwn4KAF/zPC4bVdczk2xPeMLvMshZw9XjuHdUmfn
7sCVHNHNad7rOPqV+2IsX0lBA9rH536uA4Ke06HWSW3/XhZl/1n5RQ3WLAFZ8AlZ
KsJPjwT1CPFxI0mBMiuyZdw3YBS0eR8y+OqAFv7N6Qx0hBIewhSkFUGTg6flcOEu
uomxkLRl0Qz8hHKo2RFVGWkko4WF/5/mnRkeirsEeoloKPFAx6YMO2cb5LUpe87L
Qnx6ADMNk58ByS1LhFVfgf9uFl3PmMBD/UT3wn2TXZrlQS+vgGHBReWWyAh8MRhE
C0lUVyR3lB0LeNYoSCvtQdM0r9dR9jm0s3aYNVypA2B7SwArHla9mLHQuce/aUdb
TlvVKID7GtDoWbV0RlJIsQ4XfzkoUAosrhPVJ8USCoBI9m9ojq++yZnr4jukbQN7
kcUXNRyLKe+mSKWCJaiKOzut+UC00qYX6uVGCLA1nKL6QZ6jBREjy8G3tRE4S3nj
cN4ZeXiqfj7EPY+nCets7B2DYYFUYkn7wiB3MYkejGqDJPTPnM0jBdHNlBsLA4Ii
ROOiACKdoGjMA7gkhOUtAzu1LbEjFpjLNMj+4zqWl66LX10yhlyoGsaowQ7gm+F+
OlQNzuBH6fA4Lwa6KK4/gv9Qg5ZNCl9++u3vlBOKV2D7xdV7Rsh9j8FproGbIWzO
D3V5JUVR2SXdZKlmYm2IDYqhhu1uN9sS91d75qQgXsGofdmKT8TidOHXnbx0VksR
1pJiyvvNBk59mWAMwqREcfoCafcRixkvVSkYl6fJbddKOHjZcsPAc2XOw+2Bwg6U
O6HYnIROdihVZ7ehxGTeeCio4WG0wL6uB04Itz9rzUd0xr1/b0jwUv5Rr+o13mDO
x1KJ03Q7NuNNIsWG6AgoIxyr2mJcD96uKZfjqCcXS3+U2RW0iHTMZL/cV2eFqDmW
pAk4PHgu2/pPDVAaQnrULb+rR7Q4eXSl0SxjSLrVkFFZo0EOfl2iRbdvB48A9J+o
iGnEtKlHQKJ2YW6+eY6OVAEpZosjY/V6mO/SOULrf4IwgVSZ6+rF9wAbaD8plTm/
iznnHBRDfCnSgfszXRJktdQAMcSL0mlnHOR5qlEDNmRW6I1rhKH+NrxtjBEnFPqV
XoA7GMv8FwtHwEJpZsXZFOmnjLbb9CPM82tBEpwi9+1fuo0wZ/k4KQAzK+nbccIu
+QFS4GhgFMaK0igj8UNE8Du0qz7vPfmxLZfLfUmD5ilm30CarUB/wZ6Ay7pYLfbM
Qd+zoPRfR1Bf4dVikV3dKIDdWzih2VWuCWl/Sm4/fNZe0c3gOgeDrpWR2FTqIeDp
xbbB2/ljAqfXKY5gQRuYYw+lj3+99gyWjEjBDcIzvuV+4uYsdWDtR9LixEyNsz8A
deSCEdi1PJi6XXxBGLfrkpmzmeeeJoljRkGF11ts4JT4Pd8TMIBo1Y3n2Gr93sus
QpsqWISrjX5hWi9f2XpEiTH7Rf0PKblCGsshQMA1oZmR65vIJ2Vs2pMdeP8wjbZu
Z5+WzjLw8AX3EoffbY/An/b7lOShgjcYADqXljZOO+r1yUHQX68JgfGyA/R6Fj2k
K0p4jsB5l7Gdm+h03eVw8dBEvF54ukqfhnuTqGuVlSmWXfR9ht3uu7R1PwX3ajVs
uzpk5UKQEJbyZ10vj2d5yEXLQWtl+0vaCHuGo8nZSyOVZqB8E45Ej3rCpfqJzO7k
CB94PZtAJE2p1evZ1J7+pSFrNbwS7wSg5g+Kcy5BKipYHRNLcZnmD5EeC6pnXm9C
TMS3SAJxdYAlcDLDWY3GaprOEW3AaAb917GTwK3bL7zbJANHgj87xbWWkll9DcL4
wVUYlBKvjedJQoq9oK/SO/CaFwxP0kNUwLM2YzPmApg/9SO/m2nhtss7cGHCvA6r
3NBEHumfpdlIkj9Q2EZh0TO0q1w1HTxDnmbRgcyatQm6fH/Y6x9PQ7S7tKDZBPEL
loMItX2cndAa9hVph/d77a/p/9DQZXRwtTprSzaUw8Z4PBI3R5pjap8bmtuYfQ8J
E4S3PLUzTMMMQd1+73wDsrtl76nTLkd9Fym9CVu5nniKi0Dc6LqrRt3UYBxCvHpm
BhFrN/kjnW8dgH+aj05MkTJoI9SYO2EVFRS4hvubYTB5sAuspgqd4ZddX41HAyFq
HBnlyLZCEL2r9WTo8Sy5xZKZPYZ4rqgW7WWIVeOa/hLYfsY4li1geyoWa4olCMae
4W1kyuA3P4Amz7veKorGNKT+yySqpDgwPMzm5+W/nkfFqHzNoJ56fzSHOpnwiQC6
609rXCYuxyegzaYekKvcvBd5rDAkmK84kULacA3nc+oEnsbaRkkPu1yniD2frIlI
jyjTa1DrJgEPLJeLmhecwd0hXzoN1UQO2Y3da0ICTjN1msAUo9Dkv/WGghxb59sc
phCSYmzqckgw9wWLU9enkhbf2kiG8qD558ogEFGR3U+6/8HxfzDjA1S6qxf/dPNJ
75WPS5phK7ieJG5MoHO12kP+ij5GwjKNNj1x0yuGnnGA0AIeLaZ0yMpDmNuNLgnG
gxphC1V0KcJXynxqE334UCgaFoP9lTnDPvy+MoY+bKPfgrt7fEfujAvnyqMW5hAP
eoGPQYXp30mWy3X9LscEnoz5WXplm06ev+0C5FxtAwIRLD5M9DhO6JZC56nFExI9
rxfsac8Y5GAQzNgD46kV8YgbisrWmp0cbWC+l/W6NdnlUZUgcCfNH/GI8e02sXR4
sZCzbBUxwoPJD++yxDFv+tEryXP9/AtkYQCTBOTpc5InMjbS5TxyDkmBbC1a9MwF
vTxt0GYiAl90ZCoItTPAycXS1MMQYSB4gcNBsB4aI5xxVdOp8poF01ipTzNacYXB
XYeMVqjUWxLvmiJrY+Xy7pkz/gbqT7Ue/oKROpqSIBAWWnt9MNvkejnkODZ0afWR
icEhmX3AF2aG9iA13WMaNSg87UrMj84AZYvHHkdVovbHXygxBGcitdLWWfLBMOv8
x2KGR5h2IRaFY8iNpjjuYZPy2uivbxyXMuvGAnM77YCs1RUTP/+sG0d7uEC9UvIS
Tv/w37BUXSBVb90XFs7dVQHZFqOP4c/3vAHOOhn7VdzP+wW7EicvRFfLaZJh62IE
ypyJFITUuWdZ1oVjKQO3mS8Wx6KBdkISopL9CKToGzVGTeiJidNLRs+b7NEBnhFE
/1N+5OODzOhoIEGcptvj5youGMOIJG9pOelyfPBwRNpzc0M9x5y18/t13wbgpmwT
H2RFzBTMUudmSWfT2/HOdpUWtsFvoXel7QIdghzrtBwkucyp3TWODcYuPmw61CfD
G/bdPzdSbewy/1qhY3Eh499MBhxJMrMyKPRHUFxjQ13IpcwDh0+yI5tfKwZC7RWp
rXIVJhdlyaD9y1hyYofCVKwzmLIn0wKzmeZJ/BpqkEjNwLCSrncTWGVfSAEv1uSG
4QLTwIdDyNesFQS552Pb971axs8fugoY8PNyFSGomjl1plx4RHTMwFUgUMyuLJ4B
0UDsB9f8dqhKtxjwAsGwitCBA7gmmuofGWQFhmDvHnlg2wb2IwW7kcDIN7ghgBYo
2jyx9FM89HWyTmQ1JsOQvGuVx1pIWMMxpNFaEBgfl987xALtdgf6+mp/vmEYVQ3t
v6sZHEWSEo7NRXrbpnKmOX31HnaGVw1faGMTWzzyO3G8dhvsxItW+wVktA/Hetyt
WGO7Z/M840oQLUgQLb9v6g4liIf7tBb53RimG5ll+PsRWsdWhOgXDAcMOh4DdEKQ
0oMBJHSHGa8CVTYLR6Mn5krDRIQsn6vhGk+GdEoDlO+nxjimmazoObqr1odh6NHS
U1Ed1eQtQ7tEwOUONVhjcyF1T1+VbGolYD+38EulILKdw17jsB4rOS0WZlnABdSj
rM+6jVwWbUQUXR1j8EwKip7Dj8UEPf+5u/Pm20BgxKj81zILLNi6/XJ0FBkq+c77
u9/Yqnu+yfW14cVJniRdHkiiIfPHhCnJ398rThMvwmR5GQSnVGlzbdsV5YQljTH8
/MyN82f9KdicvNiYbMzQ7YQrueFDH/1cQTOaUw41NDEs2PsVvX6gWFEuwIZx6c2v
DQ5MgHFD5A5yGhXQzNBkahBVMuez5CtK+H5B5nYfl5jy5/iG7nwUdNEJ2vEbjiE0
WsXESI/3vf0Yy2BSLvK7C2Ve2D3tzGzx2ceOBQ34Lczyc8wu8gMpInDewuhklpSv
AUTlffLs34+4VBl6ng4y7uc1DJbaocMmd6EIC18NPHytX5CYFSXw2vVd3424A0yY
1jB/h9KK0+xYjE/TPeD1fjOMSSHoiOAtv6qB6u51n/tpaqkc3ZPm0rpEYA7DqioI
I7fkvnDQvNyvPPtR08SYheZjyjnJPijExQjV0DJtwU9Vy39SpzZ+HOAmoDkQPCE9
0qJwwI/GKxSU1fGholc77k9ukubnRYxx9gevt12Afy1n03cEEKraahbmi4yeoHBe
HmvgkyNLPxAg6bfrVkNa+GAKYfdgrKejHOrg3a5IsW0ZbblzJC58hMUYngY5bIM+
L2EzjFDqTyBSjjDj8JA829IanXYCNhfeG4EQ9I/+3hdFfqQ6yjDYcH7lAWD6rNvP
3ykjb/PwBDaJKPmdOAg0lAOcXBjoyqn6wyIoBzhqLqf+gJxy/eosmSQuroeEXk9g
F7dHS0YKl2LPtY4WvDlYPNj81H17PHhb5NpVpwrFQ2UYiAKBCiF0jVFNuyOd0Pgs
Q2tD/T/UezbWml4lQQ0F3U174L4zf01SYCxthPfMsbo0qgHG7zagAQ1nJSvheid8
Mo9K/hcaGSXE0RfXhj3BCEgIpawXGu//eMJOCo8in8gBLGwUE/BCWKI3bUY9W2DE
seqI82iH4d8w+t677/OZLeCA+9bI4+4UsKrrkdL9iRVKo24rDl9ozKMNroUnFSYq
o2UGJ1z15CwSnTAS3R1oTalhxXB/KyMyRetqNvSBjlkAChuEP1yOe/+GnPGHsCxy
LYw+/5iiF1xdcv0rkZgzt18KKgDJ/Tb8OOQ74e9mmgtk8/aO5Ir1XLRHPphpUtY2
eRovGa1x1APHbNTG0tj//YC3hwbyH5BYmmSjjloWKBJx0ekUQdH/IyJimus2wByO
DUFMlfdYAlrqVFx/vmzUEceqcQRPHWedraCrCdiqYasFWV0Y4V0j8MNNw6+SdcBV
XbPjhXRW9BwlI9mdWnemO74b07dv5bBJWux+9FR9iLHMwHjuho2SLaZcI7auUZyi
xSgGJlngsRWIKuJ2XxBrN1kvE1u+03c16wyse/cPfGRK/YKTWUvsAPeaFQZrzL5r
2PckajQV0fT+2HCwSdAhGzr8SOlJP9YdZWxevPt16I32oYsaGaX0hFavy3v44xCZ
O9jW7EGIwZLXFUIBWZax9mg/PQiwBDEshRARYW5BIWa4ZVzEEkASkpnGoSfJCC0g
ygUpJ7TCgfO8q5fAwQhlnxoE1UXikBU3lHN+bfE7+rUN6115bitdos4ceZaUxu3Y
Dqp+Tb2jc3eOonjEl7T9HWBUlRHvfHtLuDjK41wapREJWVa4zbRN7bV6JH2M6bVw
aNBA6gph/yrQUkSjJGM+70lMppkM1qvFL0WVs3lgggs0uRP799bBzEQT1IXkduke
7XZ/reND3ojfOKOSSd4aqLF1XHN72jWFOFYA3M4H+BMCfllfgB1t9HSCL0pe4cQD
9uopKZ7SAOakWKE4NUCTTKqwfm1mcFzTTQ0aUyTPFaadZBYw0L6zYy1fWGPOE7Ws
N41Tjcri8qVq6RQYhLmJcttIOLMKCOdYcKvvrChac5M7s/WuEImMcBKmAx6iz8IJ
zBXuhga98wmSg/haAzYOXXd9JxWjsXshnKTuoOHb82mGqDHSQjsJYbZu+KD3WuQv
7PQs8TcaKB5kJj3q6ECtRvVJkZgIFZqAFBHKJIdt2UyoqizsdYQwZ8uN3DCABZ8/
hma/n9WgGHWeALGdAwYHaXOwzlHMXBMyFFeryDqMKVawPP6k462Y8uOMa3ZZa0zY
csyNAVhDtE80Dx4FiM9PaOcncr1vK00nhnz2iRrdwcOwnTenaEcI6zBcATJE6JOZ
ZagcqG+DYvb98I9NEyngNVzPs0j1d2FUCRyQulm3oHC6Lx2PKw4QqL/JiZ57Z61l
XFokQHyOV4PbdHEcPfeeq4cmhjwV0klPpwxCtf/+9eFnutU8NUqgElWeJR6ojxOA
x1t/dT2AAvebY79tUdPrxPU0mA6bUUqQBG15wA1XhX+tp8DnyIg+srnZoU9mL4lp
aSo4cKG009Q5hDsyFGMCMgfXfBhqzHTit71Ei2/pk6LeCRGy8kSfM1K5TOL8P770
IdLs1Ql4f1E7yG176In0juW/4YXbpyURbcODUEk8LkHtoseMvmN7qW2S4gltYkoa
wDGQp9IUZjZ/vAl81ntndu2YO1sRaxmUYuiAgaWKNpS6lgJPpaBzVp3NNs0CQLMl
Zr8FxpNvuE56aqtYoEDH+9EFw6NwCRDMgQ+c7gQK275gGRaquy9ej+8vv+T5WXkM
IMkN6B5Y0NwFWCA1AJf8jS249Gpuc6EKDHUZH8fCdBiuDO2Vd1pNVat3MZZ4y8Bj
PVBqdhm8kuAvvN4auQTzrnv3tL1HDg5DIVsT3EzC1NlhvW8iJxXTaEQhmXNvTgP8
rDk3Wp1EQ4brNyCOzJyabx+n+u5MUOvejVLmJa4qL82ZTluXsHae+g7eBYzT/4Tn
yXbY9WcJUvQF+fVOQSgrkT5xHff8yrtL7qIl0t303+cXlG+CxVh3gDn7pHzAHKSl
RP+VZqq6vfjmX1G9WHa66N+kNwdjCpKS/Y/ribX3IH4Stj0ivo/T3g/lsY2XwuJd
WkWEhy096ZzJ6Ey7VpLP+hL2AnjkjhpRJv68P8eAaScoXOtzK4I35MUI3EVoCnMS
QvQr/3KNtyZh59VzCSqp2iyHgr8S3T0smYfbxjFaGDuVC+gZtr5wLfY5fvxK2D74
THjUzFGEnuDF3bjOYGyBfyYDu7ri9PEh1zzoVqe1vz/QgithfeycqGJw/6E/EC5Q
lI1gW8ZXRUOZg7jg0j64hOAW/9ykobkKqfaJgBxnK70OGlUw/SySQl3/S9xMXASb
91IEJ4XTXGdHtJ8mObw+0LwQzYGBQN1CelLZ6CLElbooGBIsdjfTiXnxcw4LoK+H
zk+dinoXnPLpT62Z8fJaLHcmPgsXfV7HTLI0LE1ZfTbtQAOIZfOhhRLjwNRF6Kq/
GEwT84ce2qXx11gyKyEsEP75Vbw175LjgKFTCoe2b2l5h+3ZPXUeSMXWXFibuh6B
iimx59RtCzlhsFvlCarrkqsw4iNHTP7vN70XfsJ49aZixTarNMNYPV/jOSI7FF6H
IwYfg+Pyb0p2hrwcvDKXF7gedaqLivBBWaxuzbUeaN68yqpINqmq0r6TFU3Tq86/
wT53z7rbgnxzisyE415MABlCJfPBjL0jK7e+lM9Tp+zC+trxljKy+zdlw4iTWOeE
E4xcK80TzvnlHiTnCMYz9TloqvrHvzrbynoy1h4zgqUsVsGbGuNNBaQrZqB4KQTD
W+PLfFZPC2FQDTin+BRMjOlTm6QYkyhcRxeCHq/Uhd8wpsbbQX6FJpzVQfs81JZC
ur/5e6h1xMtmE8cWWYuXTxwG25deBkD3gsV1iL40uGPbqqey8y8lAMZfizBogRLs
Sejs76PNVfdAa+uf/xhpI3JBKOb1OsV+XqZ7z9a9bxk945W96qNQtCR/uN79XiIp
60rqWuzS9Rdi7wOHCatYshquDmv1ThCkPGtNcslBG20W2kVaW8y0LhpiC8h8mppU
7QVIpDUZZzLeY+M9p00fzo9376xan+9Q4/UoX8pdzM2zEu3xD+djn9gIXrY5WYE1
eRaNKBH9Pf6Vox6tWbbaQP6+G0+TRZKl7xhGcswyVkjE3AaTYX/oY8MSY2d5bFxs
IZJ1aqgO8LrKlLUuogo+8S7qxcBrMVZ358LHKL4/1V8MfxbdKGl2aRrr54yzTobl
siNQppg+XC1cbfi2/gcfDHoitZEoTADH9tSsprNs90N1ael1b9lcH+LOmenlJLjX
RPbJBXp2aeLnYdC3K1cQOX4BEIko1zgWOEgs8YwsdMDRwOrkSdb4UxPwqKKfROk1
IPDYSXq2pUnUPHeEhZ6tjdVUcD+IGI4oCWgpJN//qhumVxOo3tSG8jjXYGFn7yhT
yIgTG9RGiqx/kwAP9jQ1rL51zBXHJVpdpACl+9yWjHoZKn/hH6gfLTbLgAkK1tnH
g3Ca6mPxPpGf6KGaLDJ0aM57dmYpAU62mpabDc0LWbag6+wxMRraZObhPQxkY+0r
gGewRp3EhGdljqkE943ux+DPu2zWS+oWiFcH5vx4r2huiKBD+xiIPBHswhFN29Qm
70Lwgr7DW+2o40v12j0FoIhZxJYrOdg+Z2xEWK6QUb2ngiXPfYgV4kVQMtb4TaSX
YI8rmC2ThRvaeQ7HntQPqQVwkmE6zslmMh1YWfADBV9SW7cP1JLu2dswE1d1XGeO
eWjK0gApIpPNWuhZ0IK/Nbc89VABYnRsWJUkogRXUibCwfA+yntsSNCgh4ufTNDX
6Mdzd/u0L2gwIh41EShbUmb5ECJgawEXHZ6C42e/x4Cg/LWAOkauZ73bxe8cpYiR
7qwhoiciuEPzMWVSsLVxeQeE+YYzIibQF0+3UHEjpkFHQrRxFv8owNEGoQEiil4j
Pj/RLzVfdiorOhtNjyXZp9BzQuVNQKXYegFUyrsCn6kmMfrsFanKPd87Pz8qf4Ka
Jk26LEFPVsNK66ChAbBqFI9xWcCiF+qzRCyner/LNxtSZC0vjI0qvEOo6BLVoRtO
h5gg+63MEff00+an+T9goWWug8krE/LUtFQ0/SEWXy/hlctK1VgQCLZTi1DYQUh4
bjHHnM8IIOIX6+xOYNuLKvdoY6psAnJy/xrzzZYMtJN5BqKPLpGcsl3/D+s14N2I
NgaizUtIwnHKvauIMss+ZDl72ELKMo9qPyJh0qr0CnEabyDb74ysEiFfY95D31To
97KG5RD2EDaP49waAChWfbjeGq0oCcorn5yw5b/qn8ynALVrUrAgvxeatVVipUew
N92ekdJCAmt1CPLdBvvM+xzLd/8PJI0UUUUDRrZMUw6NgsNrdPzb5uYGwEFoG4jh
hB62fbzihPpZIwbVKg52YPJULh4bbOyt+/LeCX+MCIwM/5SaorH9Ii64lwt/h4Hi
XEi0+atPjpcHHFx68TVRY4h4R+SlhC/mfN0+eavRWvJ5zx3L8J/2AwOMQ6UU2BQd
BXQN5u3W1cMLcIQ8UqFAtHInEBTW5muToNiJQGmqo7ypYxm15kUX4KDGweG95BCS
+5x9TyeSzwYk4yCWV4TsBia0rEJKJWP2sHvmByRRnYxJkxx3sev5ZbAepKTsaUgO
ZFciyBRRsL9GKs/BivO+OUltLeNoUvj6H5op/KC/Ut7em9arbsRQMmx1Fp7Y/J9y
1/XKTITmsxJIAT0Jw7QR1eeI+22dfRXBYuifpUCxV7I0shsLc88h/HQF3caekqfc
Hk+p1sw1sw4m+E6ZRx1cHJgGE5/kWlDZ7CzHK3ml5y9tlPlsD2BmheMKPsut77FK
rzvWzgPXm7ggsOC/hud6ofCFTH5oHRXFLFXNrAvwrh27Y0QN8doxK35lYjVy/Dh1
8p5vFmuszVs1xyoPlP8g/JKqzABkpxdGPykZlvRssXvz+4xSG1wZjo7po8aPgPID
rd3qhV16ssAyqNT8YbL4feTazyXBndhIxH1ofmHNvCH7WkAbzVh4CAugKRE/46QU
MDDR6lDpbBdUNeC61LekQ+78Ypv164QkUZkuL+mOrVrk8/wAuyFSTdW4HOK9v9qJ
qDoFxiunBHjiZNCBHmxo3v16cRIh6m2rE/4qrk77CvyQTCLLUoLj1UGbib2M0zY4
T7RyZyaBpUDs/zMr6wWguBy8n4+DGBBIHGzTUZXOZ5AUSpXd/8dWSyuTiBUfBFaW
m4HgVfTPQnkHoO9t+2Q6z6zuSfjKUiS4sVOcGbP+eWAWlaRrbAtZ3MOfUqgy7AGZ
KGaiFjO+OYvmuEaHB3qSm/xLYvMrBFEFeBQe0BGX4GkTCRIas08lQf5Ce/E1Ug6A
UgQhfZbakI3ZH16cGbkkWINPvi/2Q7ILnQmwKcZRS5Ng7LxpWs6pBPTurvTzd9Am
9UsypR5lylx6BluHr2LVl1fpqhW6AJ7tsbvUauj/pEhM21DHxr/Aueq6bbLmMFsJ
XjPlwDOX14eQ+7370X+gPkgf4oDIXXRHpM0+jXikyAvUcHetPnPwaf9EUkn0Dmz1
HrF/Zoc56BFDMjF6qNCNDzxdKEZ5geF9Rr4EfioX9XXk5Wjfs0thsrOL7wNpcMin
4R6VMrGJHk/M7lx5cPWpBSQX8fjill66x5bI1fIJUFigJ/10uRm+NcPto6Q5+DCl
8SmIvxZJagNUJFTkwAw+bfTiV5ioSz8pOCnV7rnLXaesrSRPwpdOqWP0m5Bson95
njcOhMBgYZvO9v/U0mn96RXA1wI1Hs8EthC/G9O9OWK2H1fyMgzuSftErep76j2M
5JuI8BCQvTCCzKeOy2MWqGRL2Lk2xR4Ye71jBIoxRZpmiMf+SyX7dwBDIKSS7Bvn
Y/3rlQh12BGYmnGFxTzC3kQmIS6OGojh9mnYa8zBR1C2iHYNz/RKCF7xydU8GpVG
RV4cd2PuF841k3xZaiNXOz97eEUdURSbiTVOu/brtMnix6k9BOvJvqJF4qBfURop
LH5i8ARHZEGhvBGR8vkDLnHxH8FHxFlH//sQT3Qi9GVJ0MQPpYz5rwvv5/J0MKOg
7qrgIC2bhM6U5M4apxl3bjmf5vn8soWKFWVXeYns9/brFMzSBBFq19P5+WKBbSDX
d7ImMDklPEPwa8QW6jKNFGgZp2MHmjsq3kzMCQYR0lF6p5AeKRP3X6UnoxiBbMMt
lzxAlvjCe5rCXrd4Ki/8VPyIdFsY52T7YzHJjqm97HImxplEnImyecForbI8mN/Y
Hdymx8jnRIMWc9NHlHtPM2N6xnEpLaukGJ8lV5Gu4zoqdof4wsldikXWt/1o4qmn
vbcUNUT6TVOiwxZi46koN7/LneMNziVZbUeFMZC/AeK+O3uAHxoiBDIG3QkTm/Nr
qbiFiJ4ZFCAQ8EyKVfkTRzOskQb+1WXknLznfFaCT3CIIhPzn7EG8Nztom67y6a4
Ul8i4vpSLaMsALps7hIo63Q3+qo1im8bP88jMtxhZS4Vu9G0Qv9guRA7bpdd2tvO
mbBQsX+hSUsWJGEYzMNcjD3vIeFwBh+cLoCjQDDa0G+o7yJTAwC/9gY97067w2Ei
/hnaR+CcUowT89kNwhmxqftOC2pfG6fcDwlpb+K/bud9CxZTaEzfWeUTW6zdVfJt
FspTxch4ld6lzCe+74KveYgNZT6gUdHFJyeCs6zSh+w4ndWeNDpiBlAVKeGmZ2cQ
kgneniG4TgB9pKd3bWQDCz882+wrDaQCoVb6dA7yVY6zjlbXROWwh57IPp3K/Xbw
9DThs7eG3pjo1LP5jbMYYMFOH+b9CQxZnyIByrpiVaWmmkleyp3gxWUdbeJ9afr9
XPaD9reGoG1SC0vfXRxyJyWLLN7LtANsFiIkOfWeQNmfMwE3xP7paqPqnM5PEizr
/VSiiUOdz3lZDDmVUEFUyVE2yWFsTpZ5Auzr8nfOYft9uoCWLome967dubkcgO2P
vYm2Rcils3FE42jOwHFGEwEkrLXD9+1HdU40lxyRRvh6W8opSFS/07QDU4jrG2KI
e5d3XlxYkDvP04cNI6U0ncKGgDbE8QoeXg7/JH9n93xmSQVQzBow2YP4DSTwI4LE
Wllsu+IxVmzK4cMc26UTZIxmMuGV5tP7vVC8r9MouPMAHA9a9qAOLggxD79OPvh6
514Hc7GxKiHOAVeP5o06Tom0q/S8mja0O4Pwd3uEPML3z3F95M76f0R2y1X/w+dy
yqQJCmMt8dQf44Gkz7XV31c11C1yu9QZ0KefHHt6wTOgeiTO1ngmEWA91CIZkcgw
zdvC0nti4G2TWBZwqolYyZhEHaBp54a+NfpfjAU9vTUoR0tyBFXsEsq9PmaakFbn
QMjPxhMaixaF9Nb2Y1pGVAuHYw6i8gsUOHEWnXWI6s6Z+bBXWPgUQC9CAvcoak2I
Qa54AO0BU+kQ3b0FK7AvnMPvEs9GvzKSpnN9YFIOgFwwaQ9md7EUzK82YGAmRoVY
gJsAcSENbkcpmlOZ9//tRz05GaxfTEH7h+f3bpaESht7ChCM37a5He5QBKxo66iZ
m9eQQbArZG+lOS2VaXjyk8hZl5tvP4uhGYfN9N/hO/3UdzeYSL3SjaMSnKR08zym
PwUPl1G0YKxbE3bSGdO832QYq7i2qK5LPEWEB8EcllcObcdKjN3MZWOlk9qGYXn6
Yk54drPQQxfbYkIuOFFmVUgFpcAsP30ciqoMrzU1l4IFG5oBI3smIbQgMtk+lopP
GVVqLGdMxma88pZ5GnzPJkKt8MvZh0nEePXSLm8EWXw2zOQiarVZcesWRmxrczD5
MgY9G8agjpEyy9O7gGu8tKAclLIkx+pEWzF+y9aSq5r+C3O/t3l2n6Rq1m0Zt3BT
9o7kjkbbklqt4LS2jpx43tDFnm9mHA9NNPFHDSAgf3iIMplNvEpFeQvG4XDXfjB9
p9LedgsBrFh4a6ARmPwqi9RE7ar58QTHptWLmxHFu/yEmJxQvSl9PpV4fI4rsXCt
2ARZlnmyyYTrM2COxPlY0Q3gn0fTZ/ABNZr2CHj2MlfSI0H/tI9rKlIh2e3qO5K7
wdxdhn1GGvp70eNA7+TvsByoDcJJlKFQ6QNz7xrwu2hUzuWXEcyXlLbm+IEjMiTh
X9s1q15PMBjbSks9ZSTPc3BNdZQjwdalUJ60Maf5j5aJkPKhHTHw7A83X+5DKeA7
sbgbPRFX3fWurddfGul7HkiETzZjbOT214TaCdkb4xkc3qS29j2ENe56pNsTi1id
4mx29FE17W33mVLTc4rNwjTVcQMY8V2GLt5efyU6P9DRbCSDVY5+C3uV9bY2U4RW
BvPhg2ke+WTx4Pi7qQCITyruTtjPJKiq+L2OnmV7msUrUViM+c8CgXiYNsyntgZ+
xV4aFf/jGXKdHKKhiQMGm+5pm6Eapq2qNQ9r1VC+qQlgGbODIpQ4AERxXNJoVClY
ROxkwNs40q8Li6bAQutxTLt2DHE9ItiL8ir0mSppsjTrj9VoJ3l37DdEtVogsdTg
Lw5CdM6SFzNfwjP7siBikK1svS7IoDuzwisQTBHyK8JxPdHhxvHp1dHFT5G803Ay
zzVEGkuqKur2DExl4RjZZ7fPL5BSqkNIWkHpNV28TBMOHSMBUJmqu5YVrz0RdkFu
DaYq+Fg727uArzbJGCIA84HFlNlAbTY6YMwPGyYqle/usSRLx9pPDx9rOkuCOZ4Q
NuV6WN5dPnAnQJBdefWV2ekDaXzUq9zZol9SN6CtmPTvzZNIRLxO4UUret6j1+Ok
STmdlXj1m/1eteU4MEJSDbC8NKsMKZITKm9jWH/0BfL3srViUBNTI11B+K5xhpdH
1ARi1a8guvyTZqNZS5GVB/ermOQK9l7Z6Wkis/OPXS3XxFbBP1d6Lz3QNbl+gEDg
+RTkfOXn8XsoKDYWt984afxxLsejGqa0apIBuOjvBuUO6GfNGkBdF3BrmhHZJ9Wu
AujkU7mXAWQYbBo/vujfrimUQKtThtQ0lag7FMZT8jPhNlV4sl/lisitPWYhrA39
S+RtF8v/Et25P36gK/hzG4uH9M9DjX5ER9X7+KADuqA1hEzAU5aJWSv1Kj3J9dCv
J4od+Ot/jj3vpgrv/1M/b5/azhGcPx/9nZky4pQKqxpNcPJLLzenbgHsGTPTPclj
VblAcHx8cX7zGBs/AxtIhHuaGDRv9t1/34hnAweM7EQIKNc5aa1zcyVbVncHLY14
uwW0EfdZ2FgvpzbwAjVeb2/WIQZa1kHc/c9K5iGKhsSpo4FrivZWS4KefFDqOJ/K
SdKEtkwvM1XZQxALSijJPLJ/YchbzCUBYv1FVdfDhBV24bWRxn9UTo2fn+9MMcqN
i5og2bMYI//fKi8uglgpbOocJR+kq8Dxp+N8zr3v5CXGOUlg1DWVfvnOWTP/IM4p
h4/ZqryIxqBK2/haWvYZcaytcKCCGIXmZKAIhYPtBg/LE/6GkfSaoJFD7jheGjTi
FBG6egQkZw2RpHVtIk4mKlTFUUPunTHa4iOCI9rsTacKVUS1FSqlxMnRi2f60vGi
6Cj/7s0kbr7KNy20XO+e3urtxQpjcmy3CG0P2RWoONpDRCJMsbkz5Wa8c5I0NxLl
M8Gbdmm+sqV4FfmzcLoiLogM3NHrBvocPHTNBVEYI/l1SPRkhjwAWavtZK9iJ6gH
OpqmGGlnza/kAY+7+JFi1A7Mi6MeQ1Gb51JHBtww1fzuEB/mZOrBMFJjR/GVCWvQ
Nl3/tK9z4Q0cSWriK+epwJEyTHV5J5+RPVc2sfZUerJArJl2sjfyLygqZDqXfMn8
2bv1lFMs591QFojIUcP6ZpJXUOx2F5D4b4rSS4NLoRN3g7Wi6CZV6ru2TQltD2G0
LcERI/krBuifHW/aR46OdrAsM91v7qwyvPYdAl64q0O5RqqrVccn1k1Vdrza097b
DjvYQgZdjKC7E+zZMEcHO1mp1Jb5NIguHDD+I43mx5SZdyDnv9cxS+Avoh4vT8Gm
gYWnQHUmSigEzgKfO25+gQNg5sVY/Uu0GEWnUJCtZ9W4IkE/bwQfOJvxYqTH3U6b
icdwtIA8QIuN+d4f57ylTlfKVzIRnoU09L7xAvvGHoKEbfqjD/aZTpqJbugQvo8L
CHg4FrYCxb0gwFNXr6SDyqSsxbBPBrZxUHLm7vRqUyLu/hGEw9YQM7ng6QNRLI7O
/J9nCAaXjElKJIyWIhOCywbmdFU85TPUpLJEuk8W5MXoE9A4JV54VA0qz6ByW4x/
L/EtBRsDG4cxFDOfvVspfzICOTufuA1CQoxJXc+86kZGrfFWbM3gVQCixiuSXbfG
e69+IW2owGA/v5QSM6nVzAS7HB8DD7PDhyyCrO42ySC4VwGbrFlBGWMepbwBzGOd
dLMb0QSchWfaagf1/psM+RGStFxsz8l4s/98GUD/gGOO13WYPzD2bZLg/gTmdpcz
1+kD23F5pwPTVH4V+yS1drXXzTIDttdF9gclrVgH3KxNlw17MBfYaiDuKA3/QvQn
Wo/AeqLTnDtOaQOYMYXx5edWIbRjY73e3Ayu71M5NvS9aWWm59AfVguQId/cOP9/
VTYIvNCsRzQ3h/sQxjXpKMoVuxc98LTPX0qkuRf1DGquaOWSpRNRwkcT4DzdQyyZ
7ggmqt/W74Lhiefm+8wGdtlskhTGjxmASxc9IvCheyB4lxV2y8HQRDvRDG53Qn3r
YPXZwzDWSUHNeGuOPs2NjLc4qG1ZCfUHSl9pBrbuwSEGzQabslBKRz3WoDFZuAyJ
0vWIdWTrWeQ5YaXJgPAebkLy/nyYFT3i141Pxccw/Gj9cWCruT/GLW0xF2DuM+aN
sMz0e+NeZ3JJcComfIfxC/iQcouCxZJ/GyTrP0aQ8gn35MiZ+KS8AYS89mlYBs+e
RIcEG/kGj56t+CVMa7Ladmczxq64p1JypCtTeO7+vLKdr7ouv8B8BAuu7r6pOFTP
LAgKzhvYNkL9dZe04ISqZjFn5BSJGu70NtOBGEhLftf1H3dCzNhW0RTmYHqrFFry
lbzzuUAsbrBMZijYEz/vqvXG4tiYeGV8nhfWoXDUwwNV98VuwoL9/NvRCyrtOB2z
g7DBVUHhQp6AW4J9pU1UXMnccq9OTqwLZeJLWrLl1/qYMZsMPwszX5EKdqDXwUUw
p4IL5M4E5kHbcAejt2ZXY3qij584KUV+yHy+eL7g11UQyrH/tdO58JmnqLZkcmk/
ppYHOR9i1cn79yXbz7NV690RRVXfWYEMgN+u2eVYcIiBzXeMpukzOiQOj+PN7xDM
jsGCXcrKVLb2PrjzEzc/v7yXibEkdx692wmRg0Zm16Yp3CrD0Fqu5G3WnISUS4cw
u26nCHVcM95rhr+qhcr6cIfnf8HmsY9YuN2s2WGpoKTTllH6Ql9d624eJorjK4MV
xKLmmdB8Is93eQzZazKK7UtyOysaXZHidFp3rjANBrTHZfVYoA91UmX6pPmRELuF
uq8KomMaGhm0bSWcKOeokuUaoHmlS5RcyE7yumIcVZoFVw6efjdwYZci3Jdphfav
SDKuLEZnjBiOabKmUoHm/F5AG4iHlzGrLTQxSYrVqMo5NzSBb8SNacRhgRg2RduL
xAav4hzk92MNrrQwnmA9piO1XUnVlu29JubaOmMTSVgRajIIeDVTcbH+fHzyiy2X
Ml5mxh5ekB5O6B4FbsOH6mbQkyQH3AnarF9JZ0v7ThLBKTKC9tpvuAu7jN2F82le
TKBpvO8N24BX/BMms5apqaOb+FPj2c8SC+C100axaR8xvtYZlmjwHX4i7K6nUqYj
sUYzWSfb6IWC0MdqUSJ2HQvdJ4lDEdXKD5wkV6IUSSAsPzIJybvNCkOOew3MnBBR
Ra0uQKumS2pNkJ85iHfNHJLJSU/Gm/uvqDeuDl5e3D2Uo/Hyvuc6XaKHVp99Q9Jo
CzMxs4vZFw+ZuUyF8jEEsMZgkOex/pTX48ASt6BWqhK5VBNn/e0tXqyuiH1K1rcy
R06OFpUZsKmNoXVmNNM68fX9kk96LN1z/qioJR3SOxciW7gPPQEUK1QAHlJojU7X
Ml0s0kZgHBGDSLquBTUEpDZjBDIXqQY8wfg3JjZz5VMLZ6WVRgNE9hUw+PgpGSTH
Yz8WkVGYv/PplBxR29liYpdRPWbty08OEu8Gq5//QVTALPYRMPdtsri527Pya+pF
8WiJ6GohqJf+Fj5t7nhqwaGi+yMsCJ0z1ZfyyuG2udCuASOZQDS4p9uadGPMHJdR
9+PeBqEPjXsCg0iwbRJVAoQnV9WUOUtYMAqjTSeAhxuzhaeMT2s9Avxmy6k1yOe6
0MvHWPtA5LrvYOeFtZ3qWcKmV/nbICZOn3BHTFsxjCt42pUnbvgQyRRfmDovvH6H
e7uw2MfE3IUwU0sK6jct5aG66ay39faLMoL+99HWOvBxBtU4UAPPsZmZIjLEQAth
c+sZLPbqJcjrisdJKUKN8yy/ZOAE0yR+H+l8na2MNxc39oqWE4hzXGEK7fb5Q5sd
vuS4cJ7zR4YzW+qEhFR2bJXynX9WGcvK86r9wquiG6RLZIXUW4B8opinO+yL3JDD
TMxMoQsh/BDKBAzVfz/j/3uLPbgdc0h+1gxoTp1iSro1wMt80N4sOJ3F2KO2T3Jo
SgAmsqYvGF6HkmKdGevR7d7gwdEuKlIKN4cdph7HDFtlOZjd8c5kbEgdLJBfQ2T2
SDs48P6xdkYbYvSXJ2NSrn/3/1j8bSAY4A/Ay/3coadua2w9GiV5TL+i6enHT10O
qZmMHBKc4C7MGxIiqCwJO9wDsSO+RxFrBP2zmLMOkNaifvR+EgTwl0aCgU3n1sQ8
+xDZi/pEmogXZK9RWrxvJnI703FWaipGwCw2R7jAss7Zvpi5kq8kLT09wOZxOPwT
qMDOYTnA0wH2PLm9ChMfTjxzh6R3AghS7NEwJfeU+kQDWDmzjWIHT/6ocyGsKRjm
0OXiHYy5K49j17BuEDQLRB9ZOgpqqeZpUhi4xQNIKobGdlLblPm1QJbxECL46ww0
lW0agokxBDrnXYckG6zWtzHxQnL3xTWMtRFQel2zHR2K56zdaX9AY44yZm4XQGZ+
EuhNaZifjA6fkogRHW64N9xQiaSa6N0rUD9P64IqRVw93vNX7wZFzm9YChq+0w7F
WukO2dGq1gJePxt3UQOO0CEuoDM86csABEA1uBvzBAK3oK2B4otDfjBreIuy8ddj
eNgFm0kzCzQBMJxQjb/2oqM0BhZC13Scsqrrq2jMareCpWjTPzmIsKe62A70CT6a
ckipVYSVeQdKc+u92PU4RKzZ+HX2wDLOGxxHgc64TEPH147TvnOsHmVJwUHnLLS9
r8OX7OXaifUH2mguYUe0EokiAHNdsrq5l+h4HWZvk81GB0oxU6MWg7Cde52Fj4gf
N14IQNAma6y7cp+BAJRirLRrMBj1rBU+W7gPJqpeJe6QWxP000121WC3aAVAylri
+kOdVhlbRxpGBRSd6U8uf3Xyr5iemnA076J0FIWCh9OkryqyUCAlQBKy9HeXyQpv
edKwnyxr3gBWLkZ44HfXclppRniSrzH1HtrGNmljrn9aizLEBE40o1iLqJ9p38Ob
6Dh3B7bjPuUtnt1+5/CW2bHlCrFrAslv5whJb3QgEx41asxay6zfhpdmJlcbh5r7
8uplRazfRpWuvWKhN6U+1wfIS5nvNwCVEfqJOBtjQivyhoYsmeclahP+RZWLfan8
b9tn0/Diq2zjRsUB0+HIpRPrcDbUvZuLLAWu8GBs5ggyzHbEZI4Lo4cpEjEBfr0G
SVONC0G24NP6ebBMraY49gPppxWyXeaQapJAfBVrzfiNN3n/0Hj2WSqDkSQlEe8y
QEuNVT2Q6xFpsrAUPCWmbevgCC5FTFleA2kwADL7POsi3MDd+511lNDcIb2pzAHw
VS2KCGgRPvF03AUwO1bn8VZ9fhtZh50DI8VvefQdf8LfW9+bS9LL0d2Xw9Wjpkxd
k9OZlbdSpWNYc9IGoJ+wu33KvDr1dQynq7SBGpRf22wOyx99FB2BGAi+REtMpsCx
y6VnCNzoZdB61p7YIAOQUBOHdbNG3OJW+dRCxkcPfMbSFC+5s/lnTy2Z2srsBu91
+XCWNxI1UhElLu+CyLahkttinBXwq8kia9EC3Kgj1MEWJEVu4ZAIRazTTh6kJcRn
0K5O7KFt8jAyuhMO6Af4yK4MCULMTpHnftv4w3RZAjXFJrLp0JNBaAcQmL9je56b
MSdO06U3ky6HdAq097EgjWxl1tOTo4SmV2XTdhPkDkcOkUhmyRX32Qvy3PSvbaxW
mc86njPyBXta2C5EBH8ILIefmeygghQSEJN2Lpx2r38sUrgFLLjK5htzngW9Apwg
RN6j0bwA7zZdhqyRGkN1TkeJa5Y8ft7t29SqYXWN7PTveqNot+0YPtKxnhNjfBw2
ZXmCHiq43dxjqWW/XaB/5PEUUym9I03gNVRIkvDJNAjHUwzTP4aFab32p+61jiJ3
LYkO3dWQUi5b7aGcdDJz5VaQtasvGDN98cH8fd7Xg2V1y6ngzoY3II/9wKGIXEq2
zNtmddFrShDqZ+te7fS0fSTgYN94EMZF4KR3DehSrJA9PYdy+nxBFhZ+6vQiBTPI
/X4X32Y58hiTtKUHmKuwAgegN3br7WyQLogZoCQ6kH8lzi+n1HXuohYK1N+H8cRz
9vDdnR2xqj7xB/3PatzXm7aFe+ooK4k9UNq3BjvQKImuIK3orOJHpRbxF6mq8vSi
VYqQKq+BGSeRRgTVVRIyDlZjN8avHWLAaIhBDQFli2LTNoBB3KOAXHbDrQGbM/pP
9NcShvwgSBBisyEd1XCWIIobvie9WSMBi9PLV+Wj98HbtA85EL0o4uXNLA2+IYZP
Byq63W8JXWRVSj7zDi2AqrHedLfng8uMvIOHqHNuMR/ED5T5GXUKd4p6m45Qic8S
o9sVBWRGE0uYrutyg1H+GrPHqxnzFjrJtxEJ3hSSi1hM+vXbTy15CODtzUhYprP4
QdZOQLIuOTAbj7a0KQrYwWxKpiZHQb9zjUPBbEnWjAsPG438Y/We2THrOjTef++o
0QiATtvVTKPXbF8YmmHVWYOlUBE154tcbnO3FOEYZr7qjEO+8tAUfHY68mztawUL
MccGrYW0lMsxlLVxg8zvbqsVnPxUCIfyvx//2TQyba+Y8o+DDKIIrNpS8ejgiMAQ
jUVydteSIjvGVyp3H+3hhnC+EYS10rZY24T++tVC8v8hqPCBVo9kCyGRT4xpBOnN
6FecYoXpJKQwyAW0RY+xl30mXKb/guFB3o/FQNnqr+DGAcQeh5qoOtF0OL/yjX1c
6/wOBeraGHsJ2zCY2VaVzT4g7sFgG7xGIlv8dTKqWVG2EyO9tU6XeW7EWWeCPuk4
fvPFYnI7XhOpihaWUq/WvyWQs3ZmYxKEN00T5NcI/+Q2eqhiceQObD4/sJQ6MojE
Px1gbRdsoLXk70d4zKewNXTaq2JgliJPeV6g2S6D2MSSstyZ19+xHnR6UQkI8d8e
RdQN3lgYxkP5TNzZIpfHrlwx2aOTa2ugpgdIBwQpNtIIVHhFfM4wsT3Wq3QV1ytS
5ZPYqTXAUhY+Ly+n3ci4MeLEJZ6VUdOTJyfGRN9tyHRoWQ+sg9cgD3Ndok7qxcsi
1ogKOaQPlYp+gJVNb5TPtGb+lUHarxbdW240exFKGx5aUsjMTJ013mfeOqDrzFXS
4sW6NK8LEOfNsZcJ7fF6/CzgO7akgIBitV1kGawdI7naoDvOMtLoL7NnJuLcezx2
FxKlLF4IlhnWmQ4PMjLIxGpNhNMvSfWhQtAY/TqkxFK4Cgqs1vhO9yDMrfJ+4FKR
GMWPX1rUGR+KC1TpMVFe3LTrAfD55aTXJVN7fVSjuGAxd95z7Z+HVY3YLqtFS34s
f87cK8HKlOT5OSSmPSIvPsdnyA60KANf4USZXfcScYKYjX279eRAPAR6R559Ib2I
BfYh1LunZvsL3Nn+M6Es/5DGyRp+7NAPcbuIt/DM27+yurlGbeehgjqmvsNYagw2
tlyk58kZIPMJ2V2d3W3Yx4jEsAaoTGQkbKxMEiN0pn6ttIHPhfpW26kow3cMFh6W
B71j+e75dUTaOERDBgqXcJrbQFxoA+05guJ8eD2QndjVunahVwHx6WkdDLLAnZt6
JqEYSpfrePdRU8tpKdd/nD6szz1x3k3OcZJMbfbllS6oaK2Zjwe+VmkuWZcmn9Y6
TOkJc8KTWCarZhd7MVPd8zbw0drbzfAfw3uSPxEsk7mXKGwjeLS/UC7CX2HGh1fg
Yyvo+lFKy6lAoRiGE8PQi1eipaSoEaMocVxcilq8WZ1x7HiA8L+RoAo7cY5FjUsy
vFuVUQphrrcFvjpYSvIoIfC5Rgu33h5+GmxvKCTLkYhAN6x+2ck2tyAouMUeiJo1
2c+zbbUlVU9dzGSODEKJy3gEjosy+fl62yz7nBqkUbkARitfT81/Xc3c96b4wzdW
Xqi4u8q0Uv40LnURBfoUGdyHtXB1XI1K/28KL8bnGwUPGn6IeqwA7lDShTGgNzPV
L3LRRn56Vy8skUnqeH1+SRgYZGA3RqiTGr0s0L0C3/bsCBt4l4egQmliajuurMsY
/8rQWiGRZkGYSFU1sg3dHq/An/7dBmuz2eCrCnMvcwhx1+EabDwgdkNiCoaGmDuG
vEZwvKB5+cd7yPBwvrPSZ9qS1V8dq8clXpWqbP0nIy2mE7M9KS4Y5lAl/STSzpMx
byZSipC30n+Q3z/Mmk+oBY0kXU9HFujGs3UlW2bLFW/S0C2zGL/43aEB8h/9auvk
PpQz5ePJExnHGiVJhCehqcZftuQfi0/BhS6bRVYP+K6EbkPmmaIgHCiTmvVZpU2G
qzyypRhohTrLMPOCFE0azLZgTUznQKhL8GVRUYbS0CKsJvUxWjq6az80gdgVb8iS
KXa68i0FN0VFQOQzTu+3QG5G6haLNQyzTckzc/F5/h5CbmkmN8coVDpFSX/my7zh
FpZFSoC6eYVH64oM4VsJoFyep0cqRp5oKPDjQo6RRdQKPdztQkIqUPuzK2GFVoZg
mMvaAhAdfxEyyAHrlG4rWynjzF0mCBgubwQ5f/voIGhY5Hj4G+8c/q6Jx0ilB1GX
Uq+jiq95DxdUl5NkMvi+VLzbAXtQdObQci7rupMLtVilFAgLBCZXKL80UCA+eGd9
zOLd9KAPv3rBsRf47tnZTi5WhgA10d9hMpcitLgVhW5jWeVUvMfsOjSz4I47OHN2
Vs4X8wCMBBaXVifXwm6K+3Ar1qRuzdqoHoOL9Xqsm8mD+Kfw2/PKh0WdjkM2cXqx
AjhxkepJAee/vh7xfTjFlQfIRV/24x4iq4w04sqJsS7NodJ64mwrfpmyLUd8sC7I
Z8Nm5x9V2r6DI4SpmdDhDuqj/G4Iz/0uVbPAu/YGjTt5D720IaoSRiffTsuclIKN
jYDg5mlhLVcYp9vZHONx7gnuL5vUgiatQ42R8/KFd8u91+tY3h/Ocx57A3qCAnnY
zU+APgMyTVGktEaXOLIaSgLzu7yM3z/3qiA4Kl3mNZiJmUMtQpU51tW4jXodS2O9
P9OndULgr9r0wjp4IjeJ8aXcacecyyDPjJMnaWgN8nODMlOktE6kkSi+0JT//+XQ
J3LBPVwaYPOabYZg5FN73YYVf0Xa4RjQL7WCTXj0REo4XdjFAwYASvjYs73sSmUG
S9yrpiutfI5hPi/zWlzbX4REQ5ckY3PmNE12DimrjHNT7KC0U8qTCNJA+necXjRr
4tNifpt1NXPJS1GUExe0SLhzZZjrhzqieytyJ8jCibnrGzB0jM4CfmVJTjgJkc1t
uKpXjGocRK+13qp429x406eO5htlqfOfEtj3nhqCk8KYNhwGYkfsJ7VPEd1PX4Zl
0OKzAf2rAXbYqmN6GL/ny9u62VbKUwoHZEhimATksGXEwx9CvrW3YtTRl0iQRpCa
heX5ROpxunHhDP0XJtZNBtzO4w4g7laVzpzus/qUKORqUucSScEONU1qpRw03RTH
6VJ7YjFV4C7Ch6ygsG5jpp9Wx8yMipnJFUyLvN8Iz9l8h/y86+XTCRx0EC3fJx2u
Qy/5jLimIsEoykJy5YK+0nwjNoVbHoBugionV6LrRZPhbED6juKUbo6M8QuKjgc7
9JUu/BYKuvn9Wsx4TMrYlukxY9NWFQ85keO7SXLu6z44STlYkfNC8OH0gH7eL1QS
v9CP50cAQtt9NJIzuM7tfaGzVSkcDBYImBJ4K8/qiv3zFeyzq+dlvpPBT95ytsyE
DrTg0WmSUvcVnTFXhTlrngxXfQRCZj7i5HBJYaWlS9YoZP7/id7K82QY8N5YagAK
OMBmdaz6YEr9Df/sycpV/HvU6Mz66U7bM+Lx0o1qssGbYJjrVui5xEGpV2VFiMEP
LSBkYtflDtFINe1ekccm8qbjwRQbeICRgQUwQXHszQmCk3L53smcAGP3ODpsj2z+
girnEjwpjRN+J6y5OWvOGtSjfszjWsauLWZHvTB9Dme52d8RkYAx0wZPCRK1cJYZ
WZ9mGiDXD2bKzTqLIu6RFdY5/QGFHZXm5lV8wniRseTf4J9ZP2amQ4V0Qc4xBliE
uyih5RqqsDKKIkn0eE27JHiv4Rb+fxLPq44se7LsXOuemtSxJbLpIKMTzUpqRCJy
t1GvxjZoshjkWh0lY+oiLFuCukK2QdIFWN+27SWLiiyCT4IPLbqaut8kTqiHq8O/
kGVM/EXvCI9U8UPCnRjXLAwdKpl9K2V1UJX5acqY4ZWE+kPX5s1NhE92DZ5DBVW1
4uZVpWxLzFjtc+vtXrzEyiRdbfBefeAd5juh6r8kaqBnHkWeINSfpev51eKSUmn3
n4F80AlGEVlrNWRk2pIaVlYU8ywhpQSzkktIni9QMeq6ph5P2fmP2TJ4MLrxOu6b
MvRAinN20kr7LabK1zdNrsN7x9/kuQc7C8/vrfD1snzPXIyR4OiS9t8YiHUJQNwk
azq3XjEWGXkCvTSfZZHYnKdfQiijKl+TkK01ppRe7dH8TSzmbIQcnCQHym/5MiqW
0wbnMxY5JEHtPjNy2lhsgbXx9XuplKF5Ey96MXUT8sJrlCVVQ7nwCm6Tugkwh2hU
tKf8jkx3GWrE3nOnc2LGQ3p9MNhj74LHXbYhcz3356/avvAtaowcXWUUGGI67ZPF
UqSila1d76wBIfW7asMVKMoq7gksm7HkwzSH9SGZCLjWNlqxV3rFn1CD5pkY58eW
SrJvwIEJM23suI/DgkPZkYbEwW8GkhUlLAxF6KBZik9n+b03tOZGGDPn89rbO9RY
hRoCj8mt53AFHBO0AvtRxQjkkLeFs6RXkg+4nXO0GqubrYXcyzXntPXP830II55l
0VmU13y+nZs0kdMaz4uuNL1NFl/PudsXmhpfyCcfPpWgowy3Ee1VvJ4J4zl2ukch
Sl/hudniE0q9DQzy2SIrQBYUjiuVPmUxsiORlawqoCFsoHAteqnABhj4ephhYIvF
W2L3N4YUK687Ndd1hSUjVjxWshRuq9b8IcC6mVk203GXe6IFO7NDPAFzq0rpFMJk
ZnoozRLU0tqqfPMNefQiL8CrKSSBuTMELEinOzOu5ok03AST/IoBSQACqOstVq2w
gvsSVzGjNJLpB0gmBY89saYVb6QuLjhyC1MvSs1ZaS12jT6cG2boLIc0bmjCTITu
I033MwZ6agbDSNIn+lH1LoHAG8k1btnpb7YZG+D3mQJ5GTXgeHiWkwgyuriA3SaR
XENsJkQlcoHzi+fIUHssG6IyQDzIhO1899dqD6wKyK34XBwSeVBz6B2H6gecG1FV
3eTsUe52aPXFtJmkfCJL3bhrFMmyWZusDu9xTsUFif5j/opvj//yvP8XAG6TegQw
3SRSdKI6kpSlxe1WoPb8q5jF0iX4D6tae0Ei74sLY73voPb60kFy/Q45PYWug794
8O15VspMisHOZ/ZobKK7tAmnhbuH5Z89qVETYgwh271PbpsK1Fv8895CWULbyRxV
WxmynUQ2UDmTBm1AMozJ7yiVZTx4AIiz7B7ZkTui1c4mw7cHTyBYGG9lZIRQZFGC
mUPsD/sCwi4eHSUiQTMbySGRONbOcdyv4pms7/nxcMDWkGSq6e24kPGxs8rQXHIm
XKCYK4OHKwOMGzfVg/QMk0XKb4JH5uKToL74WKSCdJk4NgUjZTaXGtn1jwwCyRh4
ohCQnjP27xmSIhSvow9riPYxvbUMx6eSae1MSN56HfeNvRagpn06IKkvfcSn7MAT
Gueg18bylLtRTLZ52Lnke+eLOI06h883Tzi21i0KsMra06NkKsad+MQalD3Cco40
KvMta14SldqwNU5188eJi4BtzlSeHCWrpt0mynpifnostGfTgYfNEr9PsfzoE5oW
6z4r8UCpKkqkFZpHxOJkYHLIxUK53wHQhCW2hulyYMMstDTEReNxNMvbaGvnvasA
JwNdXVDWRh1nMxs7qUbCL1hM2AKgcShnDBVrCgWRx/HpstmuN+y/KUQTUlcNkoQC
dR0RXLtpbhfqhmf+Z2BhmgywT6ozWrGBy3St2ZNJc2I1wXY2cTEA6YhSf5D2NMjh
BlYAC7zg4PhfrnPT5yE+8mXWHXbgWgHNbWPIfhjBFV485TzHKJzrUJT43cXeuZIJ
aIbQOfUr7ZMpUcrIKwarH8rJzOVZrtNOc8/QlcULx5mCd+iM94icZyVFbslD2VL+
9D9QSmJpdXfcIcPGvWysM4ewrqI44vHaW9xLhBHO3JqfT7MYajjrcZYtV57z93Ks
Av454vg4jKeVqJUweO7ossDHRqGkqu5iA/9v4QkVeCRl4sn1lW47c9H7sBDNKXHW
fNXe9apea707RBroyIsfsy4vUoLP+WLkFlsfZtkU6h6zs5Tua0+1mUm9fbbKSj3/
CT71zhN9yj8afiC3sr+z/JoyNCsdzWQPthBUv9ZyKdDedIXSRqZ55rPff3Hhzk50
mBEoUdZtZ3mFmQbgqUB+gELiSubxHzydJHtK5IuvSS4c03I6VN6u80U8HGq4D32a
jGwVUHZZmiiPshnkvTp5jlU15sRzDfcy9jmm6ZLQ16DvqvEkoT75dMO5pT2EQQXt
Bg52cHfZLMC1vK51m79Ra8Q4vJIbrYifxdLDlPpXL2SluZTKlJMCS8PUANfZqvIt
sSRS89Kn/xDcI2mnNkgsVeGI4zbWAARcsVSDrRIPZeAQ5XKRMvwtLZJtqQpTMG0u
2qKTKRyUyZRsmJ7azebOxwqjWfUYUamxfsOnhJRUt2afLLNARwWnp61aSNcdsUl+
TDXfzMI5Q6gPWdPvOTqG/lghKQArBWAZ2fWSvGI58FROQQsOB2b1qKDnTutbt6U9
eAJE2Wt9ddgkrfiAz2vgWGLdo8ZrQRk+0OmVd8ujjRO6yNNiuLbdDctavefVapBR
htoLFYYlrQpMLEZ4qK4w3o+eRKOW6oF2sOkCkjksGZgAQiu+D4PP71cWbMagiI20
43WkzWc1eGpHVziU/tmqqDEvYPG3cN9toPduBdp9ehGGewaZLPRjuWJPRGurDke7
BI1dtE4dR8fivhQdEwSCZKp/OzY10WASWMLgO8Y7VnkdkZDaoRX5LobDn5fkNU3/
PCfY0ELEnBwY/PnMX92nmhC6US6fj9VNz2UdBi0CApq3QzpR8/Ve0BPUO/IHKp0t
Oy2WAOpqyZ6X/uVonSI9LY/n0uEMGJVw/MNSfIFErzzaeewSey2BVVCUwRiZ2gpo
eEp09mWz4TWUTCw+hdaI+Y/tgmlkkAqVdaXJ713dgS+CPsZd7IlS8YwAStY+oc+D
p1U4EEkZTlqFL6FLjKv4S/+eaOB0uK7Fo+cOX/kuPRzfwwRv/uVGzUhDHh/S77Aw
i0GYVNeKgEhC9cz1WKzalgul+w1LzpgwDG1N/y1Dt55o50fIw1X0UBo8JuayxeCn
PDNK7wpjvHZxuwPaV0pZeYu6qWJTyWdP0r91k8QnLi+x7yO1lxp1TjTgDY/LEbSK
3gvoGQEOW9sIHI5yFQH1VpGYyRRuBlZr4JZTqot+a8zFuMKOu1YfB8NWH+Lli4sZ
iDuN5FJ1sxQ+AL0T3Wvlui370hxzFzZNOQDklmZKPFBtGmplkkDakzjeEE/Pog6I
rNhIwLXIiefD3EA1VzjbDqlLqOcbyFxQQQSEvRpeIt7GtNBsSfBkkgDuacozs2t1
r4uL4qVQJTJm2iC2PKMfQ8NGBcwb80zRKBOZWi5XXJKokTrcjoAfHDOS1fNv3vWp
TkkoOXsLcvWaHa1NXGkSp9UVxbWRHVKK5Eq7y/0EZBf6VRMHjKvpeC7PNnmfsQRy
M0VIOkDg3z0+IpWIAFDa8t2LZOEUVMKHfPj2B5M4X1/M4E3bvkAtpQ0RVNPI8gd/
mNnxkYCRuYNNZJXyYtAhGzs2AB0kOW1e6sXG3JzyjuIhaKvkWDK9IKBq5Y6z1+2G
hgstBG956vSRmBeWmna6dPA98DgsaSAz2EDvHarS5eZCsOoxo/bs6k4csI/mVVCg
0U4UQY7Dl4UPMXZpUpTvVyOAkDCmhCk2+QTSd89R+cowgbv0zQgth7SNHZAvTeTI
lnZq7HU6WUj+yuq31SBN8q8OEDW1JHzPrD3grCLDfnC76qQpxJ2OCvgA/AKOH+SJ
Ia+Y07xiGYhiVYBtFTBDhrfU/OA0ok+S5LcQ6hh/c+SGTSoPv6FwkThGYLYcBRlC
XJMVD5mYaqz5GL7Vy30txOxdajgJQ3VRtUOPi0uNvy0ov0PrnvEVOiD59tSy7o3z
Mi6rhWerIq3Q1t67H2YAHT022+jQKgIx8KLK4y7uiIrFeyoytBuIaAUQDnctFUFY
cneAXnDgLs/+/y94+vzFoqkjY8mc1pESbIUKPIMMmGY0Vr+YNktnjpAX1tk2kzxC
NC5t+GJxOYH322YevBTyxydZxJXryGeabs39jza3Z1YYOQE6Gnz1gpjkw0ugYm63
A7AulttgQrD21JqSVj+4OoizvgdRSR8eEOezUgERmTpNGc0OsAoiZPoL6ofZf/Cl
DAxzv1L9+ABeXqCkZ0MVsZmFb8Z+1e/nEQe3488H3RTQMz2XqN0fo7yef4pqPjZX
AupX0os0rkRUB0svB73Qm8ZkKhIx5YJNwnBP1O3R1TdxLOsC+j+L2Ob8W5XzUesM
/1uwk9Dh0pfj8YT6zUhUY2Lz6rduNb0ENUtCsEaoJJwPVYP5aPDUBjK7/dBV2gFj
/3e1qw0yBQgfZ9seIJIhIO8Ecf9+JTy0JX27H6f/HwRU737cwfmDJY9Ef0u/TKSn
73uqozaY0+WEa2TdOGEmIV7CrXvOH45nKwjT1o5ApIFJy4l7nKVjkLMgqRZmThMW
G19MX6JvB+U0kiXzAeCIFRGGXHDsJV/pErWpIQ5DSoWzksRI//H9seMvWNl7ejKf
8fTggC3RqDxvTIQdhXQmhGTYZqhv1Ki/LeIZBpIQHcXUcYTsI71wVwRZlJH9iP7T
CkqALacjhVjXZbcZXkjbCfHSNdaezUEnpNQbJUv9aFJHDAYWskxOiJToMxKtOleI
/GbjrbvLwxWOViFB6nx+LqdpAFaByEG3mP12sLA06X1JJHOwaaMfcYf70KXBY9gR
TLsdUFMk/TMnC31pXvhb4bdPQhVzo6d/tXbpIPriGFUftUzbTl5IsUvOmdrt4lko
4LsMPiXUA+FnSH5KvpaTsyl8ImcKiEidAHARcAv7lpsAhMfdvio9boFf/gLSDHhc
a+NUJzuUTq2yTZWNnVFQ4VhjbjoGhxRSu03ecRtl9slEjVAI0QzsVSeocB3rRC0f
rkm8Ae7FiEGWvzUaEenwgsFhQhammZnMGqcREuSOJIm293irV5T3mxOUB8WI9S/m
0coweyohJvDiDOLyCbq6UKeVThJETbST8a0d+xkSuxW2uHdEJ0k1khI8FCtgr+t7
IOYfBNtnX5u0j1zl7WXxh+AA1iKgqlGFQmy7O/8CPdZs3nBTD1pyzdj9b2Xw5j/o
aetpF+noGG+GyOwKkj22N40vcXsYEvOCiX5djEX0nIjzCVVqmDhDkM2tz6qz6O19
Y3iZPWEupmHLUourmPoxQmJjl4YQcUUNdHOtWePnfbYaAV9SID5hJ4yUELEgLJ2p
46GaDEFjkiDDUKzKHzzZB7ASkdklZ5WHJbw4dbq4y9YDDggGz5SDF9Z+htav4/+i
L5Yb7QUzgS9rH3exXT0a4b+gvVkab1ieybVjJS8hBEe3BKRDUgMr79JwRre9V4S3
4iZ7Hak0qMF1E0hzH7GGC3PD6AlJuMtPxPtboOIydspLi6NpziUVsIH+FKKVexMa
XEVAjIqTFkHjUYSgFTUTEFr7yhmecfY7k7+s7TzNZ56BzcuQCDnIDG/Gop5cnR4M
TkA48jToAePd079hS5NchVUz63DVY4cd3QhsydHH61KRl7cJwaN43AMjSOQwuLmo
YHh5LvMe8UGFM1N9kkFUR0+xa9wcDZARa4JxXxtfNMB0U0qDjWixY8EyuZWIcBvv
7gz/JQxNYrHehKlFmDQlMZ1ot7IVpgEhxtxVUZMFF6QN29+rkT2ByHuIutI8FzGM
TyFVR6UYKIRhQu9EkpoeOAFJY6zsTQ2bZqwLoAQsp28eSYG4CcxFZhROliFQu6fu
Ze+sOlpeBgYwQYHf/UqnXhkgBWNa9ZmILucjTspTsmcS/iSFse6v2c0eRECc813E
4+qvrw1OQHrAsCCQKg8d77GkdLU6qbKRqmXZZ1N2AvU9tJWG+D4KNoFUiif5VG+X
VpKJaaq5DVDwR7lG0Vf8f2MOAmbyjojPVjeg7/0leCW1mzf1bRQ5WkpPioKdtzIo
5I10dHBfpnowN1jt4ENbda1QOogwgKg0culNRqYlBuZ/lh/t/serKwfm1LSwZEGv
6Em2QAOA9TnGGyiqfhligLz4xAwS/fi8Q7+71LN0j7UCixuHtrIafQTRnJl8V9iD
555J8d0Qb3Q76pexYrgQlenf3l0fVPhl4bi1jD1RJhyUzfBhgtQSJnGwliygd9Ms
g4yGHDFCAH/wNWvclcCpdcrwF4oWVqBhDPYHaxKcYdzHgi2KC79aDqm18EEyE2Eq
xiNl/c5BlrOQgMBZ7M0DyeJDxmwnCd8ZvtkjLLYT9xAp8tBpz13ceBgWB+oAvreK
Ss8f7L3TszzZRGiWbTBxfef2aVu8Dd1egAPfFOBEpVh0kYnAsLQ3PxKkafgNynmV
lJPrKpIZnW00oipo1VfPYSzNWwfZUKIjosAF8DN7aO5BuEdSWsoojo5WeCuWaeHK
4lg2/hnsgAWsvpQ7Q+3UFH2fLdQLGYXe0xHNcmdHVKb2YRvMtBhHcW7fQZ22tmVv
HAADoSUBX7tzjq05zhq7HGZltO28x2KBu5lEKFjlstYaWBdAbpQrarOQomzo1SU+
fDn7xIVgYOB9NehzYuVHw7SD9uqdMYgTHfee98IXVUvSWsnRUOeBlgfTlUIIkSen
22VUuqx6fqcMwnP1U4b1onnCyZ3U8uk9slRzX0J4xO6sZdT/RQUERJUyF3tuowJk
eTck3TXdxHKvOhbHzlQZwFia7rfiGDbB9MKGLr/PGmkyts0+hlv+iHuR4XmrbrFT
JO4QaudoOTGBz8L9tQBGFOobHDW6DdTbX6CAdOa7+w8/8NpVIMwneo8OmFzseW2k
oaAQfDgY/qMcXxk1myichEqf7kUZySq/ZfkoLIVl7GffY/2pyZQRbzeZobd5BuRO
Q6KCpyQxd5UVmcIadLtPFt9TGaWD+iIrvtURc+qL1NgkuG7obq1cZo8sex20tO9v
SoNOCnZJ0h5hEi6xvjeZTw4xYiX2pi8ZBb7ZLjJW5HpLNZu9ZMu8zCSKMOetThFH
/C2p83eSLlWpQ7i4L6CXNGqsMy5lXn0Jr8dkucGkjCvurba6X6crOW8O2q/Xa5xf
S0RcSOTDfMFbNOmp4lby/MfGtWHWzoA4yBsskZxIyAPOrDDgJpUPsPl4rYsnS/7H
P9ml8fLFqOjBMj92xVWyREZHOC8T6Tq+GgpoJlM5iB5xgsv6cAxs6iEHNx3Ycd6H
qZIWMLcGxvmSBOdmjCfxqqC3WMlLeu2RQ4XvNGhZPYCCNPDbdpCbRmxchyj399qt
PVdsVm/RxLn/eWIU+AjfeYTDHrqQMZ+yKQXBA0K/F2N1cObr+7xIe/Yy4/EMBkuH
U/utOWrmnKPzqnh9mQXjLKQ6MJlS39mfjY5CIszpMBjVr1Ss2zE0vB/l/a0mPcDq
fu2iwnLMUx4+NfphV0h61JsZBxy2Gt30JTWv//ov9Y43oVbhko/MVDY9mTlCVGOt
TvcT1JbBKtAW1AWfqBPJadBz8q1MDUhtsynpQs5Xp56jdNIxA7AqCPRrxorT0aj4
QRgDvYeOLbpK9UuajiaJ0HiLGPpgac3W6s+EjlyoX1C7pxK/QDKyFpuvhibyGu2h
MkVJQuiJkalULJ+qHJeobhxDVOrAsJkyc+35JLbvAQrbfioPQLUpizDege1FaDwz
YGpr3uxAp0C2SThAk9rT0BQTVlk091NI2W6n7u4VU4sOPGe4911RZnAqOEG0/qP1
sCLWghWH3rCDThtEzqC/S1bGOYy2GoQA3FDfbvb7L9TCkc1YI4ysNusK+QOTFaoX
5CYxv+kHvKO50sMZhErpFYgjYL7vl5ZnzTfRI+il3Izguf5hRZ4Pp9fINyrry6T2
dycabTKUt9DIPQqxGQT6jlo8c7MqV3ODoG7Aabfw/xUDEqjDWnuAcPd7MN/Wk+8V
pkKic208CYlOoLYdV/4qZckq1tg5xFmsOVLWwBERyMXR+1scl8mzeiFSrpA5Zopf
SdkPvw96T+mdsWXOeZ3chEZjFRPUy5JMxyNyTKWCK9r48qUJjVzo2GMRB2SL2H8L
+Bs7BpcQXEYXXGpMR5kN1iXq2zrZ3/QBho+QPPQ4FMJLXPiPTOaTVOBOmkEyZD+C
R9yJzEudeEm/jLqSAljGhpDHYuVH77pciPYCm7e32rJdGbbFJe5rFdml+70QJqEr
z/z4K5t0LGExgGN0gPkCiaiVcNSn3cExoGEXsl6E3VfKrlMPNVPjQhTUKfcZipFZ
Yrueli2W5ca6VvQknmqqvhCgzNVViPQdj8ebgZXnHf4IVc3YfT71uWvsZB9UzalJ
iv9Q6V8IcXEwcVB7VEUTJnPR85DrMBHKv5AC5/n3DynT2hyYnlN6G7MMIF5SE/j0
0RXFy2uXSNK+7LfjdsM7wNbq//8ZvczDS4/pnB7Q9xRZJ6Yy17tYFipuuRe6YvtF
LUwLGG93YT8nxsZefvRfebyxTZRizYgvsjGs7ryH/sQMHqFDdGb1JFYChnbaa4lQ
aDsP0bYNmL12fU7NpI7ACdPM2T4a5Hcdj5fSslX3EHJT84SDIAGyTAxWAmCWF9XH
NybFK3mSJAbzZKJ6aMw5Te68sZCq6/wn2IY/5g5ZA0Z+UgFZGT/V+2RcNuE6O67Q
wcJb2z1m+a1jNDfvxqruOtzkWvanNw0/EMDgySFmUUvh2rZbDnlYmxSvFgb10EJs
0ozugUTF87t7WNLF5yjPQrnVXNa6xVd5KnPfHFmA2J0KOyfifpcXsL8b3z7MFf3i
5TJfHW4yuso8SXTit2ALLzg6G0DSmKvuLVx02rNu25B5bTZIZxMxm//S4Ttl/K3z
RzK90f96jxkTYy2wRaQWyh0kHkpejIGTiCrWot2qHqqHhWYU7AJwFBQfR1Cgn/7c
37TjYvZRfuqaHhCj6usus8xjVoeavJ41/fqrhfHZBFCuAQ3DMPldp+wGwqun4LhU
hO1qIgu4FU5lMCnxUEWLgckQFc3UPBK8jRLmhNEMqsa32cU2zz4frt0dnBhoVaFq
YkuobAWO8zDjdZJP5ZDiTIy42EF604pWZvadR2he0PEfCGKo3/c+CIB2sUvoqx+f
/QajJu6HOhJYOBRzSy5QJWrmTCnMLP3vlzMkxGidXCw3utwd+lkbqmY5SVXz9Ei7
alnUA4pNe0vyaJ+hJO+9MsIwmLt85Hg3YBUxlK4Q71kpp0fx0XOcWny0JINh9UYf
6f5D2kCXjxSqZ9wjwSenj706Cc88gysBLIlaIWFeRXdWp8jBNlxB9eijvqChHbhQ
VLEAIifbIbZlqW752inZUZsRiMZu4u50f5YcWNvif3hw6J6+tujIUE5bnb+PMQyN
rpJ7cVB5Nj7CToSkX8/n9gSQIc0/OAQBeWy88Re2YW+T6zRbM/XzmB8mwtLmu+le
oAOIjK9Bbds1r4mOU+2rLr88GC77SCIuKO4kGhyxU5CDdjyZ2wBQfcn9VjAK2dMa
keQvPlZxZ0nTcd6ueWFFgx+ReW5894NDD7IxZA8RPhNjxUNczBmvlzUzspgG5hwQ
3RcE+d4huGiZoDSKJPmrhBI/5RuQEB6qKuJz0h7S3qj6L64hcVvzCTNnS7iZUyU9
9qgYLoN1sU9kXwM0wRsBUVvwQLDP5EJskerhG1Cg+EprAmsxnZB4pZtuG02IBp6K
nbWTx8W0U0DgDFCNi5pUjM5bmxM8As1uu3ux+wKdXzelo6wdTUaHBxkVgwlCeJ0S
wCdc7TAzfW71+fcQansUAxNWq04L82hnqwMw6KtvInUNt1DbTTWzYW9hi1BAoZhp
k7xnbq3cdabvfv0flAeRbCHLQMmXub+Sfk6Gwos/OxB4kXFoOT27A5EIO2HSd4UO
UI4cRFR0R6TccQOdrLoyCtY08sqeGWjokRRv7ob4rxmZl/RzHoSjHXRQJInOCe8i
YRzsRSIJaZgq9GFSmZqW4ptAVCr5Lsv87E09Qq1T3h5f11gjdF1HVbP+FdlsImMh
wyk88dreZSONtCI9+7cSR/gbnrufo90bOam6ymHuXvlQVFmrNaQ8fFx/EWmV+wRF
1XnSJNfvJSf7TIH1y5labEnATcFqfKdFqzGmH00KoJWQNLdVMHMp0KHpvceZJO7L
VZDqzj07R31WsznTEv8xofNWw4K0gg0L6gKR0YOYO/4ARfGN6XU/0UnciOAugx+p
/fIEuIb9XSd9uumlEmkQPq4453Ra2C4IDaWbv3fXmuzVxIzd7tGRxhrZavfdFpLa
INaJsZxTWx3A5Y2Ju5JQB29REJFbcaXwR5lQg+gVZHuC39NrS8dWUY+JB9QL2OVh
Eo1J58KlEsfcLykqnwleYMyrJngTR4EGG9H8pENczctravNa0nx8pfwAwm8OmQhs
WbcS2VxHSZTllik4cJF6Qv90yOE78/WaJdeNVkEGT4STHNkK0iJmQynC1co1rb6K
NhxxR5Hv/IvcGmmS2vo6VXI10jZ3IK5Bi8vzrtMpRK8V80kAwUtyrUC9ESFAtvKD
ePf9OD8NVj5yx78eRF1FUyRdijuuGB7fjs56/J2dQptmUMlZ+Fg+x1j0lKjys6Fk
xku8DwRluimO3eRdhlDiqdA7XxkiN+jM4VZvLxXLnLAUBfYA6o+NmDd1/2D05nrV
1iGRqdVxQPAHC02550SEOSZEzytt+grn1sC85RrgAMtDXPRRe6SDebABwWIIBIbO
iDGY1htnh0f01316csqSqVQtBEyi31vVLG7taZbFbXzdNEgTDTb1pzHlxrFlsKJV
s2oVx/DwGG4GCbEsgAc1nK7h2YRnqAp86xsV1grzozjbaRtOkwPL32pUX8AgXsPT
baajXwjDqw2zE65DbEBViudgfNU8Y+cwa22bUenD6ooaqv8ueyI8dc7SypUO/pND
EI9SO2XQhkh1ub7u9AhZyxBExKCW1PL+DeVgp30gTaR8gnU3+SWZy69TbbYuraVR
dscApAwHDHYSfjxcuHInohGYUzs0Y2D6BreUOyG+HvozqhNZxe8ORKmpOm6udZZD
UCnDHU0HvE4cQw5XFUU4rmArBYxLHHtS24EO2KyQLlaAVAOj0D2kUMx2ZD04QufB
1YfRxTivPApLPeCTC2SOgDNazMd6YYjhPLJrJbfkkLSUV542JeTjzkfmR6JTjh4n
56Iu7pPjliJI2hdXaxg1tpYBcCSG/vInEtn5JodwvLl6jByGI9gTWbq7Fu5tkwbm
3wUOmPo+26YXccS7+1rkQaVNiMEwHSfYB3voNV4n5tGaE7o/1uM4nvufoDrNsvtf
CUGC8isF24BX/E6Mh/lEvac+exVEhCtcNUp/YoR1QBHICOSnas4t+pbW9T4xH+VF
zfgSbEkmDey/yiIgtiUk1ghV5rQkq79R1FaS1nfACf4+1UedzIOr3ONIDuydD+oh
ECZUATpjWglVq2iLgDAbN863Cr8eQGqdiXlr0INq9F/vWUoZt5m2iGy5s81nscJq
2PoCtKLtvTckVy6F+fG2rzEyScd0OBYcdCSOibNMQGSFtL5JuxhBY2LDtSrc1ANl
uwgof1pNLovhGiDfdO3qr9REC8fG1Gb4RCEFNQ8mK6Lrfv8FDNk/lM8GnCJMKW++
UFJh53ciYqfB5OwDbfzrO9xR8af0tOoaA7H7Puia/FC99LwmV6lPGpzJssuP0sHz
j15bDCZLbtQMigqhrJy06qyUsclIpFJ/BKMxcdQMdgDkAAR3+a7SE9+JS1/pQqaH
OALX3VxOE+2ljVr2I0BTPUKh5vfmU1b4giDDR1NC89eMJKpFcCFMFAvGAIUPQXix
ATigl5lA9BnhNY3D45+FAqPpvDK5W+dZ5kwgPNmrDkfZXKGW2TvgjIMCrcg0X17/
DJI0VcDrrxUPRr4DtKP6+XuKkAVul6MisSPfd9wCtL6y13Ao0nCVPJv65TV8NZzc
c47cHjWa/xoRnSu0LpbC37rvpU0cjGWEEIqKFVXLuihNZon+SGKauEHjKQgmuHY/
vRBIv2k/NxoTSPNr0+fUqmJ/ZDMhtijID10apsG1Heh3CIzADXiLp/JakmcW/7OA
bz/yCuMZj50LJ9YKdFtkmE1jlZY6KHH476rIPiuiWli/iUhOCmHvJ5FFpaRlA2Yk
ViGISBT/nO7HllFp4Sy6PvmFD0X7pUzI73gJUJROPDPUS4rJHVnX8rFI6Al/xjbX
DJeaYEGM5RU3JfWtmUrQjU+KJ/GMI62KMGI9nOf9Y/sY0mkQALvZWsHeP0B/nddz
YQi3k6/MG7cDvI/tIrTrhkP0HIsyCqrv20dEkby6YlzSXLBhQhp5026+qTuIOSsN
F/83EFku1LL7ttA5GLJO+9n0pQAFjGAKkyAVhgxD5HOgkqMbPwd/NVbui2iqUN6K
270cJUHikQFg4VSvIbTBXyQ3/aR9oWrsdHdZYfub1OUsWmPqCfJMnwAPvaVryz6Q
P2pCiJRNm0Vh+uOCXpuBBGzGxGhJPKDikNcPwEsBsy4fDsr4zt0pG+JodSxQsByD
HtgrzLw0NQrUqMePgJnYIwXpYvZvECuJGyju/rjDDItLGerOulL92myL8ilURxTl
wILLgxQovqTSrEi4VLByUY0/TFOo7WGbKPX6XfmlDgxJ9ZMVXOBtN1BCkWT3MiQb
tsi/zAQdr+kIS+alJADTM8DHrDGQuAT8vP9bZG2GT2oQ4TUIOB7SH+FtDKHtk0+u
SRKBTPVb6IDo54qTbOyDix/nEXSw5lX2x3b2f9p+kKQVGpbHU4Wo4hkBjaeV672S
v5SrZWbS7LMQT4vKYqiPnUA4lInei/0GtLKc76IIMfXFEhMbG383zWb88MetRflp
4v/Pj+LH1VtIeeiJz8eQCzBW/JtO1HdZdgPSuNtf0WoWmnjCgsgfIAJFmhwEWEO7
+LQJq6VuoFqCEjw9wC1jNP3UOxhLfXcDdjIgEGX6/12sxQffI+A78hvOvL+YF5C8
p13+5Rw3R7Yqzl8n+rXEcwmpbUpNHyRBvui9PHcty2D7cl+rSZWGdMM5GiERbUXL
gX8lVEfNxWCxJ9uanKtYcNMantYMg1r/35+k5Rpi1Wap84ur0oLaVjzwZSrftLY1
gvg0fHGPK+lOxEi6pNBLMbRnFIqXHLWw4vsahCUo+Vf5pnhR4KSLuX/Tsv3x/3yr
GPnR7ep46MGIh8v8JVuoZStPEE0JWQWNHiWHI2YftXzPpnTchorqKCuy+POsLh6S
rR7Dng4AcmMPs01ArtE3+o5ZJDJvMiVn4mHJ6Wi3zRy7xA8Drikizab3LgGm1Zz/
bQotaGZWbRlPdFmMzyndcx2UEfg7R/Wuzg4N7eRmUzTumYe9yWgjpoK6NuhLVNOv
G0lqmVvSfd17HM94gE/BjX3gYTlS4Oae3KbrmtEXY95wBcNk6fe38QT0D8MBQYy6
EZ5i8t7c5zSKx5RzRzhZfULJAYZKQ2d+kc5AWk7xcXt8hRgncRG2WNehiox1El/X
qDR44ebmYF7ZSEyvVaPM272Vk51lBo3ib0WnWdPWmq+UcTQGr3te7Dy/xC7Cju1m
nLk+pjzJBnXJQioUh5BVaYaiI2KiwN6gqEaK9B8G47nKpVcrTv5EZ3MoVYR4ZOAB
SoV8FOlYnSOVaqLnVqNLtYfcYDwMv8WusPVnCJEaoLLfXTYuA80mvbpawJewyuVJ
CEnyV1yJMqgenrZ2am3BUlLcCFBAxd5LB1SfT6a4Bya0eFYCXcgg8iiDXWv+Ls5I
YClCBymK1LJAQ6WQ3GzVXjtNwV3JN3ol/RjrGfCUcZ8QMy2u1zMH1ufLcj2dBGGB
KfARH72S/npiOPkxxKxdYJz2KAR0M3cyEDKEvWj/hr4AYFL7jgcxgkkV2ZtOReIT
nNkg5S6MlVlIuqOr+ez+o+kiGK/s4Wtnj3p3G02mjePe8GhXIQ6xY7O9S5RXnb2D
/a8dz9Zbvj2LAr6obASUXxiAxNZ9DW5EDLVVItIuoeuqz+lw6CWXT2dxQPntxg21
55S5ZiTfX+X84EQMaxOuPVD3TWlLgvcBWWRmI7NeLgAHOdWPns71uWF2frZfRPI/
M+GoknXBr3CtkKHW6higPD7/oNQuYdd6L75FPB58bJBdi7iA8ji3tucuPeIueSPO
WjQdU6En5urJZWnnQahcckllbodepzAZSEdyQa/yYoLpEBDhuz3Rz86RKnzVmZmV
kFLQRXuVDFPfXyIz+MAwB73oN26UtaOXtWlyoWyG13jh37Z9II0HakTbouQaoFJa
uqe6r4pSps+p+V/UMZAuIRAC5aHFpjJBZpAHQQPcwdJalrEKingy0cwtKjpjAXR3
P6ffmn1ZGJjxTZQgn8/20A1Uut7rSJ1d/ovJ657zXBL5nQOwdk0p95c71tmN7CVz
qR1fZX1ZmNNsQcAzjt2ECEvVNMMkFDcK9KNBLcXNloG2yf6HCaFGw7QTXHGvCNPW
aB4MiIhs0+yd2D0S9LhdxGbKa3fSB4dtq8TPSiGNyoqNqr1gykpLeQ5vji43S5i+
2rAo/w+Yvzi6KppqRYAyU7ODnUFX1Pwa/hX8jOlsnDLPw7FLctbfcQx6fdNjfbK7
SIF3Vwv+ChSuBiWnfeJrgEq8/FBY+SwWZykH9Pm/hU3FgPKqJtgSS6u5gKenDVZV
/Ml7ysMg3bw0Nrt/x69P3n54iJBAmdvrs1cHrRFH3SBUrCj/2yep35+oR8tmRGT7
bt9iD8+rDf1HQJK2CEfMKNVVLfcvWPwGqwVciTnIixOcIEhTXLxgaw/6YIOO/wFU
xF49Yrw5DV7LSt9JjkVOF1yEHnNepljbVsjAMU/7fsJCYADfb5UnMg4uqhUjFzO3
uNbOzGlugTEmlGOdbFS224FALDH0en3regfmkFJbnqnVG93JDuh3OSs5O0fhAlXD
nBAbkjXlSCRZ8cZh8XR3S/SuwaJLk8lWYewWo5m7BF4ov+Z2iP+kLRk7jTcXXpBn
f/w1yiOmTYxJlVaCsVlEWHcR8rfapZeCziRPx+jyb66NUGtq3v3vXXK2PUHlaFth
v9FdP5IdE9t9l004HjcdNFgpFcniJNrjno+WFXvhyfqdQG0vlOzI+krlwJ5jfiO+
2z/hlCGQ6m8vSVMvk9JoaWwQxC75hF796pWv90bc5UYbkhHsmeAVXXBvoBvaHfMr
v1cP5mZNDglD3u+nk0F8TRC0IX0PXF8TEh9/FdjiQkt2PMEmlbEJpdWzm1hHpjlc
4zlljL0FpJuiWJA9ffOFC0YS21F/9XN81Y70A+yPNsSlwRpfOEDXzyL2tlyXk011
1mHl5F/spsolXhwF3B/wXVfkF5FD+HdeVKaxjWuSKdtScksxlo4whqe5S1DLJMkB
t0w8Lih0H0J4gaXgjBDR4LrcomS3bXTSbuT42zO82lg077J0iHndRpSFQ4537eQH
xCS+WtTnoxmoyWFPG/hJ7s5974tszyeHhGpChM1z+0PjM6NuMtQ0tO9MZnSqA4GX
uDxpO+C90tf662vKBrciglgomo2r/0qKiq28RAjPMgYIhGTeVFIaq6uxGGUVzInx
o08OaG/jblpvjSp/qT/g1UFjibjfTYIdX1ecteflkRozWLb3mZdx8Ggl0nn1eCt/
JTVz6l+LV2DqKaWLkGCAJETYfVD8XB47bTnmLo2DYYycm70THuxRapx2HEhSddmB
VOZfx7mePyj9ZJVSzh+Grc7IrFfR5eVmu/1m2yxI4wWg26XB9x4dlLFGZEE3OyBD
g8z6zyTQTOiSGkQpe6h5RmV2SOxqNMqvZN6HRbVDrQvPP/OF9aQl6lK0XU0CaJHz
4LJLBkQ0FTyWLvhEirnGpoKnAoN7av1BgfIcbOE93QNFVpJaIyn+o0eJR3YcmeAx
v3bGA0lbOm+iscjtqrfqyN3YO/Q+tJ8hspBA9BimlBRV6PIrYsejVsGihyoGarQB
91CDPGWl18zIcslMGzFCLZoDdS95iKF0rnOgpmNedbcC1i1wFRG0an99/dy7XURe
5Cs/D/As8e2XURkfa/lyIxB8Dn91i6YspqMpWdiyJ7devziwTTJuD82UV3aOzFZb
gypA+ObyY4w8jCx9u7iQcr0EaM9St2wZTqCC518Tase1y1O7CL4w0LRHH/d1WMkA
m9O9x38WBn7ziHAQasIJts4GeQsR3Aax9uQE9Qs866C/dINFj+MUM22ionUZI428
yWj3GkI6pVdWLfDSa1MDVt4MJUepMj0lPKG9CXVyt1WyliH7Ax1t8Z2CdQHpI1fu
ZT2qYL6BmITttsJ5T3DHt8Mkzxyoc7F3pXImI9BbgQsmyST1WKqF3zu+go4W57j+
ij9+Md0Y4PZHdMzFdznPdb0UItC2ry0+qZFUNlY8jy/5sVfnsmnZbeyj2wDL4idV
XbKmE+KIzzwjbe0Y3eZ/i3XQLmWFQBFmpbL/5aK/sQZVPjIUM8o79e7DEJWIErPu
7GAet8sXS1AqeVFgl6NahqQyDg2AW+yYNr1uzYDEA/C4+XpdQuE8YWJ+hd1Dqcdk
DX806xTuTBUB1hvK/gDAQa2SVi+7aa9v5ZPzNr6X7/WVDJnG9bMnwEHiP9O9JDe2
+dmQZOgeguZ/BQcOg1ow0o3pCx0AyDXjXprtkKhL2MoFPtqQ1rYrJ3PL4qf9BNMJ
bT+WOQQkgfXDhE21ljqEbKM0FeiBqdmpxAFiQuThqPW5AZBxwsIRBk4Lrg5oEKxT
UvLrLwRPijy0RWfYanEriR8OcsYEeKKDjW2upvO+2OP+SDj9u+QvQWZcIuTBr1Zm
1Zs5iOZSO4/dEtnEvb+W5b3wj+gUe4oUJ/ZZ2AGKlRivizCiVsNFqWV7/Keh64Dr
pk8BMJ6Cug2+W7xXS7zn9JyEaBAvC98hwaSByuA5REu69lBooIJVS8WoucEUlEv9
OUAl0G7mRJ+OOv4lBPFwG6jOPu/6/53qXSTN3tkyun2UBGP00eCcetIR8b3cg/wH
x87EpKEIIvCjZnVtsfDSXkMzYBI2FquM5SnJMgBYNiIQeXXvvy0r1tGjWN81d1Qn
DuhNx4Pf9hv8NVtaNaFw7frdNsUAR29rfChf1PZWHtzkY3g9qvt5B45hehePdcYi
g8GHbux/iZdeyS92O/vcCJ6akuUIxhQZVBCdkJzziXWXadU2Ajh7JDHfYFs2FhuW
btvqtXRo/IGZ4K4+h1uCUQICvZRlcYrtRzZmgPjf0u8aRqGTnf109Qxgq3l4F1Rc
NYYRPzBQoOZ2bGjTHPqMyaZ3iZ6qpTCpqm2sW/RTedRz3o7w5hx8SHhGSHhkhydd
j/+TrD3GJtqFmPTWTJ/h8lYuzUJGceVkucdClLTNPRnwLYugP6MwASrH9AassB2+
0Gxu9Si/xVK0YVnhcISxiNhujSApiYm6GQX1HYkZg8Ox4ekfhqLLFtwlwws7Sq4F
oyRxWiA8kYBmxegi9ini3Z2NOiQ8yy3+Vz+yCupmltpfvINAbXcoKWR15CrjhSQH
lwptQLzQBwKrl7J8VJzdeHjD38NNDwNHD2QjrdAdMC9reqlo+L8iLGT0bZ1rsXPx
3GTJsfvU8yG+fiqtdGZCSXKyJHRmW9c6uM9WiPsowSaL0eeJBg3cHNyWI9/Emp1Q
/JRd19uUPEkkuxroUdAaTFPmnVuQMhNSQKSkD2MhqP3tVu+azqpF2AShE05/5ZfX
ujvSzrqdeEIgheHzZD3mGw91UexhPVT0hu38xQuNxyYE1lwtkL0EOlugKoxsPTks
ar4WBK4Lb2d3L5Ba6aiVeHnmJyjfrEdG95udfKOb+KSXYLuylYbwuYJwmXiClrHm
0MstIAcXWBpID6lLwg3bfnij76kMbpar32Rdtg9jrWF1yU0rzD/8O349nYAY6LQS
1eigPYK3bIGRM04xAEwkWV48Bkf2Rd9gUkIM28bBm1TXxVIHtkXiKpNwqffqjyYX
SEWB8/uonTYvSpmzY+psLt4Z5XuKHo7+WYFMAmIDq1hVNfOd0P6/Z5C4Zr6uMmLl
88ulNQYeEZxehHlDla/OQHsLrLRJQQ3xa7FFvPznvkvsblLVn/6c9C9P4l3ChG6Y
Dc51QDKE2ecPpqpKTkIgj8L7MlVZmMNOKKaL8+gs63ZxHd1RkujRl76izPwlIQ6R
rmakwr2cr8u+5GdPxz5IWoWExmdWoJp5E90bx8Hx3P6x4RTdKq7tPLiTVY74pUCF
R8qVdi48D1OhWD86hDN8h4O1rmkLW7pVBNTCFXHOjoP2L1wq1DYFpttChW3aXjvv
19kqTCaFr/eROnYrYIhSBNQF5ytA4F9Bzl998RTcw/qqt29PTEmKMRFr1ptjhTQR
IYyrX392Ns7fj1yNvIhUq4iT5TNR6LKnSVQ0bNmQ9xnESvicIc6EOqvwFIlcV+qQ
C4QyOadPHyZuUcJ14AZB5QzI0k7J04iSv4NFeyf04QWiWjhUKH/TZOFhJ1z3ewXu
wF2wW6CnstNkWyk51GHPFde9unZHExBXIK2d81Ibk92vbV6p+7ip3PeH9D9DSrN4
oXu1i8rpQTTRUHPwdm5dYY1a6lUGktUFtvJzwmNpc155rGoAktKX94Ppk3BxuOo2
eZOBIlwXT82z4PehkWAy+77+UQHOCAIVNxAAuMiZcPurWEMq9+GeBMzj2oL3hZP2
DXfvc2xzfCGBtgqQU3ZeA3HU7oKD98fl36B/QUX4lk9mBNiJHl2uavXO+rjv0JrC
BvEW7TkJXrQ9h9T1iunoe1ZCD0JAu2yAWYsupxAQjtoHJuJu9pXVzbxeK8KlvnWm
ZJ48jza+xQQ7WpdkX8hzRi21joBM9noPegb7ZLtQ7A+qrrPeNzhb28TKWnqH9ZTU
X2xVsatNRk0nqhltqmtCk9ybZuKsYWKlLSERvbZ1QcyaYVW4fBbLPeu6zQ4DTMng
Xn1EtMAi+1jSWVtJFQDIf9eaJfIAsvDCkUrt0cNCm7oYb0UScRLQwnp5sevqgimo
2oANuBLb0u3Zi0+MJztoZBYh0DobSBYSNpS44XYt1ZY0fo6P50JXRL9kY5QsYdbn
JuEH806g18R7mgQEsOycowN1jBYm4PVwiDc1TRsGIs4maZoTky11DkHvBFKVz3W7
ns2qu6CUo8mQPOkpS48bmK2Xj/oBkNzVix0BrYevF7Fa/MuwPh60P8qH2vXhapSl
YVqt8t9owr04z21zC2kfrr14kOpqMbdXvwuby/9p/tVIMQAQ1IvtTFwhHLRcDGLB
UYw02KGGW2oPz527ipR//AQieUsmDXHklcCv6iksBF32TFD+LXwuoujKSFax1J55
R81uWX7JMM/rq1XUQoeD+t2zesUxNPwOUNKGCTFxBTG0oy4KxauKM0jq8GPVXiUR
P53lXY3Owg5NVO08yBQGdgmGr/9Kfcx6lm2FIgBUUXdp0y9iYwCNBPXPiQqYSq7x
lueIExyq9ZN8TLxG2VARBwi4frKfr5xkOxeCUa0cVJG1ql2KTxcQ91Ovv/PSvUav
g50JFk5kONrOzZaIOqQWXnYSqkSPrdJFJNFBGTC166PtMYb9lYcI6B2URDPm84bm
BdWGYRKXYF/KQjPWMFLXcHi2rXvn2+ab1ZM3ylonS3iUCh/LyDeyk+/3hCGFOqxK
2Cwme/pcZkOkzza6crPJHeQapD6+CNnr5r3bHlL99vm4bTeN2msxG4F9rGVeqw07
DKD4Pv2fZIkFh6TIbqjm+ZN7Kql6/3+om8cQxFPZP7eDdDhmSWesVrdkBGJUHiyU
kemcfr8xveE9TSAJ/4i3+LsQDv/1SQsimYuDL2vJxe6QO2SiP8rhTLQSkDLGAAUT
FsAouuIHq4nNdNUS26f0HUpC3Yw4z18waHkQmYrBVZPIuk9+EHiYKWfASPyx3TXQ
YDUftvZwiCOvj1A62NscVWgE3l+CT0kmxOWG6gyi4CozbRi+BmDD3IhA4QTZ8OvB
hkki+veVplm+CqctX/TwvRY0dAPXkOS8QSsrWG4xz6Of9kLZUg5AMhvledZKZDD1
Pqx7Ks1hvHwSPenRxF7+UxIyhjzaFoKKN0qAI2DAj5CbgPoehAgNodn7NoyhrVVk
Ido8s2LkqER3P8E/jtLNeGr9NQ/7d4rnpfaX4EE9nwCgj5izz4xZbdh3isI7Zo59
d1hY2nXhBc2532/1BosEenhULMGXpu91DOp8wuVZkXScWjOvBvkSnT3faBbTaYh9
xcm07WQjdkMu9wAke8PUYvkl4Xus6qQ88nnKF7r/HiiwHQg6BLomcdju2Lsqyv4F
1VWii9FP05t+xQ9KPPJHBWbhRfvZIGi2h8A+p33XZhPj+VJ5F6NAwStKKAr0ocMP
M8hWlkRr1UBxB9WBH2yNCn6n//dMpMPP+CchL3Wwtobo+cux3TbrDQQGnygXD1RT
MxImq7d7mlqkhaZbh3tVhtcF1mhEG1MIbVVXxWFA1iEIyoLJLkGfXZu4MgLZxjwe
OVBWE2RyqUHfIkeD2FpRksq5IPCiogRmxaMAZH3YnCU/cDkw5fLxWdwzzg/2Zns1
sSVfdQrmmPtFKq2cc0Iw5enjwvkILv5u2dBdJZZnqRhPLrqLED4/q/RTYEX5qFkq
ACtdT1zLLFV9HrAkhIZN+LYLz1XJbxy8lBI4XwlUbpP5I8ujhG7gz9cv3yRP6vHz
QDI4cVn/bVXAyKUobIRsnPFkFHIvsFhhDUXyPLBRo1UIjnx2xatpPsohOo7gCdYg
rrzAvIcwekBa00cc9yGHWayahlYAWNQ4XrBnMo4u7hqRF9m7QUK/Dw7Tu/qBJaX/
d+v45D7nCsp0wgkflv/ZjDXFCoPh5nf7dI+sfTGXsD28wosuzThI7mtL/l/egFoc
UMBOjrFudYJlLNZHFhbJE/u+eLy4smGmnWne+bF8geNOCxSgTcA18eQ+ahl2zPQP
kCl6Cqk1OeQE1W5y7ob39SoHoFXQd4utJDHw6HLI9PseT6EhNbclKkm2T78eRMn3
Vq1m0bQ1rrqm78fm9ukrdt02IzvSV/8RvzJaQUYE4tsjhxJLS/hu8GWwGG9drYKK
Q/sj6qbZeqbBniAR+hu1mHlJDbcT/zPCJ64IsyZTMVgY8ZPvU73XaXsg0FhVL4Gb
Iq1YCWZiuPeLrT/dxH6QSrBWld0ngcDf4940SuVnpc9Mg2Idj7QR5eogfA7/8pV2
6pJyxH0LrTuB+70cs9jIcGy8ba1sFVUfUbaDEv/aM6HovTW6yYg5oSreDmLxkWWu
1rCcRMO74iqFdx5f6WwjaFQq6OV0R2GLNRcxNoUk+A5pSVsQNH0eddrcDxrwQ3Gx
gSXc2xACjvL+04J2TyB6vevzmjUiHi0VCFiVS3+sjrDtWhN8AkeJyQiE8hYJEFGH
ZBqA2k74TqGfC9rs9JWssY+3crIRagC54SlD3ttOTUQwLvOsFY8FwXbHx2oQdtf6
560h/FyDm3cTnN2TcbKacbMV0ggY6l7t6NKRj2XXduBbWHs6nzlYosKHx2CIkY2N
qauz54BN801mnZBYkfVIqbvrJrzL5cAFIyjGyjKx68csma6DSEqU1a95t//NOsyD
1EP5dMpMbe5wUj/YlM+GaVGKcsmkPhdpxLOuroZt8n2e8cYutLTq9QlajsdXSTIU
+l7xva+kjklAr6LnjZSM8I5d1EkatGCFG0G7cHm6w0qyLDK9yA0cDb861bDpT6Rd
AGwk2HoZWYMpC0TJ87N4WfjsMnvQ0E4DRe9prZPGrQ42qtk2gpPJfmvPMl7X1mNg
7FyN5R/fERxjNZsjv0mjToFkmfRvQR0N1BvW2Lb0mPgq1L5uC5G1WH50XSy9Fek5
uSeQGiNBFbtCMFYH6VxqfU8CQmn5oDG2LUa4t7xXVQymdPcRwsQQOuY9C5OoYnZT
6xAA2G79ihmuP0F2PX1Qd3BwFk12v2dMnZ2ZKBkcy8Vg6r66Xls3UYv4zzfERgmJ
lX8SMNB7OZ2Unih+if0I4Rx6Dsrj7E2z/5BzqwtQPI6UZ0R6bQ6UatliW5csGOTN
Etcci5aRC1cTUESv0VC0vuHzYwsz2g+fBzr1/L7VFDZo97Ap87JT2EUzZ0XpPQ4L
RrKo/nOFv4CBitK4lIGA7+EXGaKk2talD3E9LkrprWbMe5W4NDou7ELDv0ay4qtA
oXh1+iZ2koJ4Ut7p7qV9pEiLNf5K6QM2wcu06hmhTDic1b4aXMJt2rkdWaSVCubD
wMO92R37JRkb/9mYLFvCbHuS/HXu4OGnvy0WquCcWVG7TYo29OPdWWo6SOd4b+SV
Jlhm2CTRXRPZCVh2INgCUXmngb1bRc/QX8m+aIM8wTTY0EDo8y3Pjhjy1r53S+em
SrktFP6RaGL8KbyAjUKiyEum8DTK77npNoKi1uUGVPNuiIezyWww9Cil+s4yP468
kizuW+YBqgu/qUftooC2k0yRNhUSe2oex7sVx56vbT9spfe5GsCpIt1ldQk/FA5C
flp/44/q54RgpFAJKUUzJsqOVLDrRtsVEHuzmsHbekvNm/XgUGDCKbqLFpncISq3
6nPagx3YKbunpdl34GdzKTCBlJiO1wkrGc4q8z9DjvsiIsAK58yVtsqYhvzhN2az
PLJrC16kStvtWJO+yL24OJKMC3gYXUTKHT3t4B7/HNBm6XQvhezhxP5m8ztjwYcD
2dt7Zu14gLyv8li0CUAuIaUY7mrpADvlHNktZcScIXh7x7SHWZHtrSafaI6H99Hq
MvE8JuesIXlEHmmBC6FA9xnP/TlXPp/dAAjqZWQSLZrlhqyI7WPdCS6Rkh2d712y
tF55R1mwTQwbUqNirzDi/9V7W7e6dB0pkHdp6r3M7c5cAOHMcuVVBRrgU1lMMakK
dCQqNDe4+uKaF3QTP6lj8H94xr1mBRoy4IsUAkgW6LBUvPvYiqfGkpiaxYDgo8c2
k2GC2pUHtTxiq6Lcz++NJvogWOM0JLlOnAk9ISTJ3zY2Aq0h+ziIU2+a2WSGMbyB
8NazCfcrufGqMW4b0XiQd+m88jAQGeZbOWs7ZjqYYYFUXe9icL2y3UOdUIIoaau1
6gkGk5FcKFq6+p2fg3f56b+iJ0YRfBfM5GT5Qufn+jncgc/8ABzzXrrtPwAjNHSB
ApQj/gePULsc31wLxwYCk8TiyISVh2udbH4O98jUFkBOgPLqpHzvlNHrKw+iYM+V
wSP9BBN3LhxvAyvBu3WfqZFuyVJA5peJ6qauBnpEWLphPKD6649h16nqVnwh96CV
8S6TV7ANoVSA+03CUvDCp2ewkABMLotf+eXWILS6Wwx8R/dqn8A0LOUtS7T8Qk5W
lKfvA26ILcVMIBHM/AgK12M5b3KUUUVfzLFJuXCJ0QeIzU5J53ajivD1Q6FU8teS
VQwh9LgGbjxURXml1GCb+1Q9mu5CSuGkkWQH7NVzNYUBHzUDuGZnSTFilFY3Zbo6
F+Ntkur60Vmedh/wSlXVMz2uZVefA+cUaVNgnA4uIueC5pfbU2mYzxwHRMatAikk
HZoLI0ybYEjWUH3P3VqPSWWiJPn1HW6SpqM47EN5Xs2YymlDht8xnRUHI6/HxhR5
hOg8NEB50oRWX3K7bhCOuP7rRY65p5H4fHYUEi84dBRFa+06PL5V7bQ6l/c78X6F
Oym0uCocTRQb04PMY1IraBpMiq3C0MXwPgDknLY6r6mjcK5tOqNeuJkx+DL5KTnn
+KBfcsZn5EXBUmPDmchWCbAk5T/HFYRHvQD25BAUq4HdZ0nfLE2qq6OOi8rpuNlH
QZyZ19y273V+IgOkGuCG84nxLd6UGcfrKCcljlHpt9RW0iA67w43BG3tqlZ031Va
6hnNgaegWvBzq6gof6g31Gq7+a6D8EZrMqPjOK7kxTOTpS2bRF0g9/hxLwzq/naV
Kq9N90MSDuP0ywYu7cW5XMmD1MssnxvlMDg2Kh0A0R65iL3MOYUm4jH7gpXpsf7Z
BzqYUNNU4JpjU0yFm8WjY5jDph7+lB83vaGu9mTCm05ipne3bjHQ94aeQYdUQImU
fPWqw87EVfGkNdFOh/shFBAm+hfu8A0njBEylmPUa7mLvoC8hIoJXd5flzAWreCd
9lTICWh9UfmpzN2ouKNoN/rX5nfs4d4dhUFzywkvPT5JgBi74BZtMWFDzS5sfLnq
joPeb5As6NVlW6FoQzWZ530nlGV979R/xwRcdUj6at7p69Mmc3llZDJ29nwSix9a
i3diQo88sxYNAyjLK2pH6XDLP65jFa+2MvAoCfFoyyfmwi6Qh5nhmplFMKTr4XsM
eu9ifMCK/mAvjlranXW2NaHKjTsQM/ayFi+K1EZE22nG5znNCadmb2FgpHjVLsSf
5CrrFs4w+ljE73yD3xnFbnqxIw+yFsa1q8d/SA360ed7vsfH5rWcrRjVRmwHq/SQ
n4Cu4BYEUkB336N/xVvwTNx0671gALksFqxUI/Oo02mrVObR7MH/uM6BVIYEoj1F
LJuZIkJgjy+eengrUfCY9a3fBXY1yYEEG/OUTvKrLiT7Fqbj504yNPXO6NFOTfB4
0XU5YsOUTpW3KdQGNYe6DbS3uQINL5H/v7XWWFAapF2BBVh/EtbYQwq8Lw6CDCzL
X7Z9BqhIpKD3VBfdT4ytG/etL6RkGlJ3LNHcKnIjXzPCF+CDRx6d3kY2/PoC/oTB
cO5BUhHtYdgQaGeRMC40IyjTz9PVjBPvu0FVn7Zxd9XD0loj+p/lwV+FQG77cjvL
vzlAFmjLF9kUpY8GrNJM+7Eq4TrCtC5Xz2ypRLxHTWrYmeHb/VavJ1for7Z7rqsM
6v/YJR2kr0TMcI8m18oo71ch/qae4ayajz2sKmzNePZQvmB42Qve9HUNyHfaRXhO
phvz1P08ThClLxfY/5C/YsZOTPruFPPwXr3Oy2GdF8TF36SaVCLoYPgMF5qpTDVk
ujJSYIXrPCaulertQcVni92B19E6t11oQAu3dS/kSY9/fs3ODUa7skOX+IubzeeY
/KuqQcxm76gmRYedzobHLjnOgpO13AjOb21TisUyN8ptgpuhFXY0dLZ+/Gc3vUPN
fQprdr/03uoIBM22TqPtv8Se6A+ZyvnRnaoKOINoHFXTlvXh3KvrnF4FZKGGrZqV
EBUhLwGaslet8nVi07rnqI3uv/GYlmpMH/SyysKWGrS2F4PmIwE2/mJy4+Z2FBH5
4aPHC7c5FgvK1APEKYM4T2zALUz7KSlG5SoKp7wf5BMMoXyaApAbnny3tt/rced0
eAJVu9VndYkkj4A0VTcn4VDxZWhqrZh54EMyH03ZUIdtxtwlfwJAxAciJaVNnf3n
aRApXg/ji5qpEul0NqZM1h4onSwVSu2SXCeBgT2KQYwtttkewZX2bC+yQVsTHw2v
+UqJq8K2FRhUDJpOX6V0n2Fd0SRVwntUSGKxU5mmBS6RPHote49NXFbbkV/il8hI
mLRYbAjbipSl2bkjnCk3Yop0LSbH7en9s98rdN6J53mCKx5r40H4Dzd17JLmwUm8
2OCom4zmzRMpRsRN5Lp4KDrNvM6roPijqIDn7ftOPydYuqns52dxS3/lFMkzb8aY
cRO8zHRqpwLvOLYTyTzRw5o8gve1DYbvwidtD0dMFy0d1hMR86VghJQ/aYHXxqly
BNfS6CRrL4HVQTkFH3V38owWOEY9Rl7WP/vvwxzdNJ339SQWVicn4OFXsd2MmW9e
fdw0wzSSM8HYE7W4cCXD0s9nkAt1zGrv3IaL1symAbq0yUssho6VNXkD8hx6cPpB
t/9FliNUW/IekjIh3rEmT8e9Rg3vGFn6UU31zwKtktL8jGP4qP0vTWvEAv/mLkvb
3qn237hi2GDRwF8nc/WVXXq11LPpFGoku31xYAmZ6J4yiQaw1+mbv3xOnna8azT7
RvhQO5qDo+AbJVl0j9VKgT0l9X6NBaPXEd3hC2JudLBl2atI+TL4FzPFsldh+sok
wv02/ZFfkMH0FoxD3q6oW7pi3bqssm6sBDv+zFzDQ0NlBeVtWgz8vYM5j/Jsei6/
ySikoR30fd/zFr1MGq4IgXgMn0v7jCj3/4mGKECgRHpC64kxg9YY4YVM2hQJlwbY
ZKTnDNEwZSYyAgyp7avzvR7DhjX1qktzRuBXrDQozgTFU/7w/2iYPF+fcpWn5shs
HLEv8PZ5fuEK1zUKjumMbSUJP+jO5iOmcMV1vW4d2/k64Bs5IwqaylQPy7Jce7FA
cICtcstUX+RQrxr6ZaB4JYvGIgZtoAmCQ+/XJZtxQJMbMhnDo0byzoBnegKYJDn6
sEUxOIvb4nuEpLilAv9BeFSWxfUUUL/eli9EAuHI8unpdwbs3IgO66pFv7TcXDaf
8yIquY/JN1nFhsFoTwYpVQr8iUSV+TOXSqHyzSIgg5sKg9t7VCzUUCEt/zxwyHhT
LbNFl/AlheHavzlgg3+NDjFWZuTC5Gpw9B7QCsZep5bbMFjmsw1aBgfUabXhoRQx
l1YkBANLs95oLdgcLmbr5YhSo9e9Su0e+Yu153btFkQGQ6NYFyaHbqwujP4PraE8
zPhAZukRji3/NxEX+7geGKnhWNGgFcde8cB4DhxKhmCWo79xoCiqtPiPX+SMrd1C
IYsMMHrg48hLI+5OAt5aSfj/RghncCht+8Eynsa3voanEXLelGK993oQVr1e2S0v
DnutIT99V5SticYnYXPRTZ8XkEJ99+cP9ydgjh5aWIztBDcyikqOy06CjNFkSTrN
bECm9SHMD+D2LZBvyNSwuCwfwcUAIjQlqIllJBQxs0qxls4feiaktBvV905kfy9k
76p1hBr7bnR+D4EoI8n0cyFrQHAxJWG3DH6Z7HDcQMPc4rR30BS+1ypEi9Ag3hAi
HhYcS1THujtNhPAga758htg7Pk88Kak3dorxFHLRBPcJO8XFWfTQgLHdBAd9+PnW
aDa8KhjiUSeJUWMPQSJOz28C35XvmUyPBEwIHF98k+/2FQUPq7jKUe/PCtfyc/2r
gniILU/0ZISVxsupPvQ2RqOdOpvPeSddKMAagKw/VuvsWfITOaClmfRQO1tM3oX0
i+PxucHW4vfkAlB7mqR1ZgmeZQeK4QKNimLfAywvQHtOrZZCXlPUi6WEZ0bKfstG
EWuHt2n15pYswGg+olQaP1Ce4QjG94OsGr6KGJ3/L7MaYmuNMkAh+d0Yf9A353pV
k9ypwBlj5AQpKXwai44GlyEbFHEFDuedarpUZjKwqZdySDWbFhMREMcOE7iL/Chg
OUJDoQdPBLLXWfqw5SCiFOFAMbDrqm0vQdxaU8VvkEPn8dP1KOoUrXyKK0p52JLb
pvmZbZ9UR2K5LSuVIfXLJHpnCAuIIlhPLzWl44x7lDz8QIeu0qZgc+6a5CTCJeF1
qqzA/6NcbL8yqEnUEgS1Rxq9JU3bfDDP3oFxbuPJgqzkVH4KEl/Py5W59Ojq7O/b
XNi5fMg8j0IMOd2neTv1FktedtdT5JpGWgMO3MWoXqRHF851FwyZ1yLUSTUq1ZBO
qZ2K+I+r0P+dVhZblN841vtD7NiprlUqQYpyLFlZmP6nHimtpFPNhGDEwGlA006a
eUgIM5JRmPS6XXvK8+ftsu0wVeQdW2c9QQ3CKeu75jhL8ZoJ5r2+4VOzqdGGlM4c
VxDtxBrIcDLJ2uy55gGfZBNuV3so1b1o440HOjbvjtqcVxcqoGAK/thKr54H9zBC
aQKgDbJupFeDLuBdNsXJAs47KHinC+jPr5fYoXgsuI7VYx9LAhJBczgTYWLlVOvO
C3TL2AEz7wbv3lUemuQIXSwslCus9K4RdzI9H7bhrJmzj+OL3kkADI7WH2Wcihi8
tvZEcgvGpXEg0eNE8PdzMnY5c67iL5f6mveB1SE9Jirid/KPPHWkc3NyrpFuOvYg
L6Uv6NFuJXsWJRTUN0x5zl6v5E2qt6nfUq9L2AGongiUja3/luNwo4sA6YrHwSUT
ZNFYSLsNz7cYXUypxfs7Zsin9/hF4PWMfEhMscDWxbhc0SnWH9sY7axfsStUqS+z
XGf3YZfWBnPfrg5YyGyyCUt7LrFQjGGwz4Av9unhqVo9wPbBIWzevYQlM3zvj0jz
GcQsq1GAIy5xN4Q1NnkAr/dzJ9Uk9fdwpSIvIUqGNPBhfM7VowC4I/FdfUVUhuK1
bhRZWvHbimMvyOMwA44fy00hnjuPYzivh0kiapZnwYnIbtkR4MXatSxVaZVcuaJ2
/k08cFUcqsVmsLf1cDPvMxNHz1GMWLIZM/sCURlwvrz40k53av8vWRcrzLUxMnOe
MN66ngec25S+WXGte2l0hX1lT6K2fHKJuCL4Tg/DBRmVhTMgzoqW/x4fTIzb81SL
Q7l+rJ8aOQRVMp4zfjRT9KYIlWe2bbCXwFWszqDS5F7dJ1sCjMjM4FL7q6HHWaRi
IaFNTZSxeZsFQifJIyc4j9kZt7rBANw5gc454rIQbYDZiHSoWh9FBv+h92XakHiO
IoHT8Q8aAXHC47b+kbA3erSDPleDI7ShR5dSjMZiS6UVubTJaA31FuinQ8Mhy4Xr
u2zOqpl9t7Bu3UNmH0ikMxvKkgg73E2FjVCM7+AsfcEJmJQlpVBLz7gAgYm9wO2u
TNXgLQq9QN6Q0oUf0enHJ1tjXP6HCyYnkHG8RxeBdxX7DFurwCBNAE0sayoO4tRz
tiTIqil01Sb6VP9wv+aMtdGIJ0zC2fLCIx+Mx8RxmXuVMhGntsbnHv1W/wLUtzQG
Hledl0tSthdHRis8XowkKK4YMc09eYk7QtK0u71BYf04CenxAYa1B+P2Je+5ZpFQ
pYdWkTDOPzWEeYiKOQ/XrbwuF3PJJIs7cbtPmLyCQuV2v/BojHVau59rCHNOnbAI
1WJkTjt+7HyheNxfHinahwY588qBqqQhprKwCJQ+fEFI869x07H8Xn8E0uJzpbzs
nV5Jc+1EiRkHsJxg6zWwpiazgy7Wcgyi7VSOgdFgImffxfovKf+JLX9LZFVRhin7
gi46xUWSFP6Ki2O7vm6XsFHHZQCl8dle9HMkPP4f6eYirRSznUnCqvRVmkoSIgaV
mK02IjH6C+FDMjhb3eeKO/nt4Mb1kYuAFqOM7x5Oib63htVtfpsxZDcCMS0yo+fy
qnL1vuz5HVx6j31CGxpqlB+Iph7bvNzZr0WjZ5FID3/v0a8//Ge77f2GlOWkJtku
9+zO8KLctyPT9CSkAQnkqIc7u4trQEyCAYtUrgn4376qoDfZcZJn1di8UTXTrRun
1RtOps/NQ8UselGxLc4hCb90rT49oA/+GOfpCeMTOhU0Ydpfo8dJ9qZPFXLP47/D
mQhtM3N3tPvY0Ck1d+3GcdPvQPD1uS77gClTXPGmZdF/OCvciryL/NabCoTeGxtT
OOvIAyN0Ku1Y0FQAOkPcWdLv/cfPc4xtUfBURZF+1sORDqpW2aqMeywqUH++o/B9
2J7zQnGqMtotx9vOyFeWhyhMl6YnqO2aPVCcSZBGmc1z/aYbJZz+EukKzknjPulN
YOMwetH4c7WdMuwIfOAFecKQQg+ETH+jiyZkodDVq0ikS8/5uq2DVBxVf6bIswyl
SqT+ourtWFJfcAK0iZPYEfvT7ZtqeDvxu2Kabo91RuzQZpIz2ocMEg4QJdN6lnAz
v87tKxjv4X5cvXP/PvnnqbEAVaCeIrJjHmrfpELsEQ0NWE5HlG5Cfl74EdSclh8J
Uf87NGpiHq/99/ZFgyb3W1MEk1Qpik3OlEoJrZmpY9915xvNL/bol0nRiBIArEXh
q9o/eelTIObwAUfgsy5B6a9KE7viC9OLZYurEdrLqI58PE1SyYDK+ka4p8lbud9a
8cnbbaoTebM81yHt6STF8/A2vKDjkXAjVIP12j98WygkR3nyau4mGyx589lML757
lNFFF9Cw01LbRKE9wa46DzfsFekyz3XKNzdprZRUX+qvw/6myaCYCOwwLyTg3WOs
2JMEoG53VWR/rLorWIEHCUt+bzxyy2q6Bb4cxz7eV/C2Fqecp1i7HR2Mu+iXX6xz
UgWyRhIL4NvwkvdpALePPafUJdHSG0DKAcE4wgmdXTDVBj8nSGA7iAziqJjrxY5l
ttZXAnByepZsJMz5XFZDCidEeJDVY/oRQA1Z8fJXpy+u8MNPQ3voyUl3a9mRWe4e
3FAHspqMzfsXtIQLufoaHYnyRIvDqyHAf2NFV0L6DHqysD3YM8cyDsiEAHcX9M48
Lr+Bzn3BKlY2eqjfCWZjwVbGhLTJ53pLR42AOVc1f7FJM/O1UTb3EIBW6thD6BBX
0Pk5+iihCGSqf2vnQFL4QdgeP620MPttPoqkasRkG3G2/pIIEePB6eT6fT9xK/go
ArBRnEYccBpT6IACCc/eHwLH0OIgYy2G+qk0mta4At8Bu404WPXSewCkmMtrnba8
Hgm6Ky4W+CBnkivWG7Pt5CVhc200PoeRKW9SD6GbKsYOTYb/jGmFPIxhuGPVixZ3
z7eRrg6+HQ89yWqbNyt9Tjbepw3mHHmbM5ARubOxCputOl0+AS1XTnakX8mxdGur
LOizdIQCXHSWQiTIHYwGKvg4jZp3p6uuK7znltZRQ4E4MQ+92XzNsKZ2TmZEN+Mt
l9EInHccq9ywMclUS14gspcBc2dovFgldA49iKMBzSR1lQYr2LVC0mjgkDqCuzH9
x8ADePKQi+1jdYuZelGUCjdExNF1NYcR4nFVEn3Vh+wo5eY5VOWvQR90EDg6jV81
qJ/84O7lLLxSNerKnSvLM13vLXmetof8eCS+YrgCYXdHj5X0lrlroOFCngV44v1+
fJTMERzDBr7gtAdTn0+4bREZsLlwIpCBEX0NqIqKx8xtthiCbu2P4dH8A0YdlA6c
DmokjoFJMxSDQ7LXgFI7m69qHFO7blW/bw7XpsP6NaV6p34wnSYlMLsqQbHgocma
IJOqQb5c8Xice7iCTbWHNq0oRKtbNdhBzGjBsB6ouNmrItvct4AUwg8aNR/0BZrR
IN1prSWW8k59lAvID10Ck4xzeoeiW1XxRN4WGb9KYiyB8kXjWmw9i0XnyA3zBFpP
9P7EURTjKlk5zrcNGoaStm8ZQYjrM+Tull7OBX+9jVrdA8rLcCDvtmFONFyWwsUr
eO2phldeGUb8dprYX/GLfbVKD+Nlen17Q3ikgnXoenmFAJVdNAk/xittxjaLB5BM
DV8iPeKKSf0yANwHBz7sho6bp3zUf6Bm2a12N4cV36nflvMeKKJyZZEPGvAKg3+b
1Al9K6VLMz0EqwOTSaN/pS9iszIqWVPOn/ZTuY+g7q7Jvw/LpHXz7xk8IniqBamI
YZAPXxc9hAl42p6Rsydi22bMxbXikNMnVBVJyCmRZqgTZSq+5lNlYbFr+Z+U9Plf
30Oc3OZDB/tXkGmQ2C4U6pT7tzfbxkmyMJrDI5tqy73DB3+cLvQyIxi/lHYVRFyC
WTH87nCkIAflgPNQrn5aLY6YN0md1KYAb0mXFeSv16FO99JeOxNQq/hKicrARBqM
uC7t0k6LEIDiat1fhBCV4Dd3F9xmFXi4l+3JMkanSxa/yum73F2caiOz2Z2zZ13D
yrJu7L33Tnq5zF1OxNFAv6pqsF3RdiAUP4cj+IsV7s7C1LgVKLZC228gbB1xkwKg
qhUU5vFKvWkuLG9xm0ZE4ZXjU9RSrbCnnkiM1i7MZteM666UX20isEzpBi78Cql2
iMHYfq78UQmgCvkpklPIN7w08zQiCJaaFiqciCh6sso75XFqwMRz1VNgB2H/eC8k
jYGLGUQPGDHMuIm5v7jg5/YEYlecQC22SB6sJB9Les/UZMJpdcVbaixi0fGExpat
aGM9FIU0pz/hTZssFw0UlHiCmf2MGxSebyfWhjgWUuLOzdmjf1wen1P5ga7eU4p+
NlGsUL6L6S+U14rhocVlgz6ZuUDPxONaspfdS5z9mWZWdgDLl41E+8s5aBbT14f7
AqwinuYeNvpN0PAkM8fZ3N8nSqznUG8RVTxpJNy2MF6ALUDX/hlmMSKA/uP6i8pY
AXBntFQq/NvLa9WvguoOUECHw02bUHzBdcUAXfkd31e4EpCBWJr4F4iVL9Ff6b1k
j85vdm8AJpvi34Jd1JdvwnLwPaK3zwFVsJvMSQMPhmovHPHpITmRDCD6jRnml+II
04ThtqKDPRlN4gg5k/sIF4fOzFrBhcBPVBKkXATB61D157oAT65ihXTJE6WnVUcr
CQ0UsVdCLGn363rbYS3S8Lhn3K5oj/4D/2IqeMg9mdKUZ0sAba5lLvc58uzqW5zz
f6sHf4Y+EGUzedepUKBvdQduw+9vyxHlo4icLXPlNenwheOf6zxztjv50m75Hatw
4MPlpZgy79XYgKrPKUIVjcoweFia2IvMRjqLknU7+0F9WgWSq+b0XvykQ/KVlQ+z
zfW4IpK8qdN7JwbJ6PHlZOUEKSm33pxfUJwMUf1/EE6fJc9/lotfwznTzaQspwDb
Uds5Dw/k+zEJjQlTeZ01qPM4UmMzo2FkkAM3K/IhhiIcfaXbhq2tpWEpOM0KpTxY
bHCsaooM60HpzdWyjEANAKtxJkrA69qVK7mHjdPPpV9szPH3U3TkLoZ4V9LvK34q
6ycor7UlN1qnJg/buqwDOGhYq7/JcQBKvVVTLGNQY4qTaHH40gyuHHd+za5P077e
nGy5cQu73ai4bxALaWFTg4+7ijngDxKVNzvEW6K275G/RUkR7kgQEwvVVRJnaQNm
RUQqv6ugCoGkwjpauTZEEHb6YsZpV3NHwLDSL2GUwQprSQiUUXsehCfv4+2/0pS8
V5/75TtM0jK9P5R1x2/uyHkrcoS8YXS4NgsCBy5X96s8H3iAnFylwkAW3Add3O+Z
P6v7z8hm9aiebFoC/Khg7/SSXwBsFRQw+WPsiSaPh3Iv1oJLyHX0MUI+RAJV8gC3
EygZolqj+4ZuQc0yZSkGPgBYQyisrUOv9W++tWBdufWBDHrEl2bzA0/Ca5l8OV/3
3ofTfgDUXqhskPxdU+VGpDO0JvumEvJU9igQqw7vMUIsdVvVQ2yZRwQzWUzfb0B2
IUK+atNSjo4UrhKZXLBCTJy6CQetnXgBlvOFTaJvUufgpr7FeW9m7zxQFenuEJ45
7AoIEI0F6p7K50sJJD7HIq6m8GdLfvbidHaNjBJ1wfmT/37lfuqLvq+tEYLOuDO/
jcqgU9TiNbVy9eZvUyGXpJn1MWt3dwj2DuRbJePUbmU73F0RroJxMG9w+wUq/R2o
rHiUjSQ9EQM3wAlWzcvfodtcODxef8v8G4u9LhRgER3WniGOGQv0hus2Vbna/xfR
5jsJWISu4KxXyPvjiRF60yl3AGupqusPzGLn5EjWLxfl3G1MPI3NZ5oebytQ5R6H
ttmmej/SaPS6AG4g9DQg5IGa8/sZmf4moSr/B91A6oDUT1N8GYUJ/dcF69KwTd2M
4YqMfR/fpUSVqvlMlX7GKpiYkbhF1iwKnlaMev3LzhPitndzB7kRCd9hezFU4965
J1CR//Ts/ylb6GBeq8XnVfQH6eoFjoalW/A09q582iF/73GvTNMl2YvwbwGFm41E
6weMUUo8mrT354uTCT+9C/Y6uIbW4oDt85+E9J4reJvW75lSe36sKfp8fZeKUfIS
YJLw9rWx9e1NY+gjLX79mIg/PP+FlbehXQNxd1M5xm3bDFjc2FSydJpqT7tRSOtT
QgnRcPAUG/rIBGJ2h5IYN5ugjjAhQZmxWFboI1FC6TK9DH/1cRFeeRM94qqmbnql
AaHWMPwQoscszDDoqrud4o0YBBVnoKWRwtROPx2pt9sW4zC9W9n2NIvMBOZU+a3y
24LIXvldKjZm8kTmLAbUbD6HAB0Yj/atcU09ajc9rVV0rXLtvRNCJIjL/7x+FVP0
dSSrSIJGywSBjC0LHlu7haOTM/JHMqDxSyqHDGKoG48K+UvOBlykhiGyPkIFaq8n
x20AH8/wGhRcqqqANHQ6hBtkF50Msk7Kmd/FNL6NlyIGT8Jy9s3BomeAwyfX5fYi
s0TKiuQP3hVw/IGt8khtgXuoORiNxmE1IWxfahUWJF5yT0kCa7VKL6jSpZHEiQOl
UBKihX0wfD1jqffpnYoe8DNdElKCG8qwOm6xMy8tm/hRhMCPEfTLA4u9D8ZB3yFF
1GLAjB3xguKI2ogkjsXA1DimrItMc1gEFcRCu5NJlmnrB/XhKpz61oeMoj64wUw4
W5ZByutlz71Wvv+KlwzcCGeSwzw7XS4yexhvFEOaNowl+two1DBXPx8clcltGOmb
EwwtZBBDyaVk58kZy2MVbsVmg//nt7gl7gVFEsOlX6Dvlerbfqv7PXoud8fVkVRS
2JZscNGPgVtIv6d2kSRpW0KAjn2xCKHlMVKvTeJSRUGkucqJYlW/+8GDfq8OSw32
dcotpmbE18b8Y9NT9HGXA06yoIjfd85ptJbs18HQqBODgAt449laGpFeMf27ySct
BE8is4e/51XxXteUeTUIlzqOy/sZH/PYOJjp/7NU94xuQfWmtfPuUBgDlaTXyYl/
6GaCD5ZR1wI5jWZoBRpQIRNLk5dQi3IwSMEc4WKdCiBYx3SCmrD1K8lEKkqVOOZ8
wF7YzEPztV5v5C/qPiA9TgeRAVgd5GvV3M7/hBrGTPs4eRSTC5htkhNLeFnkpiV7
99IEZsEOIu1MsD3NSZQiXV+vFQNNcGxAir4TU8POLI280eA66L/2XYu3AvUivAEk
3AAwcX53jPe7zA6tNNxSQmgGoK7EoDLJPWKZ+WciGrSKDJRH85/mrMr8zQY9uVgd
Zv02/T9IJl97w2sicXRT+lPjD7KtNXwEXEMTGBmhVPZxs6gQfOcNV4Bfj9ryUU4N
O4bXpcrYosrqXF9273AHNV5AdAajvxU3tlaOhdA29rvLd/BNr6x2DL1Pzp5eanzh
yaA0gVqV4z8nueDbxaUHuNNUGK3dnIVXz6EsrJW6427RlpwxwQgUhZidNTi5/Tom
2ye+g8T8sVWDsoOG9I80I82PqcxEa29UPQlEu+oz7D0gHYzBk8c4iHMl4D7CFC33
uE+B/K02vLYh7C6s3IjEf28dohKeD/MSzcVM3NGKcVJXfusTyCNM6le8NhI3OL2Y
uUJahN7WUFQi1xcikytw2QijFXItqSe6KcuuVB8hh/n5AOrq4jp4ogz2xqwvh7tO
CVx7Ym+SiCZ0ge1f5zwp31evpTPYk7qZ2MS4yB+JzgOBKJdkD77pmWeU9WY1R0P/
3yB07o1q5vyE9mX7/Iaghxr65YExL6OY6SEt5Xk3h3ZeuPqBzR4uXX7Mme5gbrcS
+OAQH8YC8jj4ngzue6gtb1Gy9A8GWL6k7tgHYcadCIF5ACNzAdfxi8Doq/DHZCOP
QYwh6dMD8yF/4EjRS1ndTE5UeQ6e6qmhH1kgZWkai7Gz8YaZ3IjH0nh6XDfSGUFd
K/GgyIA4jQPhpUqNJtRgtcqIsTYhGDKlzVdLc9juBCfnqrliwoXnCN2FQiOgnCl8
PwEytzMoYqfec3yeVl8G2s+nju8DV47V4CH4rcUaX/nDFPitPPg/uBMq58ahTRhy
KycLwzV1zwy6qaQodpOC5dzT9R5iYT3BnyLHX4a7k/USYYLTOdSj4XONgWUAABXf
df5J5Q+JnoEYxtu6vGWDiOHd3h6KSWjSB/YIKp1fBuOi8duH5CBk0GNZnecpVgYK
ISfR1A8a3CczqmwABx3rHUtJpvLIdR2IJJ5UnIGBrpyeTt5zt59vs6TY/t0XPi6U
c5XeFUkscU0pDLKbJojJCymE30jjZqLQm08blCr1dV1I8bnQyTx47zQxdTw9K+5D
ps8/OwWH/Li8TVcdgaArpfbl69hw1y14FOGofKesgn5t3HMm1rbvPI1dLR/xX+o7
CXIHEl2qQQkmkiwcpq5BKlaXQ+/BzNfwNn37ciPUy0Cw/A/PLYRMR80D1Tp/KMEC
LiIArdXa5ItTaJ4pbgTJ90w+AFdRHIqB3+0czy3c38QI0pHauAH9XmYAu2pGpdJY
rpR1V+11evr5SG0HfPNYsevT24N8HQAIHrkHM9o17OadWaM6Iqj5+GpRIvexVM3o
3L8QniUpaO/KmYYhyTld78Tt251bqHmctQswO5yCpwXCvqudcnDIV9jwMyIgK1f6
SwtESFs/sSSYmoUWtQ8fSIbGzQiZCZPZKi0xbmhxri0cKadZD3erQ8wN5s2/rVtA
CWsIW9NaojL4sN2tc564Tpsj/LPWYU2v/E3fCF0LdkUD+irFGzIZesdsFDSt3RM5
dbFho5bChFRGsalWzXQWlJWe3QG2pckzR6gNe5klB1VdHHAaq2V2JswstF+Rd4MT
0uE7Wt+I3N/CpkJsDo49Vbs8aFFWBSS/Tzq0hBcU4V8m1DcgXVj0bGDAFN2xQKbr
2eVMT4IE4338cTPuXkWF0COhcIQ9XtmBQ9NmBnhwRoPWAE1xK6ylDfkrF8fQYP5C
9r/a1/whflZq2C9nJfnCXk5EscRKxzILxW9LE1tlXA5iCyEXKmOhJudNWKmysyqN
NOuaocuO0xuuti2vqLcc8diwif0B/+AFEPnUfgka+U5SBC1JhsDJg+i90fOgVFH8
KH8SwSu23lyrxjD9fUD66Kfhe1y1gbw14mDjBIbeWM36LveavEvDT/cVbOzC4G4D
AGrCIhiPsZ+2ibCOAHPpxwkzJXB46iW4N+FruR/laN3xdJA5wN8JY33XGMBPH7Jx
coCP3bxdglmqtYgSI3Dw8TbkSPbaewkfbeklc8cNoj0c/y4wzg/Ha6jOMVjEUdYb
kzFEu7atjzH0ZluGmjB0BWlS5CVNZplkpEpKqWYiOXjv3SmeKxQa0NwHioGaKXbJ
vsQYooUYo6/vYEN733ExIki3EE4mQ9s6t1nY2fX4ELKRfGiogwp0q4l9fyuxxMcB
p56MhbNXxK7Fctk+sKVvaVJBCMFEzzT2zROAbnFIuRAPAesiT8N77dWAuBUTjr+D
9j7IK4m54kDJPkgzAwkaM5i+MhPAceRZmN64xs4t3OYY10ZLUwhEUeGUz9pBg9h7
wc6rk/VFueV9M1cRBDAWtUoHAKD8a5kvMTsnjlxjmTsSO+ZeJGb6nODnDbGmmHG7
HHFevwJtHZOLGJL/6kSeON0YN6fx7QXfWNcKyu1BJE1dNdocKI97J7IHXQATi+74
Wk4iTdYtzY1VxXCQy6qLQAoPwVnYgE8S5u9uLzAwtHG38dEAzjoFlRzF8a157o9F
/HyRhwD8i4dyAHdNhgBnGQD4zcHV4RWpxjIU16uHcvt5naMyAhojDYKJbiN0by4d
XQx6E2pXSptsP+yRDHrsl47hq+Jy74QP9+7O5RomayCpC2qraJWpJu04kh6Jqi99
H1KbyK6YWuwnoiYeO2wF/XrUrqbFOY8c2pT9NaOunhdD58hF7uugCmOn09KFavJC
lbcumiNBm/56WSiVWsrJQ6F6oNkjZygahr67vKOpzle4BYu1aB3+Y2n3TVtk4N0S
jIucdiPTN7YGJK7M/xGLoHJVPsrPcWV8a75Bz3DWuX+8EMMafGERA4Iq5McnkDZm
/+V0VLCrFLoQi6eCO5nyc+wl9QKo/NUmePSJWg5uauTNCepeHiRXlOcJn1YHIdyA
Vw6UWgSTML14SGsq6qM9dmQVnHyBXOu4MYAZ1NVY23oqdEopGDqbmY4S0YuChHcT
lvKxmP+nRskcp9xjwYj6WNtklVzcbTuda0cu3qhXi53bDdrQgyZ5qYzyTk40IQgM
PQf1ewd23ZB+X+hSoxVpD71daq9o29XnGS63yqdQ3cGx2oTLgn55HpgHQdcwMcwL
7uW2uht9acZkkOjtJgi3n9T7vTeB6KpJnXf+O0B3CLw/k9AD9oER4YsuTF7nZyr5
ai8IXnZHY9SlHXObQlU6eVv8eF6Tc1KjTn8yXJ9Rkdej5JewGts4b4JH4witJh33
ZRT8Pz96vuXzzihIQ85Z+hUt3niDn8/OoZX6mftBqittUTOzhsk87N4vzE5C8Rv+
fNI6Ze04gHMvA6PfmfhF+Jw+ER+zTcUOWL+3GWs7zCaxbJbBnWZ5dRY6P0oi7/EY
Qdk4tKY5PrAKSarehS4SiwC5wEXnqdSFWmJhiY6iN4ZzOjnsYuKFl/YxtjBMkawI
ZxD7XGRj3q2Wipioi4UxY6Ilvd4+EQinpsR4LeQzxvYRGn4s3NSim1OneSnKWmbj
6X8r0BiBhdIu72uC2jwjTCpbZrQX3uK/oKvq16cM6Wu6kQ78tC6oUoOzjZh1Ox5s
cTJ1Bkv11efl3PMjkVhDR5KJPh2m/0+RlwpGP9MxNT/oVq22Hrq1ch2IZa9HLPka
RBF+3kEhRdpCe/kxedUffWvVVp3ZvnWATZzQHmVRgeeaOfJDhu81MYjLALJOHbFE
Rr3YBaRZIFMEdRxWKuumALBnpgVS+4LQx7NILTCKFYUAsGqA1TxDqw6gxu8ev7Ax
IHticyFC3sbrsUpanzO3gZsgYZ7OX5fyPJ/IaLEDsFrWxRfA9w4mp9TbtY356km5
o+jgLB8QEBd9U+4dcMqncTmEhfWGT/Ck+UpdQHobw/tF2BYvY4Lqi3gEnVl0XZly
jSYIuiQ7F9ajV3SpB60uoxN12zwUDdqgqGMGJgsHi0PRcl4Gnk6ANux3ghRfdPK5
8WcmwIide0aw1UyJ7/9jWTf0QmH+ZxP2be9kK+CTT9L3s0cHy0sDlYPJ3kEGCd3J
oZoD6AJWl771qCNLewQrJ9bigcR6dvERTBwqP4AvliVrAKQFh/8mvlbyslB1jCf8
ryymazQgbbFmOgVZK0+patX7ObMUkaTy8R7xx6lJs8ThT2GrzllBIbZEME5MsxtL
zds4iy1+G8VAiJo41PMaZTls8Wt38F66BUlhIu/KVffyzJcNNV5pvAdthMj6PRDR
ojMzCrIairkHSngo4eMdUD4XouVZnv0106zxD+JgYX26A5Vm8aJ6kAzWgccXUvEA
7zBkepQpBbSoE308RqCrqeBNaEHlvM+d0e7CZsXbUoJoTGxYRUMLEIpUMO6e8mEB
zLEeIeHrEstKd5cfC/wACchyJEmqBZqXQlhpkzSLa5Af+58als6TxTipXfcSDLvR
gVTDptOKXNro97pFE5mKvXIXJ46Ex/7AXo0JwTQHSIT3e6acNcfX0IEgIRfJdn96
mXuwLOTefGW9Z/ZSVGUfCnbGmUgf2h+GT0RmoQXd0weBUncdo0gUm8UYZyT1RTkq
8o2uvLzY+bKwhFRFu9uddEXQFrOIlHEgQNSKcPZIS0Csy4cRgVi53+7pYekt7OCy
o5KgYLVxefJPM6+9K40mDmKrO/GbROmqNUosaB4zo4+JLKF6WQxS+LyElePvw25J
m4PNPDGD8sW1qWWZe+W27kn7hbFyOEoF9Nyl0ALhpljNez9qnlABh7V4zXmmDRfw
geC+fdXIQNyX5sGmb1Ty/VcCa7GnV35pmVbZ9gskNLk722y6vNcOKtVafICFGYcL
Hq+JKcNY4mmUt7eil9Sf5Jkb1efXpmHDs6/Aqgvbq23aOmT7Rbd2mCkeahsoJPZx
sysPmWqrhXRV/qXKnh6ahoheSsHx3ZypmpBLN7BrfGOlJW+YqWvRR/PXIZENzPFT
STw8M5d7hcQxr591swYRgYlKkKZd9CWYqbzz4Sd2wb0zPGOaUcR8xzaPzo3AUhJI
7IzSbfZQ6JsA4foe9mHKbJBcG+sEYEjSKWDhZOIurm3amhZm+YtxKr94l2x2jPHT
yjYmCnvnn4lgEF6l8002diMIJQV2Jsc1qZhbJZ9os//f7LeYU451l+gcTO3i6b/s
sBh4LZS450SCu8KgHoPrY/wWVSuRdypJcUAJozX4BR7u2tvcZq68K2w4Y8TXJ8KL
vhuztSYufQhudWq2oUHRMsAOVQ92z0wG9L69po74ZkG4NJTOBMPAFnUDVzsMfzpv
QiQOOToqmByaYba1+DXTIc6vDa0awg1TxxE46jeIFe3ZzB0RhGx61rQqWjE4/ZFd
SBoczBHw/enl8LKyJsdSwdov4cmeZ59qyaxN5XFRRiz07Ta1v0f2aOftxSpcRm+4
b/4pT6tnSywPxFYbTFHmaYA7l6wUv6tHCm2UFAiCE5j99RiWhj/dEAfSIUic/Pop
oDkHEWqLwYS4pxTGvEBVHWQfpOQCDz8aj0uA3BFm0/00zA7AxiqkfCy+Clch7WDp
1BdBf0jmGpU2KocRFwNI666U/sbMEUafn4kzHAC4/4zjPyNQA0Kqg3NhDGOnQAGq
7nh6+iReY0fw5kyjSgzNuy08FDI3OFJmqA0xFeI6nG4sNNiu15s5FI3pXvpsM107
1bq4GK44WD3vv7F3397Dspio4z3IqHh0MRm6jh2M2mnplR+2dWEgEXyGjY4uY2nK
xeukubha4qSdnuCDNINrFJxsQabV3sK1y4FpSY7kyOXywsRkPGrumjU5WVsF6dkl
rfOEd0ngAPBWtQLxzCr718hV/UkYDBprq0ZJPcUdpM1lMuminAYH/agtyw+WLM+a
wKj+AQFPsRXRjL5ALll04aD2GyjkySvFBREYetw06ZiJnLm2yYsBgZ5+e9fbNRMl
D/0GxVjURbxivnmTs4mmTYxPCXbWvNXG5Ka3+DJDE6q3YBHnXVG1qXBdFL4gjvlV
kjEieBXIjyYQvpa26MDFkGopvGNZ974h/CMvv/wTcMK40sXee2Q0az4CLjHk5keX
DAYg6zmD3apC1C9WaY3F4AnR0xnUjhaCbquWTjTZEzx75aG0BXgd7LdfN2bdj1o4
Zs4TSC45VJGmd/lujWmXw37RY8EfacR9mvJfvmRixR+LYijpMtQGjuUzhNUGAR1v
1ZgNXCcy/gHZ9B8zXkd/LmewwUe5gzZpeYr58UNbZLMp+nzG04WsJbKACYm2ISny
mcwfzTnx81uae22/HcdqBA1hBGc0xJiFZj+qAffCjDUHDAl3PmRwEW6zwEbXr4uy
n9Wd1jRRP4mXDcQ7eYa1IL6NUjAuUonEizxf6XfQGpCw9gLd2IEKAIjZWFctBAbK
wpk58YwW/gRKJmiQlZqkEmTTrkkwR41q78jx3EeHeE2zoEtMhI7L1zAxVZRqzlb/
dRzYOCHY70oQFUz13AfS5kyZ6shiWPXBvccelo6HprpDqYAjWNM1nkkgHe3lALVd
XpraTiMR/7PwwtJNU8+p7U8rWaB2ypMelpsorJKsvHzcTyOayWpwblK9CsQIDTx9
cY6kIJPyoydo56uVAqRaQgqK+lMwTOezYWj+6QLkI1POo5sZztiAK+RVcfpxo2RW
yDMAkZ+4I8Pc+Y2nbuKgG8bFJOcYROo74hmguekr2nomLGPd/yN/fV6sk1WLpkhu
sxf2PjDJT5Dwk6wIF0/g8TPbXJNPp4wt9fGoTESLD5b28UqmOv5fdOVcI+TKP6UI
MtYp/TgJWYURfOyfy7uJNeDWlG+MumuiINVexX3SJsgRMaAGl28OXDaR4HMowFzH
XY3Vq+LM3D30wgeMtJhkF9z8SodLgwi5P9JLzt+uG4nfTb1A67nRJyWxtw+2bKBD
HLM+eTa/hCCBl41WyetQ/09hfNoZO/dcWrBiGWkdxO6PE+TLpXgc3zszi1hJinw2
BZBarleZ+ueuuqozrjrUdYghYZUSjliaGTATTxuAwYQouCxI/NQC5nBwvgn1D7HK
5pzx2OSoAZs4WhpLZAjF04eyVM43HvvTL9LLriu/isIcoXg68hvxps1WEsI5XTvU
ME3Er6wFS4VyG87Jyx9ajwSCr7nI/LLQb+yuQDiT+hmMEiTjmKEQ+I3E3ZeB8GdE
GpLRqsbCCwV1tEqiIDM3Fp/4eInYjPPXIh23XudGkAIS2pNQ6TwpuDFJ5cW0sxJa
ACa9sY0ZUhEramwgwoWlMtys2jgXIYzYTuo8G/GKVrH/4qz9Lq4kr2CNVBMvoDlt
D8J18kutIjwDdP/uCRgwBNro9PKPZD4kYX5Dn11nk4MjSlLE86YCywbAHZ8WSTvM
d9/fskfXNJ0mTSIcI0DrsElaQI9pzylHs13SkICdOFcQYUceIBg1dlx0zQwfUT8y
0Bj/+BB5wI9VM1/SJk5AmQR1i6pND410VEnfdErEZsNEl/wU1G249DNdgAc3fbLZ
tKUUw61AXSxg+Hj5Y+eLLFYnFnnUZ+6jrOCrYo8KwmLLcqMgMiVkebD+/+9OgbZD
A1mRZy82hnaOQUMzB7hGDYY/z47YvnmQp/W8138CMTfPtqfzQiP9n8A6EKltajjl
PgWw4kamiY9D1RZf6kouex6z2vaJanPPenws8Enq0mmLdXdT3rR1gR6wTl7TPYpU
Ch4W6jRxi0KSDWCqKBa7pNacKIH066fibmJbdqD58YIQ1iQRRWrB69PbDcFRYTJp
Hx2B4GAFLBsWGKG6TSqEyO8h5OOXX9YOmp2hneCF497C28lOyl3IcTGMJkIyEu5h
mKfSOGz/w6nET0QlM/a4NwMXChQXwudhQ/pR2gTx3qDpp1LW4Fgg1x+dAs70x4Xy
ejpGZx+NRe/kFlCaMfWSrKXiRoXtHLyn13+SNFfDn41xlweeQanM9YyEQMv4zPvF
/Q34DNsoCEZZCqkshjUCSJM4NCvT7LCDT28Oi/ie1lzVaFNCHp56WIOhpo4w0AQp
dcEvsu9PnUCiF/E4uCvTdwIrglIoXAOI7vVydTYSydAJEgP/DtsFPhJOa6gD1DKI
JdcNuk3MJDQ5hatdeoTbV9GmNC9qbyOcaoFSTQq+/048dlB1v/+snFy5meYTGbCU
IqYtgEtzUfvimbIBPDCNM1M8Tn1FClDMWm/Iob1ipl6dh71N0gnZdO/3SvydO29V
pQhVk4MZTPvitqGeL+mhHX6cVtmVloC2rU9vbVJbGWHQW2/+IoN3gYUtIQsFSFBW
OP3+v5JXoK2Tde7v8b4We1QTR8wJ6W+mP+fQ1OKJ9Lc2vUts2yu8qlha9l1m6zjA
hWbafXiK+frQ16kotTohAsIE7aCOVi4bKuMUmTm5JwQ3Ywvb1omcVe23XldHqGO9
mfSJF5LnwL3vO6SkfLLlw7SEB9BfZs7VYJEE2YaSa1imAWs5w/Ilnhdz3fT3c6ku
0oJq0ritvkQuyvJcSvJvgF2FjiX8vovCubNGade0oR8R9slKvR6GckDgiVXZuZt6
j/vwS3cfxGUn0FUvdNP/EnsEVGXCkbMHcc3MqPhTBay743kc4LHTxChG3Je7/SZa
6vsZEE7n+PXkPJdpsUQccpzdAZdjwpoMZl2nQv4GOlH81W4MDgSqgjq9EADuGXTx
VzK/6d9LHIH3UtNnl0oIY83bTZZpSAEHvh3DrrKGAnYwzAUwfsKK347/SkzG+cH3
iDEosCpMe487W0XdFAL1F1mv9SQ9hWg/yAwQx3gGTqNR2vyaWiyJdswq0e4gpub7
Ircv64bJ+IwgvFPwHByuRXfyk73UI4qo4DXroRyj+NsNhaj6Y6tnNzDvfHPYQyRI
7TGjKz0yRJuSxfajGsEA1Fa+hFMazCRf1+p7V+vpeTRbcU/mZDq96YThdb5uwAgK
q5BdmryrWNHSFEx+uSzZ0dEouDqKUtdzhVPd2vidvy3GyAOefuvCL6M6gbGYrPqN
GclPpFT5JFehOvHkgNavMFoPuHZ010T7cCZKbokAPcGFTRalV0e591sksC+TQ1CR
2+A6NGYSGrw0/pC/PR6TIjY4YezNvHy8gxP4ZswyQDhgSzPO+dq8h9yCSgyILlpA
yfK9vXYzsE/7U4LlBwqS2msHrsSqrfvJOK5HB9a1orY2YEMZWQvRUPiJ2f5BMSBt
lziv4lc9gFV5boNcryvWWJfAWJ4VKvb258IVd1BKZRkyPE0seixyLPOPb5bOR8gI
4IvOHSxZQrMMyO7fvFy1cC0Mhp4GFLfo66VDL6W0jyjpD1v1hfZk+D7gYbI8+3UW
IKdmXB/QgWMqePZxSMckXNFF4SFQka+hfW7/YXcb8VVWPGUXiCfIWqCa8+6R6Rtx
GpDHZGxU6HcJK4A/r/Xd+5QKSXDdEWwt1wupI+7y4dZeZgrNfkA2I669WKNYkJl5
oJ5S51eFarIcME3j6bCUMLH1q8yasvpbnB9mPQafZJuknMYT1rrUZ+HD7j0ewN9N
hJouZKoPhYG5PP5KRW8+djnOcsuQYuhe6WI4tpiWdiN3pGHLQc6/k+eNxN9Er1LX
3oKOSnKv8CL2S8rgAbrpNNxvbcoNhoPwIkz3ye9Avc4rP7BLD6vsfi07Pmm6G7UB
H/Ca5jK9vTgQneGYt0qdcNUfrNn0qsR7xxxg/++kcHUUzt3mAu53O4yzeeBzJGCX
HUvMeZr8fb7vUWQR20C00HbiTv/k5tEgqQaJn29KWFfaC6huf402I8Hp8LwOOH1w
aOFfNso7BJjo6s83zWrCS1qAfgQ0J8AGC5TRfVp26AhTpUJvMxehXWqTWY+HXqia
IAZAvhDLjRQXaiFdBEQDId0dvuVJeRUAUmUM951Tdj1x7c6ZM52II1VJUA7A8KAZ
dFvkXkuzCx/L+bBbPi91OYA4WUZ+1Ta+Fwu09yDBmmK/20I8NR4sAerREP/U+Ceg
u4SJW+rlgoc+in0kloa8uWBmmz2tSd5fMRVp00yuKVhHSjn9PY6+qRB3KHi0drd7
XytYxDjsnbGXTCkRcWoB0y1T7hHQ4SHUUScRDmHXLJGIs+IR04Of3Rso8AUHUCqR
i91PrmcwvuYyNQkMIsKopUYOHW5IXm4lX0bItongItTOk0RFa9XodF7CZ0TArBPM
OC5PBVPfjaXO+pyFldDp7UsgKJ/afq5C6ifIVUIhaqyxZw5DzMzcWhnxUxil8Gqp
vTOvQWvrK08VklaWTCNjPbz0O+95Fv38in8Ho0R4JpfvU9isn85ZidOufmQIJRly
bplJNWb6fSZ/egSSj+yMkdVJTgdTbWEJe2HRsKdjsSI4ZWypOrwsKXVHaL9pyP37
LUEqdrkup+Ft7lKoH/dWdemUbpzXv6wpEM0IxU9ck67MuBSfRbR5QVa3owGh2zps
QvYCm6Nk0PauRv+bg3aV5tCvo3FqpqLQHy3x2XMZ5Qgzs8ly5Ak5E9tGgKY5NK7b
PvbDKmWQJ6AubqaTF7rzeNycQ6+JmZ6hxrhEwkyrVenxK2EJYU7PvAAN+6XJ2XDT
1VEoS76mYcU0jrcN1mhOLXvH9XqCi+U3T6BCCLD+h4VGQv4chbGrd2nSKtjjXzG3
+4Tdi+Wph/hFyrrnGzaIhQ+UdRRyHiCehFsWOjTEoE27JpfwOE71PC8WQzHq/Cu1
KKiSyBR6isdFccOmXKSEe2520R473MftsT/5rYtDY3S6KY+N18HD/gPlAG3NZs1a
Dda5iXoMrOGmzx1azlFmfXMdYubzmZr3CxUgKHfWZC8jsCRzZuXJMqpm9y/tcHHh
X6ve6K8VNSLxqQasfc5G7i8aJhrz95CTJ7X5I0zbbOSecCwtTsvPaKuon/0FvhR7
JKM2aE/wGPl+2FyyUhW/QCXb3YKFy2Begeoq7jkDx1Z6qk+Ih3WBS6TB1TrOzzEp
/ZYzFk9vIok/6WyDzk0Tr0zSM2iLSQpYc0wPNYeip0mYTI4RshK3Ev6LGMjR/iPA
HbeF8U5AYpeFU0bieXuvf2o/w2ihFiXDmQLKPsXoiP/UWjTVvnxqKDiVaSdSdXYB
jpyfei+KYomjV5GC452XtcJtLCBK7x8RN2tSpcdI5vYXVe8I+rV5HKFigYhp2NYK
gHLwJ9IKj77h7oyX+aw1Qo8J9SNdX0ty5WleN+3/+JazfYdxWIqSkvMDAddZeEQ+
E9CaQe6RXBl7pOlSg4aRO8TKyNpW8Jm9O1RAUoPdJ8C1ztiW3GDIM20ld9r2hObB
IZb5r7rGbhbo++nuOt/HaxpueOltn5R1fbAd/ghHxSsxVi+3W2EhkrAJb6GwoASC
4dUAEvy0dFimt7r6wfObG8WQXCvYENFHP4WUAzvxPHeEVx4KlhvMPXiQDaW07Sd+
j6oz/i9ZnST8OujRS1RK0inEtgKroS3Nw/1faJFWpIqss5faLuaibywLANPiz2id
ikDPqKBsdUEy+owR05JZeQ+6uLFEAccQ9AKHfgNztgBPFYYIdnudfFo5tZDK+vhg
/Kk8C6VOt7b1cX4jtE6XNT3iNDyx88pBk6cNpiGz/pUAn/ocpwoteefwXR8ufgDF
+qezTOVKdAD8rdh+HcoAdcFC4unJDdhmOPtKlCrsuwn2NTS+YGfoYC7dBwJLOZd8
/hZmum6S55iqSmS7kGGx6wb4ApPpPXgnA9J0pGokjl1KpS/gRP0jFbXsVuvrSg73
6aAyyqOiBC8/+ZsiXBxInpBCvl037AEeeBOWcqW6o3yxs9Z3XAYUY1/Myj4VbiHm
Rvr8TmkXzGP0BOrzj6rTiQTFch+L+iTEZENbYdbOsXF8L+yrYx8wBxwa/v7Qj9RU
/WEi1AfxE5ctUXytCSzgsClV2/gx+7WswyvASRkIK3rtU78OAkfq44ehPd1Hbag5
Hw868WegFinKipOcMJGjWC/3sJWXxSXcqliuoELxNT3UGK6C/JYlgfDgedUPtTQx
lFQQYLonVvciCed0cSn4b1T2Rfmyd4gdA+8hfpLbwUFDc92PI1fNC3QNwikFbNOJ
GX94CWG8i+qWat+ucFnqU218IMTeI/jYPtF4YwhAhszzh68jEFVwU/TmXEojVNv8
WyAII6qHDb8718a1zqc5y5H+A/672N08SdCcAT2vfGtrhDCuYED7YCxlBrwDbPo3
uTlLNoo3x3CGo8OcRE4Css/0wZ2SdgeuOL+LRZw1abwPSN/d/D1GoIDX0cESJGcs
dkdAKQFkTO0zffBDs/m6AJLWXG5qAACRFq4USn5SgGyMTBkcXta4WeIx7hN4AQrT
Cr3ubBbtLqnIEzXAFIhQmJR4V6nIFD4U1NL3GnTg4lOP9baf9bXM00YCEcZZmO6o
pxJcqwKezRsyyF+eaU3Mzy3rcEDzYuqkaBX2RBbssthOAG/cNiYbuRSTRM4YusSq
LBE0/4wTR1DmBOf9nDXguelsOWKw9KPcORJunbwfq4LaUdMB+GH6NQz3Y9QOpyJb
3pgY4co8f0TgYqTvtifoqUR5mWmMxhC2ScxPYywROP7QqTfkEN1l1LGeiD6pOX8H
vef3XvsiaM2E4AJ3NJvJd5HLVhDL4cbK82ZxDYvpAjtnZnLFVStCr+xzhEmeDGnM
eXwMW7Sv2R/OgL7pOhgKFQ6CTlct7Dmu8c0GAnWsOIW84F2S7FhhDrdjo7xXD+11
GCPcdVuhwqtfxfo6g5f2ldxPSzs/EsRYt5TH+3aQKbNqx22QcAiF/AVa1jVVz77a
2c2GjsU9bC6y3WbBRIbTKicotTFKyITF6YaWy9NOxX2Kr4Ea1gVw0ile9Yi/eL1r
s363G/6rzWIfevYrdowu2xnl1cIqOMnfapEzVreY7KyIcsIHt+KzUBbsEhqwPs1j
bSPP9tbhDWx6HaSKRVCO/VF1sSPVO+N2Y4zwynvyLDLjabiMzcn3+oKssf7XQb0O
YCXRaGf1ReM1e6pZqRP72R83TkqZaTlaIGG2yrdKQM2/YJjqMAYRK+UkqjNmRcV8
7b2rG44Q13YmBs1vO26a9+HExR9Gjf+QLytwO2+pxFaksWt0GfnqeI7EYRbE8Nzi
aLrDXbt42iWO2NEhutxY21OWjKo7QaC6uSVib+jDKJINXkWZKpJgPaMKXyH099k/
Xw7xIdLgOZl+he5wR6n0jUcPd5X8pNW0dxQb0rKzSYkxLBKnO3Ps/kTku9LXU/cr
q5GC4wXMLceb0WZ9+SFLaorPZDR+2gGAnM+SY3P/c8kRwhYPwqU1DFkCL+zMsk5m
JX0ZNzgAdL9PjPzttl4EasKAIT7sH4sImpH0aezRpkvFKF6Tm8RwtZUVFSzQSACZ
xqDjjk4EFU4frBPnYcq1s6+WiSpAdsVhp/6qIUdxHBIXQQ+cF0KtMRoAIjRdEYj2
+ibwcck8qggfnN6NTh6AE2/DAnqNWdo+Iom+PjluwMh9C2Q7jALAKCu+XW5POCgm
HDYQkEopXd597QTJilwXdqHNd5Cl1RxrEjJU1W7gIqmvuVFRRAA1NcRUppk9ZXG6
F459Pb07soMO2+GAP1I//0NLYj0HnoaSLJxbOc4cjK3gSMpMZWF22TkIeANQT1iy
XAUcU7ff7y/9qjbCaYWJEpGmR4DZAskYyjqVEa3VQlUo801Wj3ehsvpw9fgQUPQQ
YMKvPVdZzOvVXMyISSLwQtd1B3cw9IPhoWZxwtCEn0gOMUIwL7AvtcD0z+F0mt6d
UlKtcsvT3EZUAAJcWH8zp0c1qMqfWqE0Pjww3jCexaX9gRyGZXkovPBhQN7PnOHe
WNFSLmFfP6P6ePcX5wneDo03BSv7zSw6KSfPrlAuESh4iNfhl2OERdjq5Vde+xBj
tkArt3QNYPk4gmVK407ZRzV6LmsL1AY1/bkAl/X2CE7KJMus7DS6wB9vlAJGeOjK
GvsQcxSdPXqTiBYaY0B5RVfLiEIe5fLZYCFcqR6Z50dgaDSAs5T4szYxZJdcFppa
N3WGfJu0V93ax/3O5sMyq0Ci4xgGrRfg4qsQ49J74SPVxptSGSUC+Q3eWYAvMlwH
shUTthu0NB+kGKT2G5qKpl7ZygBlPzFknb2fqpx2sdDip13xmdwXiMf29lOVh4hb
+TH7h7k3YvsjqDTqmZys1ufu8OCo/63r+62lTh14Nz7kM7EhZ0Ji0HLeA0UkK7g/
2G/vUVfWkX8vQgiGUpTn+FZC8sLjDPDYUkdUkgk+O53u4LxlxEeKsBCyZr7rgnRS
6j7LwsBmtu1tOyQSSYldVenlzvnOE18+PJYOlEwV4ZMkkFcgemRqwzNI2vbPfbZQ
jJSpjmdTVDXsY2Ptq6aRB4iSE5Shn3DuWYMt0b7GTSapa4hGk2RKczZ5taiykJ8k
0C2vqWLlaebjfktRvQ4YpJ0yQJbIPyaJM3a/gla77POBprAyXgZIyK70Ox6oy+kA
8B2dhHYtcj7V4DTba6ilPWXmelPNjRWx0pceh5GlJ5G65EX9BpgV6+NBDEdcR+E/
V6fTEc2qaVJVlfckzqieOs0iTLWfWfo1inQSW7hJdeB8kt+Z+YDimnqy5CXxaDlU
wbpyC7VPUjKivRPgSMkoqfjKAqfyYkYTqJKZHSDEMqwxK7BFKoNMDi3bbaeL0vlw
2mgcqF4gajcOGP8rtP80OlrH0xmckEvmga/ah+g63dAYgs0ZuTIsB0wwtRo3Ijqv
GCZXeIAu6sUydrplXgd87mXoMwIobCH5jQAX7Obgn4flAvEISQRX3/JhES8uQc3V
a059DaRFfdFCNaFTcXBMrYg/SSOucdI4ql0wRri5Fl1ddsGxn10i0B21PYIZpdJq
cfv1MYnG0MC+qD7XaiT+yqG7mmzodPiqcuW/w+rBX1Se25kes6tGxnBdAfk1azOk
ufW5eQnTGWa5sDq+b9TRR7cS8aCzTmrNYzf4KAO5Ig960uX/xZ0Myi0w1/eouyMD
5OenyVNkitF69vNzpkoJIy/R6LPnwQ+7GIcUVSj4yDePCKlRKLgj9ZIisOl7k7zs
IFyoREP49SA0mX54AwSXZW+tgLgo4h/HYn5EYKkrTmEmQISNwHgvBTEvbPX1YjxN
Sk940iH0/FNoI1xgw/Xb7QK68OOUmTUAUBWXVffLFOZCVjxDRx6faBuk3YiUrgaq
+pBiezBiWRgnDUpOmGPW7C8/H1FddKDbSwKB8QckAGxskutWtyrZtb4DNct1l291
vN1dreEbHAL0/3jBqWWJyBh4NW7rUswDF1eu8qhZSdaSMOGAxVUH4hc+1Fx6OwlO
ILulvjmYD0Xolr9wEPsU4NGFXO483J86tsO3Sv/arPlo9mEul0AmqZ7JSLfSo+0Z
fLfO2lVKZdeqDACVKXVBmNHRNQVOQ82ku4cC7A8SW9io/Dg/ZMoY1q+UmGnkKq7h
0mLalynjwbYb0ygKnw85gL7Y+XKpyWmVos9sv2KU7T1Cm4V1D+MHSRBAqNhH2sPm
UxxYCn+LlHb/vNVD2sObp2vtLRJcN5EQGDQJxLR93LW27EkmXgqbWrAATxLJRskM
uA35I/1IAZoz6a3m5H7eKkpoy5dbcb/hs6hnpPeOJCVwQ03+qEskN8gi79xljkRs
cNPGCZXuMNvvWGkSnWCuVLQr/t0RTELXpYWKWDAEVuAQGeE3RuNbXBhIChYPSlg4
UCvVuyMddUyreah1uxPk7tfZcKnbFijny/IQOxYiSh9m1ohGZjfKsfWfsPCV3jeG
tGelHJt5g/mCUm4gAfsdEfeRzoATKTs14ZfATRlrzmw4NQkdnvYnehBc//SxV52G
cZ0jlbu3YwrGViopCezFyDZwfrN4BPJu6MkuduoJSKsKtQcXhUn6jwqoywB4ysY1
abbZjoBe8aj3u349ZTpD4jm1IgNIC93mw5pAGglovJGxgrDKT94KtWLKvszTsxP5
fZSLp6hexBbaU9P5dMo3pwy9uU7QzjXXlWuH87I6spFkvcq1ON7L+YLnngb9MyiD
pHIeUhAzBMl39cPGF+/jBoKwzznOSZtU2dmwfPBXOSDcgi48P0bnbll3weWe3O6K
N1c69TsdkB2ZtcwZcZ2g6BQDUixHoRpU11UC20Hav+TDIF2Go2LdpNULuTu1l+9w
Ic8TwFYNPR3nQp/b4xB1Go/GL42MgwY/UFYY6TWTaOU4R6/MdEnUUZ4fgFEITn3d
eXvIhbQ4w5aGVGlvLlcHDvuS6y/W4jfyyE0G96qStsP9LHfWOCvJ4B+YyLUeZAyz
ShQ+5ku4fvvDufZ72UiwVlMLWvgLHhu0HTmhYqRAJNXWgZ2DLAz3X6sZLe1IX3b/
5XhVKaqyF15fvPqsEpZk2iC5KATivI6UkkO38bYBHrf13XuzRqnKGgN1w081lhtx
hRUbaf48XnXbccCnLnof+JnQ59dVcph0I3+Ew0lTBlFDfx5PR3z3FX3dlNKEhlUB
8z1BASsPFueOzCux2DGfBSMgQrvTYq7rZ/v61GS+b3R0A+7ZYL8i+ieDKBuGkeFU
P/O4BvWI6KozyVtUUXE9fi9SG1MBFswhohMWqi1CEeAfl/n7ZVpadvIHQMwFeQAc
cNLY4wp4rlvo4a5D7ORYbRjiAXBCYCXkvXIekj5PFN1BUxnKkExngR5bZH/8LYVK
g4y5dOCnjQHX4frWzBqv7AJl4hIXPqXhfQNWMzjSpWIqiyN9WMy0klmJgTlgKr9t
MXOjx1W0Qnbm/nYVzhth9NcJNwnJjtflsTG77XAX6x3IfQ3BpH5ZRrq+VULMJRgb
e8Hv9eXziMGl+knj0f/chgMo7BQyzradRSIX854nqx3Xdz99Ft5YhS8FNLuGcKTR
kUCuosPW9agFxSbbUZxH6z9chaue3Z0cH/vtbXnytjlwqSZh7UlKUsNOmLBDD41Q
keYi5SL/iv+I9N8OWrXJ/ywT7EeA9MW7Q7GBek/a62hHjmf/sBmQPaP1aLFZk8x3
CTgen4OMnbYg+Rdr4EF3+EvKG+0xOeGLs99vm+y8MSxv7epYupIWcLSbzmGt/v+i
6t1CtHrKyNkL3qO5kRgPTGp2Banv55QefHwqbS1IeY8DK+7eELy5eZ3xbjTAKFnH
NIFdNfHgG4fxddq+56561LdDIu0LGOJl7zwqtiXVHlUsE8rVIRB0+SGv+iNM4Ywh
CGlwMDxfFIiWOOdzj80kXQzovpF2/WCMrdOVOj3zV3NVzHVGShzd1eDnjmlgN6fM
+HRtvE5M4lPnskXMh4GPoduIRYMVkVRQtlpy16rBR27gqglodVRzi/Nty10cpxOq
pgIUgWUc0s9cKAumR2KvdBLEioW1fXqZXyz+qbjMPriNej9zx+CokZFTfS0CChw5
T+tlKKEIjezKG0O5TpI3u9JdqwhbZ/LrYOE2SonB8gFzUk6688mgxcBs3n+fifBh
1baMLv5yDVykS9vri2G8PegD3UTATe6uQsENdRK0wxPfgxm7NHwimLOKPtVp3jVu
59XnLpivcYuCDP81TywBaz/w7QZubb0T34Pu+F3pr2JYo/WUhmnkpCqbykmOKQXC
G6pOO2V3meWljiw/Zz+eVr6E7PS7JhUg6eXnfncqFG964YSayOXfJHA7F7KUOOW2
9MM/bfMnFEKWS3quuvDJQDADhOx8LFohKtXnHaoEzgFfkOy3FAEMTyMyCv6Kjbkd
+SFJRQTDfjl0M6enty7+JiaFEXA4iDG9GHXwFsRyBNhIUlWZrCsho6Az5dewthrI
mCywYd++yawW2IonvU2aEicoO1FumKeru4f7eboiGvxES06eWjTKfaN90Eb6YKwA
xrIoIUiL5wQZbOS9Cq3Ir8ikXaQh8HKLQrFZaSXyZDfScGFnE2Kitmdb+Wv7JwA5
1ZnOIkaj0N2ybfYgINdeBjKC1vb6gFNz9VFe2j964+pFnyZBK2ERm6qTbZp0AMuS
sacXBtsLiDOMmdd7SfdUIQNPrIcWNwFLvh1DYSDWDej0FR7+RGcv9jz9SG7tuniR
b5PctcxtOOnfyzUfn8cKeQ7V3vX+WCarmjyIEnF3OmqED0euohDKsDEmvNGj8tMn
3CzlH3b5+HtR6jvgBn1kcyZjHbyGgmRabrS6VLawl5UXJgXZUCOQYOMVJIdWmLeF
sSa2xnM+nJkSJfA3Tm+eGLsRhQyRhtB6/eGZPPI3P4hxr6eP22RmWqsxdOYhY880
+bYRdACy+J+0IPzJz+FGooEdRwXdfFMbAJ5HVeHXHbvDanHM/Sr0i12RqWxCYUBt
YaZUNJVtpu+zbYBM3WIAI2nifD+7mvNVDEWjVOmii4Vv3sxRTqVHAE0SrBr1JbkU
rzsphIYs8xJoqgyjJvdzqwAiPgNMSujH74VCwLpY29IQqXl0K2WuQqJ6A8ApI0dB
agMaOe3MmHo+65UhFv+MIyH/iSvlBh3kCLvAfeua/l4dBiWu9dzJdBmnKsgL7l04
pVE1xkqX58rrpLFaPQ2PN8Ew7mFBZ3r48sIIx4UdrUTV9E2XKLNrLSnc/+jftz+K
0rd9x6OP5MQ5mZs5t2YivaQ0/E0umtygniR+mdEfnH/Cb05f4D/KcXWyD5esITXq
VnN1RFIc4VExAYrVcd4qcsC54mbLkfyh7GxMMoMJCMd/f8Ydov7jRMSKErRBWhNF
TVkxTXIBiTJaSJiJ8rLjH4LejVzuMTfyuRmor3HQh1jmTgWX5H6f1ffJuJm5ghnx
OK5OVji2jhoGizbns6gS/bZNcMFZibh9UVTMximDICv+bPEJBX29tJANoxc4oIsy
xPjLSVq6jxSGKajgeTRnaP7xQ0AxBB3YaJbr2DxTB855nkXWAxAsAyOIy2pLchJ2
YkRw86mFXvAj3JuJep7A9izJr8G9G9KJ2cJIKU7j6zUNwOYYgP7s0Kgcn9gP1IB1
GZAD+yLOhkVFIzs/92HSI2+WFXQgwybuLEeGcK/lYyiK5XT3nU1zWOfdjJT7gGfw
4Nh1Ze2c3Zr3i35menodQqnKQmm1YI9aKJiM3jdXgGvP7pn8bhEyxwAF89dBc7jG
LB0c49Y8Oq+sJuLv23DNcocVpE0+yohCTyj1+Xr+U20R/oqdPAv7nYBufsDkeJag
hXNLT+pugwvbTmeiAuEURrGIFzyZDRaPP31ZSjj/406+qRoc1eMTiqt1XoMWyN6X
45ZEn2TBQZ/NGIaNbD0YuEjECtv/Si0BUi2Jm1hA2ikfkpey1o0TzIpdENJH+u7T
PEKyeAik3tDRJqGsBtpn0fZ9mdTcpDh4wvwuAEoEbt4nzMOGVQv7wQNyvLL+KPwc
g/lWLGAFtfZU1qdERzqPr4IdMbnTfI/yKFMEqkExbxNG96uwSi/FZ3hdr28k/hfG
sxSg6uW86VtawNqfTLetsY6Be/c0eUsxZem5BUA+RhCcwm1KBWBeIEJyzJ5rxwTo
KfMoVFnjK7fNdJWb7veP+HXYHHy599hm/Xaw17MhzOOgCQoGOLWSJIeQXCLNl7Gs
hwRdYMNoMxiq3ah7cO3+sDg+27XOycgKHJuPofRzZocBQp5BeZJKGhOqYNpbtw0v
YWF+uX7amUsZe5UBuaT7VJspI1LuL0TgocMit4xpnWI88JITESJAtuRIfwMLvRX0
BT051BYlKogUiJSjld11snqBMM88DBlYoE4dnLm1FmQ3PJvkf7wz2SiocCAMhxtL
GaF+pj1c4DU94kN9J0PDe9PU3DPB3TW5HdCbaZMeoiUXW+OWVtecJX9dP8VOCJMm
hVAD2d17FRxvWcPlYbVXOQh0TtQLmPvV+vVR0m2pHGDx22xJ6US+Fjo3NHX10Qk3
BjWvRi6L2XXczaFMnLJQi7nOXjkkfSW8JV3kEF56jyktosRmp6t40DnoQ8kNv+U1
TZMHCGacV2mVjUNyN3bZWS0MFcMB+Hob/ttIKb2UQvbZhIXUt39xwGr70v5CSdzT
iGY/JBJ5rFO3UekNSRcHfl9fEBrUOl31NvSOUZt+HXa7zun78jpD33Mct+vx5FC9
HYLbw9mbX3S4iwBKQcJuMg2hhYpyEZM4iDj3sV8GjZiGIqAinEBn/2aDyB+wB8HO
Dc2r/edL08V5IuQ2zWJ1SQYkhPyFD+tO+WyFpHBnOrmiy4HQ9J+Ma4u0PD0lFFbO
8LcYqpnr/T4hfcYCmqBivxD79koMjEJ66mPflCd5g9SEZ0giOEpkpXa6zxOnKwF/
x9eckCFaONmynhrBrg2qmMSHRZzveIzy8maEb99pHoE6pNCx+YqJAp5HuRi9iKmJ
GUhFLQrHWJ7JVwFIeJLpAlgIXLCFPoU7E1inGjEtsk2mnqwin5BWV918McPhEfhQ
lacAHtX5hctpFpgoAt0lbXjOAuHgnCxeIHh2JP7MtCuv340CpvD+leSfkLIS1rOn
8bXAd5TQOxEGZhYnPjbCF3N1YJm3zxaNXQljEB9UkqvuP4Cdw4Bm+LInpvs/aMgm
7nrF8o5ax7JEJzprM8QN4qpos37QZ0qUTTvFzXH89oCobGu6PEh4J9x7/N2QiXM9
+1Wet3Eg6gRNkstmuV5+Z/Sv3eOWIGSXdoWuAwg694vYCHSSX10W9fzTQiqZw76N
tpqYWNdCBiUwL5nlgy22G7K4PlEK403OfMKB5ZHYijqxdS/16eJmDkhVPg2wSyQn
BTSr5G4HdKTje0Yoy+cp7zGyx+b0I56qqKOWoqNKfEZid5lgAzqJdTcK+Hb6zFc9
NUBGXT2G03uDoKJBtO4fPCJmXsADSsSDOFz0xy+pQ4On7aIYrtLy8ucoSZvLmwuy
DvD7/1Sp2rvYcr/F1VTQstFk211VInEg3CSmibWTmc6krN0Lf+qg1dgIcYS1DQcj
xoRtYvaRwJ57mNX4yH/Vbp5vLcNdBNVuimiVLmko4CQUSPqIRezga0Id6xR7YBHo
kmy5xhHK5w2fVSi8HwVwZwqGbbejtoCF9pOXQ+mOqwoQJfx0Xj/KyJsZghUoThKq
ARadzcfk3IxuugkrV/oAZKTXvxB8f2bF2B56m2+YKD6M+pW1OVPf2pDnJ+R9A0I9
2L6WxlUyfTBglkU1zT+QHxaH3icATpi8jGoE1E/E9MiepS5kBY0JPUYzxXJWdUxV
DA3a5mrNJFejxM3n5dFW9+8b002eo6lKEvQTeSn+oZMPrPAiZarnhXyaJIdIT52w
N45KcUmRNVf2BI+/gDp4GySvLm5fXUAHhtFI5tRmw+rDozKXe4h4ryopD6T1GKnz
sEWgR3wUfmKCmdqqipeYU36DfgcJM82ccRlba1X9XVCY8Tun1wLovMnZT2IsRBPi
lETPXCjHFPEUW8K4ydoPFCVElmH0QvIDDoLVoIQ+NiJv1aebm4XG4YG8LSpFAxus
LBqB3Re9A/nzd0uz6TQ2PM8Puym9XWNZRNxMpJ9gqhMwmug+1d9Riejsp00br1qW
UqANJlkYDwxjc7KUKaI4DupRfLcRuLXuL3LkPX9/mtGUUZQizjW0RpALyEdu1eS3
9VEi/c7jgCVACijZ0nEx26sJIZn39Ps6/3utbcT6uZ7uxWnlJV1jbNTC4HK1mz91
q5lwMCkflw3ctolxrTwjgGMqlxdr0j6Oh5551O90iyZVwTHiIqxgwPZlCFU/HfUz
2xhHpAcVY991JrnCYWWfCXzYYc8FohbA5EsD8VZ+UPeTTndUDOVpi2m+o6Ab65Uy
55PxYb3Wl0aBKQYXjiJg8+UCNs/IPcqp7d7n7DMmsZMbgVjPJTNdLwjZjEpkOZli
0R3ueTpX8GaBFd2juX6PK8R+KoVZ0WXs4a1iCmLFA+qI01gd5W4fMf2NTbMANQwg
dlPAx2d3MGhMxBb3SkUxf9qNLWUpMyBgXXo92c/iDU3HCebuwrDBZu44msPQg3xl
ZOAdJENU4Aef8JXu9JE0eFJf94sZgw18oRnVq0abMQ6h5GpWvx3exlSzS/yk6Otd
zfp072qaYfBvjlWDsOPOwNeB5Oe/jAw5VuGwJXL+/ecqhMaBc4JhgqZL9VAITaAQ
XW9b1wN0ba3xmgJoPufygMkFZ17LAguapK1bUHI6Ml7Vort0Da+mMmzI+54ri3fu
uFyZDlTEFTIRazcyxVA+l794nGK9lzGOn7inkdFqKNp97jtagdcEd2pKBRtcKZHW
uUevLAi+DVYmNXsR28nlkAQ0XrFqBkbdulgTH5BXQ1BgeNAbwwu0CxiDXB4fifGI
9+71IhKGJFpzESsSqJBkQD2HBy76LEPkNrQYRTJBufXd415y7W4d00mhuDl1bbeR
fajfsxH4CZBfvY6RfPyeOsFhft/2bsle5agqyK2xTpFHTC/UEja79lfuTjmpc8gF
CZPr75H3WTGNHSfI6LGlfadKEyLNZ+nFK1FVxOyonBimNFxAKsEnaghoDDHpb3yT
jnWsBCYe6Ler2N6fqbLyTYgVxcIxiS7CJHaVzWL++pDlM9RLHzzCMDnChuapDFrn
icGG9Ao2cbTwgOVycK3qDlvacpeMVrVKHTlLzsu5RdZKOACRMI60biMxnAWHN49x
2qbukAeoT2iXv6hgGMTOyX+XLPO8GPvwaZaPndQkT/eoE8TIbSt8Sb18gGFquUzZ
6ZmULBQwkXojs9HSzoJ7qs+SpKfT8w6WUKXBQRoseg/Nk7NbYD+HHhAfFCsQ815S
SjH/r93RHuwK+kghDnjYuDCyYYQNq62JEdtT4k0dh+jfIELbKNzBlkY4yGVSm1dA
lz71xgFjnW06xtTSGGszaqrUYQIVctg3ej9WFmNI1/U5fCOHmJ9Gmycf+5fxISuw
A/VmbTeLybHQYZJzGtODzCh1HJGpdILc1TnEZt/eyiO0UnHhG/1Loagsl2nwbixG
CGVIubT2WZg4QS5LbF3pNnEUMhY85p6yuxnF22ijNjM8xP4cmpQixP/REaqfcH7o
5URsx9mdhRWGVzCZIKVaA8GPR1jQngrpIRKYia8EiACLWS9gCWxJPGdCx2Zdw1tT
flEmpmMN4sbAIDQomDscNBV3+ObSk2Eq3khHiE1YCtura8Ln7kybN2MP/+HFdgnv
zxdUI1RfLM0WfZw28OC71QKV4DJVzZe3yV/RC8jj965+Gis72PqianKm9FvYeiRe
W4Icmrx3D4teo1vWAmMiisG9pzDbrscssAzbAT9Z0owzeKfVjvuAokGG3Y163Zf4
kAWnjlONvHrXQbbRbmyoXHem58LxaxGSP0S/LqA1VgU0lISsNkTpVUuRLoLJcJrp
OHCuGATrZQgge1sME8wcGZaoG6NyQiV3qDhq7FLod2ej6Qd5otuZ7krf15D48mA1
+yqNAYBIs32UkMTfkOEVf1xD7cD70t2M3n03rXf6OEhl2WLwYxG93h9mOi5HQn+4
JEc9f6u1s+DwNRXdVmlSDkFXdATgWwu1w+KKFvYYvr1HsDhIxMVGbMmlvAMt+iJo
als7zKBwmyux9NmIN+lYTDhTILUXm8aZ2wFsnO6uBwJ1j3iKiZ9HC8JyIUvl6wQj
40KG+cKJFfY0bBahJVYnBiXitFJiRspu1CbK+VqFmDhmJDKAQGVEaMdLFzyM4NAW
aLDXPwneHoMGWnzWHv007yZWgrHXFtZoZ85vAZJTYjDeaShJFuhxoJUG3eN+Ywt1
LhRZa17mvHqdPVIkG+8J91vdSXcmuWeKEXbsLhCyul8GV/f8Zfs4JJwkN88uRdUK
rtkDwC19MnESK/n7fmKvALvc3XVckC5nuYN0zupUq01t4f5zgUe1GhGOQMCXPaYt
vJ2/MGmLEtFBgTZFU3ltVAhqujcig4jSHOBjrDKN/RZU5Pghsu7g2GRqXkK2bRjA
NqzVW7oQNQHVWObqY/n/ZB/EqhDO5u2uDxCnYd/8U09V0TiMKta+WhKHhH+68p2T
P7lGDEiWOVlYoP5Da0qVvnoo6oO83PT8adZAxOSvaE3D5LBHV1TJIpxRhX67jc0o
EjLDJGV2o1RnPSRLMRP1M38WBEDfV4xd7yrnso+mMpuvwAzMAYSYfmK6UzxntR1V
oIa1bH/N+1ZbsxKMxF3FwDKZiDuwaWCNM5BLpVeExARI+fCVfHRQSinJzonhvmA6
7+Yuo7Hc1Nj0iLKn8WnTfpH+IEEF4L+pNPVyqkCcgmtm4AfsZENUf7MEQrN149Bs
joZ2g+CalD5SPdbpYubcVFzBe6QDR3psPLsP6oDhFc/YOCe+Jt+5++F2mBWt0qYo
Xe/KsLwizZLjBMKYYmqq0CMO8XXK6x3gv3J+A4i8LfzblydIUWZfsWAqJ04rqq4I
bCsdM9pUDllaKLREG5I8qiYqJWYSGaA2BDIljc+loTGIhZprKhXeQwSQBXcXDFVk
sLXuQ45Jew6zxtn786YQs780NhVzUsBfTmA7izlG3tTuBGLBWfW5HLCdZ/dgJVg1
iMh24GhexJF+E/GCiu+3u/WCwtHggr+02y/myuSIUNrS+2gkPzJHyLyKD91AXJBU
a7BDpwmaltvspvgSiNGpt1xIo9jzicx8RSm0W+ar6k64NBir63fX4GS+NSubnLa9
9IamOcB/DiPpImaxIdOJIIIcoeDJhZa55kx42Wy9tAQblH7CmYz6wgKzZ1Pl1/oL
YYmhPH1t7V29d79Wo6aJKsmMs1t5BwFoWteiHg119XdYUMoptGACf9fusnThmHxf
y+pbfavtMU5/xy11t4Fc3Z9b1JtJmo/2snaoVXuQFVIYUfpREVCO9/1jvsI/RLtj
zyfUL4ktcE/X6PCjxrz4ASQ709rnSEqyYSVlEenKJF/XEocogblhUrUDaePHZdSL
FQDRhM24r1SJAi4cvVUjn8AzRtIvTO2eT+uSYSGpfA6m73l2DT8bESvdnCUm+TrG
vFynwZn17sLPtDZffnwbUVEeDpL9kbxVwMFmjzxj/lzDyd6zfPzEy7aLv977rZW9
VLH2ciQPkpHry5UfHo6iXYf0Qm0qSfSvSPo/k6fCzLT5Vsw/jy+xiEEqbwwur+yE
WBqmabqSs8vtdmMCH4QCPoasKXMR4HTLdNKJ0Rl57u/tuisA+Un6EkjmfW+J4vcu
qmJzrBZRHiTlFX+5aCpevyV4QGAbc92q5TuGECZT1LldCcALzFIRDhkqpKtItGsZ
z8dh335ss0o+9RzmR2tPs5dJwvaek/RQtPjwCbkWJdEa45QQRR5YzrXmjBXI7ctA
gfyYlfP9f1sTRzc/leCzat78UyFK9B/AXF4SO41E4v6Q0Y9ZmCVpveJSZ615q6RD
qqeCl4oaIdaKXg22tXxlRRiK/3oc3wqiZe1XCu8qrS8VlK9CsvII9PWXza1Rbpsr
ifnHsulPLmwvU46IzgMCFN5YPDYASFg85APHBYc/edVWXhJYqr6/Dcjnpd9oB3AQ
CUt8at6M58/CNiKvHDy1Ydsd6Jux3vsNqXvMf1O0QZi+bd7CuAMgCbNa6qhAUfyd
ooSDsRqwPlRomT1DO7BTJes24hVaHk6DncKziNQkfk5s/CvAzEMOsAcUYKgejk4s
1qa5NrDEQ6Y1hT6PloHGab+nOtxKN6NaxvAe/Vc67wdwOMlCuVVNYpwJpCQvYjoe
Dpnqj2it6/75v5sXVUkcXmO+vKmTZBj/0q6ibrz+UOJ4caV4Fjm41+9V7efl2aMT
WqXicPugo/f0OZAc2RmC5vQ+miYCweQ3ysNH/gmWIQOocECug3FF67xyf6EoF4WZ
lsSyFCkWXSDZdk6XEP4uksqN9VMjPc9MazcwKu75548cjICRk9J/CuByRv2+Tbhn
dcfMycRAT9MlLDjIOliuuDfWSDe0UogvkhF4xbuV4Cnksx8PiTEXxVWnnvj4EDAs
tYE+vxnHe5AcOIuaaAM5aetSvJhP844KJhqdQbu2/x9nO10ikvBjIr3VRUFH3jNu
buiyl6/D8kNjD4mkJCoZHrIp4ZXGM6d2yYbv9jMxKKD9umjriSjV4Z2Igt7MagAQ
pE+CA+cEVMHC5hw4zC4WU4URE0v0qk558JP+p/l71Bblf9ozS8Bp3JGVpme7O5YR
sR2zAGLOLvdsD7uZWjycDBVN5ccvKJbLCd730aF+l2rdpEDss9jX3IbjrVd4lTs5
DpcssDuTqh7C9UgW3mEt8gzM5yT2qgtWfnZT6UKfX8lHiUxnSiEFnRVATzl/HNhI
fhwRAxQPxvyZurOjcmUk8neL12OezuTL5y9Q3XTO/a2pbqKaGE0PA4pnbVPsNbPQ
aa+z3mvGHPk3B6Na+qSEuUDE78N0X/nj2DUOGvZNVjKMckXyHvwdAzj6r6bS0/XJ
1eslzb2p6CnsOuTOlWQ0lZUnTPzRYWGndLRleUT/m7PpHF9NkRd/uU9IoKNf+8FJ
9KStYMyOLhmSc6mG3rmbA+3MfCzVrRx9Wqfy1SttRsl7zR2x+sQukIdghfJkhga+
in4+UbwZxUwxlqYmlV6BikR1Y6z/u+wAYbVxUjskkRyQSmUTm5cO3SLnyYsgCkPx
mBPaXd5OAy4QO9j4RIpesve8aStZcnRkeiyeaI29yO4lcWyMuePJs9R5RJHq1sh7
ZaxqvXMm/HXXIL0azZXBvJUyt78Xti5rKfC0iKgSb46hA/nHm+bwZ5CMC34+/BpA
Cr+AN+t7bahIdLEMeRWiYAqXQkzx3Lm+7WdZlj4VqLtKCFJyvKRabavcDnq48p71
SHoV2ROLIU3EpJnDusECZtHEG2W7X+Udq5Wul6FAYnWqaIzk+P719dJLyjCnUC/k
0eb5Jho5RmwFnBOEjYmJLi9UQSMaVQYPzK8g/0OaPNnyTefdvT8Vb0k+B1HpD6WB
JdsGraCbCOoktRf4ygFMS0ENAwoxsZRIuOlxHh05q0bsh1ty+f5C/o6Fyqh1e0QC
i7hfuMcLSaG7sZZQ/J2yO07vySPbxJdMFnZBSv85I7quh+IDYRfvLchQ5567osmM
LJx0sf5gxwbe075gVpwGqnJG2CINGFWDmkEVPHAKFgUBGGfSrtfL1t0c7i+/YoER
P0PC5pdmo0KrzR+jfDdeJM/9vqTHvgU5zC2XKlaYIKn0fHdWGlEKHepuoKoN/5aY
v9rc972DhJyu0DgLvOydlJxi0rCN/CyhVy1Wlj8Z5oE/YE7tVQBSw2F/KOdOy+j1
L9Tywr5nEUVoRTm5TQsHFASipLNYpV6umo1wqw49ii86ww1UMHUXiXJNr7swiDZD
tFqD/3CCT9djbxyu13wNRl3gVg3TCoPFmW6V22RknSbKODSL5/DeOSoG10Y6hwQu
XUzTB+Z1Pil7xQFsTy9SfJG2i7YmctKuN15+T4ZQoCH39DQhmg9Gb9V6jHnagWkW
6qA8/UfDRzVMgZGTJkTH6+JgFTnDkZqM2Kt02ZWzuQ660/YwZCv6/s0sm5p79V35
XUCzXhosFYZDvEksMTDMlXummTU1BNoBPpNG5/jYx2PJ1L7XsgRraaO56bks8wnR
VDCiBHyFfPaeRh5S2c0W0BZqAmi99tFs4yb1+FCnTDrbH3xYcURnVMtVNNq+EqEX
kKCFC94sRQm704yglrlihPBD8RbLS/w+8HewJUNu8DxDUK4y5ZP063QUrrSpvTD+
9UETA9GGCmyR9BwTDMCCOpoMSiYF5KNMffI28qOtoxeFsaGeqznkuTYskPQQ8PYZ
8WtQ/KnZWymp5rP7cP88RxMwfPqBMLQuLJjILYe0Ti7URk5lHRbNG/sVCFDiv/UW
Ui25M3tBKvDRp8LGM1Det4dMMRIOAco11r5zEaj2mQCcW/UAXFBw9IzFKcoTMaed
GmUqVUfZMrDlCYl/rvVls4mmy6luXttOmtgUl/Xgvx+8sxW53TLu+yt7pQ0ThaR7
KFO2O3FQpg57sfOoK/YfFECQ/KbySAgj+ECdxSIhRQS5Hb87eOJSZSquVJR0oHpM
Kvf85j2sU8YfEEmXjFvYb4NiB5WjiFYqLN4q+JO4f9EoD6qNpgHdZuvlrADJpgk9
szeAJCeCtlwuXm16CKms+gRqYiIYjWMo+nHKdkVFVTXf6qYFMsHXRrpSZ8/TSbjx
Yt1rql2CIOD3r0KdwL053gwKPmvzOXQ38tUpl3OtY/RAMK1v1CYKTLl+AY4kgMOQ
WWBL+E5Xx+n1oceKiYE08s7sxGgun9gPX9vAsCtsrxXUvzQhv21qLd5HzFxBNdHu
UM/zjjGyOjHAXTjTAX1D0SwWdyROlhW76QRmI/uYGTMTbjwO/IARz/uF33Wf7KxA
cOtPYslTC1kAI2JUPk3erAxd5R6w+4Vaekkcw45jmG0V2VpWKyVXe7ypW+CsTr20
l4jhq/HfJXHI6q789lrfmN0WkFycnDD6d0v2/TN9OlRezwLapFqLmjBteR1hM5jQ
fla7gMl1s+JIVeAVkiE4fpIhTIlgVjO46hzkU7LnpPWDC3E1uRK7+E/kSpH1W8je
2blN+COqdARZUYVaaMn/v1SXcHLspGueCL3QUPYxTsZGHWUV7H00bjYk8p87WuTT
Qyfv9oINGgHLPsBU9d9pNUjzW9MPZQNNuhR7tMpJo1aLQF0K9qOwmP9OIJqI3U56
NhQdQKOE9NaTOc6ZUBoJRVu7RRM74KrcPRECEN7tUyESWWEu2mN2QG+K7tZpFTnP
QkSkBm3o9YefHApnRwiuap/C3MEC3MW3VPo9fyBbqQL7iHgy/axQ3zS7+AMRV6T3
kLFJJTDocWnl43JvJ8MZz/LiVIfwTOYwry1spr3ShYIKP5SaPG1Lco0YcGkLdyiP
LZCfmBWHz5JiclGYtZu2M/K/0DZP7rhmR0qdAzuAALH2OfeAD2h/5ddqsC+JYQ9e
1EC9Bx1E9hVHtjOGUVSxHI1r1VkutLUcY6JWH77yFf2soAAMC46XMV1sPsHKUbKx
jXxmU3CbNyZ4zjTK3TMJOoPX7SpMqEGe7kFfirSGPpYyMpw/nnM9JrebEsZ9Ims+
Kt+FeYaLjuJAsP+b71GyHO0zHAOWlY63rHAlh9zRlyDuFPFrteP/PGcs95OUTz/A
VoFIFlcFiIppCRys2hDtS8NUvzo6nZEwfiqLpaYkYzFPDUkpKkLA1Bl0WTQVKwkH
W0RYMo+/j5FKwxVxlDxWT8o8i9tqYKEdOR2STFnFyusl8m9u8ZWWn6o3DmseSce/
dsm+tVdiKuRMxtNgZYdk84h7D7HTXvJIekoQRIW2M6KHBrSFssrOW8xp1rnLQhT8
gorJ5Pe33ZeRkwWB/iRfdHOXAEWRl0PIP2FbE3nXWU96iS1DvqV5pwu7hDsIz8+i
qDS2AU4QX0dEDAACluqHA1/SAzaJfq3nCjw8nGp2UVYhUgBIqN+4v9Xnl/KuauiR
uxTUFf+1f4vkJJCJLuOPyjsRD+YbxDinSE+Db1odxGSh4e6nq5A17jOCY4Vyfwyy
XO2Uuti2PYukwG9vpZdWljwDVBXNoSEArfeECBnFLOihv2XLKHl5iyQix17YTgSX
3GEnftwsxsur3tqg1FbCeSGSD3gvvPz8ZPEzma0QILlvsVlVsmj8OXxBcQOfj3Ad
Q9DRhTQjBFyrSj9Ze1vPqNDs5xF7Xduahk+joJU/vjo+e9e5IqxxHO24XUCePVPQ
fGTtc9rudsri7LhSp1uMlpJ/cb0Z7+D6dAcY+kE66cTrcyOqOPa+OQu85+WUBqb1
a1g+bryMLn0pWPs5POAsFb+jx/cipZiKCLIWW5ueL5pKPpR2Q3JQMqj3y6WWVe8T
ZuBdRkqY+Zsp0329vJZKfKYqvRjMoXRGa1/rI4lSSREu8z3eEdnG+loCpRcI2SfZ
9eu1xBHLWQg2JtiWbtKfSMPvk/Ne5Iz19uqbe/HV2iJgeT7oBKDJwPtTujbUNbE/
XOKUckiJ5vNVUiXmgj8r7+LtHrMvION6zSyQ4w7xgwWm0u9Ca+qqjI+5fo8DlLAu
v29hqPwI+Yoe+9PvHjNUpYWiwA0+/09aB2QBTZ0fDh8yi8SxSDY1FB+2OfSKMVwp
jcw/JAqjAx1AiWfRG+Tsa51OsZu1fHxs3/zoOyXyswjNUIF94tfDe6756omQOGvg
zLeX7CXuEo503QaOul738/R48j4PbseaoQtFElhVyNGAOsoN1QZF2lMXUYXOOenT
O/1sYeva0Fw/jSNcc1R4+ZGU9Rou5HJ7CalJGoRa5g89dsN6ApbwRCjG+O/4srux
Ez260HNYT0+npL0zaIYRLoWcNW04nqTClUTiGHpVfgXCCLERjSb6lP/oV3j/AOx9
KHmoEinaq8NwLvPXveVM+MMXvCuk12FI6zi67jtjB9RLSilBC813gzw9sM2d/9pG
FSW/0yH5TB/KIom37h9CyPuEy/opXkOq8J5sE/6uQlYn4dmUUueF0WXsw/nYJ/bi
84UYTaBycP2p/DzxPvRm4g81u0sy0dwputpH1Ui+ZbG6uFgH8inpBqzYzWygIdrn
ianiHxKo3UiLNUKoR8JhnkoL1hKLqv/gjerw0Gnnp8i/XnHS43uuYcJI09wz5qqC
iUf0k31GZ6CWNKe6+WaZyLJF5HDeXlOlJe+B7x1YphJdE19Kqwyumg9EDxDMykb9
QnVnUCNhhrclCI4twaMQIAPOPCSnK004VnA9NFgPErQ7XX2vuo9lX2A0Q0/ygH7Z
QKXPZYMFhCyZF7LaagoV6Sw6NkWkl1zVtQs/td417J/fifInYAGt5MQ1aum7AWE8
Aibt2hUoaPh/lPgSVGbLzUZEqqZhOjq4d4R3cboPps9Zj3Gh9VEdxDR0qd5zLw+a
AlWSTpETh4lEAxnd40vfweXSRFhbLl15GtxdHCR1i7mpoIRzcBurvSuaGcsMwnPb
XZq79GXLLQQk9nEF+pa+KpG04r/eskuBDXc9dSj03Uimoq/pvgujlmcAMs4OIMoK
PkB7ahDt8FBBm/y5XW2YaOiZFzjngx+Mw2pXNIR6tLgUsnCXBvGGzzWJyFa3mRV4
Wiwbi8alI3HpJw2Hw7Cv/0jaO8ph5dxNhA3oQ3I2b4CFeS2DytEKPx3SBONmRxnw
6ezCcBkW634ECzjkkxU/T/IVUY4QZj6f1lMXLU6WxEivBenjMU2BGaO0/41Q5VJh
TFV3WE9KPioirs4XiZcGBWYe6xAcS9vyZoSOnGJidRFwlNduQr7qepXdeU/5zETg
+Cbb5kS8YHTBhqf5aSIjAd/jQe+2YzeKKpaChq19FagrpE3J6HprSZdsOtPAirwB
7ubj3uW6VZ/hMo6kpZuuVlLECb041ndvCYUnWkH8gQIUq9q1wJksL92EgzdI2vM0
+rk7kTHavGS7ijDLxi7s8oTyG/VQL2/SYbWZhXsLIZGMERVEMfzOIsRYgISdTZ9p
6p9Loc2BYv3lueKLGgNR5tEKnLdo4PQ55zv6Np5sIJY3DleSam4RgGZosbHj6BaZ
scWiWwNVxRvKJPdMfzojdoQ7isIjJlc5GIieUS2uwW45ZCDPQXbSoQfjxVgduAQI
O9ewsJbSnvpp7u2vjikkxNk+oyBcR3Cahw7o6jnY9TZEFlX1ZSrT9G19s/NfUR8W
VajGSFEcklKsJJ3WNiigxNCTZ++UKlwGJPAYASVuMYI3tfkccuhBvEIKwbT82QE/
FgnCsfa+sTFdJ2OD8YvIq11RTmdql4tYq27/vrHem8GnPdlL7+TjVsB8iIrZ48xz
QKnSRUoKC9i19tzRK/wVcICJrI2InNzqkPHqwuwXCnqgtGcbTuOJmlmv6zCu/tpu
kuE/EITagjOWU6ToLp66muWAq89wM0JcZIoWF8kCs1etELmEG9RxcvnofUeAmsc0
or1F9P+IfRCxcIXIANtAZNKuV2T/nkGMUht16pCf9ip5X9SLox1Tir84X8eIrvRQ
s0iSRbsDUVTjdyqd0sNPvYRliERip/7QFL8QmfzECyvazZMBdxcApD+4VhCbku1M
JYnIXpxD9uxGhv5GM6KVqVSmfTicPQJFcvZDM7xq4c4kLJArGweP8lVrxqiJT0QS
pm8Uoz2oCTpKrGNW9WjFYHtRz/NC2RHsD5nySXFuyymHNGIdKcB/2SNwMuuvRllV
mBy0EU2wgRh6hTuYy5s0krk5FN1dkpfIC+KiD0xV6P4pJUkKAsZgOZDb5s5HfTwU
25OBFPdaEVSwsp0aAmSIMZ9Fz2NmE8MP6+1BSV9VQrpU5IWuMnRawPX4hP5Yy1Yk
ESQEgV32fpqQrj7lbgeJqOIPASQaNaQ712aZ+lDVIvy6c9plU+k9Zf0FLbwXtUux
9XzvbfTZUOU1GLD8zswMA4x7yv7ao+B7iBawHg6uBMZ1OFD0HiZH9N35xUDzPNgP
LOPc+4Doy3shuCRCod3r/27uyvLwAEIPKFzFhFj2t/UnGGVD+NmZJyXY2AYzrJTx
AfmFh3fJyBmBt2lanajyNTy3BMTvq/Rj86j9V81Cf4TBjj+kIcdYUz5v8r0w4ZCh
Hp8G4X1N6r3JDmLzpuseCgIE5pHmg8b/6A4iCzMsFCKKhLhkj9G6anM7dweyX9Gc
KsdfowUgZwa+iHGVq46VJWz3GUBKkY2t6R7TGqJYKTrqnODX2aFigYz0M6sH5RpJ
wPClSzmK7Us/kjVCSwG61XRwClruQ90JS+YgrYChX1IRmm1p9N/ChgPNYX5XCG+4
kZTuLhD9htAP36u0uWNuj5IWgRBl7QMrcQVEE6EDsgZJ2L6Ic7kj6wDsU62L3Tjv
fplDcBJr/yyfT5gqg3fB5nNnBEwpiOd8zBzMJB1zT0kdDY/VYbAtj7auYzHIc9Jb
S7nCsRIFW1DCpxppdRRJT4wyhjYcDqfnZHGOYiVhrBOv12jj4HpmUPNhp62zxbB6
MXf0cHQcqYDiVZQj0wT/4yF9jIsS3sJEoLQMN9KB7xfxDJ3vyngVn/qe41cVW4yf
HJXNSajn3xbfTTiUuE2qAjL4ayOw5KjnfWyTHb3xb1SqTPSD3cZa+F0RTuz4aG/K
2R5Wi+zHgB+YtcThZRx/P8LStXgXSXP2W5pOyk5ZHdEWTkPMDdXBkYa191ncMhLn
YjNzaxgPgss025n99lR3mnv71f/vIWLobTAQFjZy94owLj3ce/Y/2DS3Z13680zV
T0e68WI/doYqxOWY9tn0GXNaQrzTGVX+TFiV2iE/89qnG0N6N/GZj7xqP7/AMSfx
LDtRkSf/grLjCvNvH+CPLRgyMZyeG2QA7qAuEnwBlcel/2V+PreS2aG+wNRBxi42
BactnySKox5S+UCmQc5y0dhSvqIUvUnXFUGh+IUy53K03CkXAEILPJfO2HGZeLyX
70SlHSen3S0gieRN7l85H3GQsY6LSMthnh4Ci48T4pk5bYqlzOK6dj6hZYkl/rMx
/WES/autO40YMReyP/3NVoVDKgswDlm7CrWsij/tJJ7+x2BoB24z9KYel5IzbQc/
kxpMubpdobREivdHWhOSFsPAQloNsMYHyW4J4PI1VnB0ZhCQCSDAmSfppBQ9CkqK
J+02nlCZvswJPsIlQ2MYjSILCAnUVywQmRlY/FTyPwWrCExz3/QIAZw7gYSqMRXc
iVuERLSD6wEI4L5fyx6wPplR9lpzRjz+xlWqTDN/zvQsRT79NHOKRVAql1o04XnV
Duba7JSepppI0VPmmjGAMhsaIBMkVICw9C5P28cMW3kL4H/LWGxlQUztvlLxaHZ3
c+RL0trcxDUoK4qM5HyXtz0UL7CBoqEYpEcf4ceV8yUE76MzuvJXxlslaTwbiCQb
mzWfC5j8WBxohQb9r0hcf8RcknxabAoAuh7dTdzYoyeG36PVlqUP3/7Sh8bxytk0
nIDnEyDXhXY9a8qrMC+YbwpxzreCwGpXT28xSh0lHRg/9Z7Navx0AxGab2CFX8cU
IdkfGe0siNfdeZPa4LDJTRjRFK6f6xLXkPEN4VXr0vtMLt6czSQQx/lYTGkiSfdU
qfKPGxdudJYzB9V05f1ZNzJET+/tb5OWWEXSXWWbswRq18GeHRtJdcHaxXnVi79d
11YRJFNd7AXwnM0eLCsQKI+z+9R03zFyADyPkX7D/f7mbBOMO3+/rOIy5vrOKZG6
y87HKbpliMlW2S43nKKYDQvw8M048HC0eKy90GPOZmX0TAYCzYOMASmwhQCOxCyS
jjsE39WifUmsD2yFwqnzeiF9NJPKRfL3MBrikhItGRhgmBfmrnMf/XcvYQ3VKm5u
4De+c+uExhPyUX+0smDiXRZXGJB3dhSHa3TKw3K7y9/5R99Ytick8+Wt06GbsAri
Jl3nKzyk1eorXBFZIRO3AJESL3wZgqHaGHxtQ1kS+N7oyGqkzUMP0o87q4m1llrA
Mp25bKRz3bKH5pDWmDhuFRIdmokOATu+wXY65+7BwCFm2ixmFNrN9Udd1pff7JBk
ZOAl0nT7f6ad1YgAvEa++7v6z4Q9AmcLj5Je/mnafRLMNhicQ8WRkJf4bAeSzTk8
wGmaK/73NVY8OU3fr/DVdgQw1k+S6nVvRfkkxlt/AcPAb86WXGpWpXsFkYEQqpxH
dR7Nkufo9uo/IzT5V3Ecza+GgeFXH3Wz8o+UTTpHiyKZWatD09WVjqYdcN+LgKIb
VsFwNAmpg998V8ARfCuHU6/EiHaB/mbUw5FvhPLWtskZESJe28tBpBZPqxi9Gnkg
Xbb2MGaNVTpVKrgjgq1WUc4G8IaPhu2d5mepUOvZOhYOJDnoxdGsmaXX94jZiHBw
evYbW4woOwl6zjxPxey4brvsLgWc4R9Hsz+5+UMb/PHSBC2VWruObEMCh/P9tFdm
Iy+y9wJoqU3FBKW6bPswuNW2EI315kx1BBK75Gz25lS6Cg33Ch+6M7Fqeb5wC2C0
VGLnFIT9KiMDrmGgITdm69GKybMpfweCI5KaYBsHC7RMWr3xjl5YTjv2PXz27VOn
+6O0rd+nC9h/vrourhbscaly8T+8hcVMBMmGOsDxYzSb+4C84Q7UX0tHignAwi8L
R30xkXL3fMthwrva+RLxpZwS4nW4TVKR8BbzFvYCdG7Sz7eYA0Fj1zc/FlhnGgHa
QeHVsKJprlnXjT7UA4DQ680AzkuIiJ3P6VZf2LScEI0DdzHgmiOt+5tUjSvL1aNP
vfcZtxLTIZsfOD6gRWeoVZyuZaS1bJQJuk8oom1TJkbkfsSuLwE/WJxLAif/X+55
fR6w/mnLlhissGXuJGM8zK64OiCY248A9QlmggMn021p/D3GpatIJcgdCFf7NLTT
AZVk+khaE5W718KX4wArH9CEcCIl3JEh96GxZfvMmTrcLEQYi1Bo2tc8Nmdz3xzR
fSIHi1F0CVma73jmTAZUE/C9kzDwSgfxzlU7gWTw3OKzQLry1HU0xs3WvQdbaVM0
/ZR2mCoVctyHUyjQwS2qo3QYQDZh1oap8dl37QZB7Y5bImaejoOphK+OE3A4Z3ON
weQA8/TcvYi7tTxCj1xHkL+5PSamS3M7WvUc6ZVaIEHkXTCnOOMxegtw3e8HpL1y
NqGaQGHLHjmnquEkfAUvO7f8Ofme0ziIgeKWJWW3W7igy5N9K4+RWpwZs0PRtqK2
YgJ5KyFvoFHZATiyy/f/q7kJ+wcYRMrdZOP0kEGPsisR2D/cBpcu9hQVWVrv2PpH
JMDHnjoIdr/OdAcUSDxjFEkLblc7QGMsbWYKNcMUxtTjGAqeJpKWNfCgA+It9K2h
9gCaLBxDYhTi3OHqiwauXtsh8DEhSor6D/HJU47zUm0HLGRX7KKzVKFnmkB1Eulv
PyidG9+WyrkdOVXzsZE08KMMImPxclhpXsbNbP8CxiBm9GaopU98OoVGsSGwTqER
HuW4G0OuIVEfAJTOrSWTtA0Z+DAoCwG1/6HTodBFhM/5FY5B8fFxUysRC4Ij2eM3
r45RB9yQWJ6XyNaSu0muh/BH6vU0P3ddDLcgnZHxA9pc8e0XpIpos/f4toC3yp+a
7uXlZ83eQpJDzZoLg/TVT92N7AiFVkJEsDWJCc8W5XqLOyl4gFMC+t5RvlmA8GlV
651IWYl1Ogcve944CFPA6Nd+7AIki/6vCCdgS3z7KPStJapjI9E+STAK+xDA5sNC
lHM9OkkSbqv0V156WRRslwAMaN80kDbEyUVlYMVq7NeHzhrhVT4IABo74bYdfHYp
3F6qcmTINWXo8f1oj2n5sK+yZkm3NfKhkib75g7QA5fZFR8xP4AfrwLR26kHvN2s
IuEXO+tCZSnk49yrHTT7g9vzO55gq/bCv6EiZsj0nKvEUaZ+sxFRFAQhrqjWeRJL
m3BCALj09iZKcs/rn6hxxh6bdlu6wh81pCk7TNpMvL4xB46Pd3vmJjz6Xxg3VT+1
P+56APc1a5KaVx4mPefxYgylxpH/Tl88B1tmJxoWMgs+kzZ0PAgvyd0WGtGIv8oU
ETP9T0UrYFRIEqFUDli8RhGw9yZVdOtSkbgznTnpKjpyuRPj70D+qaXiif09Eekf
K1tFHROHtUsqPEFvOVY2L6Z6AbN1RRrHr3Oj+w+tVXghph2zs4fOSQqhng9/aC1E
cTDRpfSQfUiDzPeWRyTzOwhK8t3HRZx+Nev7TSas8yGM2Tx+lg+Mcjw9hT0sB8rX
8lnBk2cY/9rNtKVb6Qo3uvwn2XHQPpvkktPXvypcBPAbh6zSsF1toBzxtK1UK4SG
h9tSFEeCeEjqIqAFbBHvWj6J2JYE0JEsck8FVbqrdseApu9E9bABQRa7OAsumR7S
orKjkYJ+26+M+6tf2vUbxIaz516NPVXhmKs5IZ5PO5GlqR+bwJXqaIlbUeGqPx/r
9p6xyK88sAkQfTfbWk4LPloHYwVHtubaKIGCwe7HhWlZCUZXMq7DaMBnR2OEyWCL
SBI7H+0efHoCYnzeLOOr1xxwZm3cZ2uJg8dRwniq7H9c8sxPexOCKmLzWHbzzSw2
x0PjUja/hs55FSlwBnZ/czwM/X92YmB0PV5tAIljT4jcIlQluLL+RqKuyT6HLLLL
zMcbBjTBZEbRVTBK9B8fIfrXEUkHszGDBi3ZqvrSQOJLI3znQUIqr2hEPWwJyoFl
LvUXkxTskF6RK6ProVmD3Ziingc7O5R7TnpdwEV/aktsTCog2MYE3lnRGUCB3Pvu
+ZjPb4W5Bo5W6e9TgZK7a/6i40zagzVa0Op0CvAcSjeimUo7zgtpMJOJ+dgAKdNR
Ykgpnp0GmX3fII9Xl/NEsHsD0VRSzdFkMH5qfFzMPT67DY8HSJO11+5hhjU/zdUz
XRQrk3eG7DJzlN8j78N6cSGBRg95n+ZsGXC7H9Zy28lmsU+YPHoUu2wOnDVIItpC
J3mbNOHM6/FsIE7u51DBiiFefl0022EIIYhKsbBK9QXFty0Je0GpUgMlGzGXgaZM
28ApIcuHfQtMS9JoAETLxPYZqAgI2Pmp53ukRFaqLXQXgG9zhWt4JyuKu8AkNxgr
ynw+wOlbDb2HVQVRDJJrRs/AdHfoVxTaA8lRaQtufUMXkLdDE/Pbp/FJXXc1WAsc
i6mJ3lPrBBM/ai0mXDupnrmRGBhFpgwYq8amiUsRtQ2Ho/RZKJYMFD9uHqN/sKwD
EQDVxPk7IssgT2Ds3DnOltIvl6ovuomiIQziiFRjb6XuoB/MwgP70bV7eUzp2K/V
g4ZFWr95T/8cwsBacrWc/0QtVOQId5IbUrF5yIQJbyNXDCz010EMx2KXKLwnh8Ii
bpcjkavVdn23IYzIwWK4oEWOVi9uuc8eDm7dP449jeyGReKjTgRUo4MhjYJpM2Jq
E3NbXQ+sbFJVEQ8rrhM9oi0Jot0NoALFPS05jl3jo9QrYAQTXTYU12kozJlZ5CWf
KmdE39Zb9Z8w9Grlm4lNp+nJDn0+S7MQYFN/6XZvUIzrg60o6FbVJheAVpv3hnRr
75PanGiDC5Tnd+ITPkiQ7DSd7/QXxLe5AsMAS71S3zKE1C9dAsr1FWQY3VqajkaA
PZMyQzIpD++RXfXpNBQFlAlzfaxA33k6eogYHzwr4b2K2g9PqQ8iwhEk2oKjlSvn
vQ1gB49Qkmkv+SHk2HiTvlWzhZNw74GYE8NlBmRigo7wsM26wYEWavjbvGLYdJRM
tnljwmgpiuD99uKY+zLs85GfC0DoVTR7yV4Iq+NwD6miex3ue6SjIOy4NDxA/N3H
NBjP9bRQGF3TUFn+J3C/N3H7Cthhx7ze7HTBNM1fXOv6Fto5Knk49Fd7pOQoiUiQ
SMqkTlvF88BGaARtjLnA56P6MvW1MvJhELcnFp0lX6eMY0EYKGZhH0bSdiJ2+oq5
dHzePx8ovL3KrBmV9tP/7GhUNYjTUh6w7yIGyb/R+8CQCG3P8pzu0RNI/Q+9lS3d
ND+dHCKfSIOUDfkLg7wozIKTZ/stz7kIR8HniDWy5olJi5iiLnvv452kOcK355iX
N7dGqN4WPP5FEf51rOyfmJwNr1JrAhL5jOUU5gtBV7z/F/xUVQgQsLntDc3grBAb
1LYi19CAcp3PFwOsEEOEuU5CNFum//R+pPUMjSB+jjsmX1h4cELcJV40zmKAxHBM
JJazPvdF+oBQseAUL3V6BfibgehS5dpGG10BS0nZmiGch2fi0SuHdNzt/qAWP0O3
HgCITcsZajZulv7bMsqsyzKzcig3wtgxACCdIDo0YaQDk3lvKK7Z7FS8N6FKjZPB
xYdfXV5hQZ8ISlz7YilLvKJbbHxL1Yd++5vfFt5cjWbQBLLiKbqnBZ3XqXykxP8G
S65QLpOwyB6nk+YOWyiNi9PXo7OwjDd+6KzPk11m67VcMd7c84mxsWfbUGR5xRVz
A5fmO4RzEZI4pArSpg43ytMCPp/Ken4S2FNoMasoTVtXsVbiy4nzfF9vDV6OmfSZ
lq2IfGlaWwkKan+cOIFdUOGyYCLxSbHh9mfnfnSQKFjjlf8TZ9D8AsHlRvYd8xtY
OuzqYXE5UlOmoMoLY5zOgDyY5D24nvoxGk3cVFN4ihmjlK841/88FS6bXIOBG8Oc
U+6hNOMY5kWR7BN2BSnppQ5thwEzjrp2qJp0oFpluiBcu6/5/b/neyxTFM5MtISP
tWrj1wNZbsJdYUG3z9Gzj3Yp/y8dcIl6lnHsiYv8vRfNiXYlAiAhv/C64Pv06Bfd
mbkr+nlDx8whsfncKLoMgTk8N2aWBKL6e5TdGyWTOixeWbwreCje6rBopuu183eX
6qXYqJhX/4eYEUzvi2xA7hRcW9u1/OTFKyjuvxSZx5Ia2y3sF8xxrpBDS8VBEqnm
9dxf86K/VAqPOUiK6ePEafbu1mOEw4YgootlwF3z9JVJnB4s0TWgyn+ES25OrMU+
QmzzJyCy4ldxRqUncYwZswx/MlTGeg1P8j8tJTNsJ6sb9H3u9qUs9R6J/MgCeNV7
hg61AKTLBePlCTFf1gJ8bTMY3b9PwYlcaQWQsOVHpzaMMDxUmK3gsi3IEqK4LvSq
DcIKcMC5IzxurjPm80GrNUUoFu9GYvcVK8oEEwSlFPYnRmrzqa7a9PCnVwfitrIQ
eoRE4y8dw910nmWt1l6avxSL6CB6fc2G1lxTB1NfvneKf+0SnkegC+lhfWwIpaHO
w5+OgvOVfmtsriDdfIxhE1TI2tXh2zcTuJF6sFhlJ8D5YEXjFgNStGS/na4Jg4P9
+Zph5eumBTXky2GBqOWCRCI/tIkQkdp5uWP/gZ2rD8XA8ffKzYUtvWkpgc8SclNT
B7ZvyqXRu3IUzPeZyBqQk1CFnfQCVwMSp6XFff9w4zeP0088N83u04k/hbmoGFFA
grmIqGXhmmAjZWP3LMZx+p3a5xLs1HLp3r0p7m3cdiuLBcTrP0L0Daqn2TE21WK3
pO0JLMLrkIvr7/5tW9H16uVkLCah1iYeZMvUuolgQqX7FgJA89Mowy6o5BEo2R5o
3GfNzSUZNvTdJ/YCL9IiHNn94LYMQSpExsYbpeJYpELtA8dXChoEw8le2rAZ+REf
FjZNRhYWp/7TQ6GDTr6p4vqlGdUc4ceplhkXjlnKcfQ+g5lCRhTQ3pjmozk4npvO
wd3jG7peS3GGPcRFuxhkIul5A2JX+dvdGbHcpgWG9X5WVuWiyY8jbQPbDg3em+pe
PVMSGL8OrwUIRwoz4PUrhhoE6o2qUr404VnQcahR+N8CqGIYueKlWY6IYTl4vfCF
uxXH2VAOk8m8sfDCXo9GazDV5xDZuYT6wQYBzjoP9PM/DqBxAHmpRNIMmCeqrmwh
eLi8t52lwsI3wKZGYOGgnXTEU9HU7YnhAtoAaZ70Cm4lPQYl3+37qoWIQsB6I0Jo
XNfHJ0EByeuipdA6nHZiR/+WfrHBp2CkdETVgykJwPISlj0+xDszjfK5VDS6Oq+q
Tt+iRYZLDYjuP555G4TyHMo6oPJor3qWSnhtxHu5B7jY11Szjmv962corvFy6A/r
Z1z3DTpaVSOaChcuS63kmtcIkDKXEKY+9HY3IcEpK8N/pK+xmjzk1ys8+KR3Wj0U
fvlzbaztz5rLbvLS4ecrSv6it4zR1stjp8Ki3tcmZo7J5nWREgXGnp6G/yZErwk6
J+P2tgvGGe+OrmaZm2IgX9yx7WMURI/DUgPYbpqx3p49YdFGDJpSSCkB5KlCxAY6
onBSScBPHsJqwCgjuu2C4Py/Zd1K6JHEYrSpfl4ViYpkOx3zH0d+zI/Xq5ex5Uax
YhCSaS2WuPyskJGcLkDBDdgoetvWMx2+lPsNQIPYnUx9Y+wic45s/H0hA4P1sc+K
yC7duWgnpRnvm9Pp1ZUWhCM1g4oMgJVgqdAjKRrjxOu85eJoEsCToCLnUyyXzv1s
UlkDhdnWSzJuM3UA0+0Gfw/pHe2XakhUHuMyG1UdXsdXWsBkvF3cE54TZJWVv1xU
EWHGAm8+mLWaUrHap+aVFcVSfVZ/uZWDwSEFBe/+vkE74RuKKRzx5XOIH6Im6e5o
eogZlxWNhKZlFa7/yRfsadf0X1rZF53WL42P4Vhjk+YWAAR3XVTeo8r4akEL60jM
HmOKNdli9/2fmEyMQFxezLD1ua1vFX8D+kn/3MgwhRPBfF5N76dQM2nBHvmil42l
fDsItmpLGANbMqTwh2NzpDBjBIFcRQEHnX73YtYw8fp/6V3usFlDNND23yHpf9lv
Mf17+ZDH2KuQ86B7Ymd64Lz18XuS+XaiOn5oi9YCq6qOGaicnifepQ3oPe7v7S4F
SDTW9LE7T+jdJC2EdEsqtCebmmlwM8IiRXL3kWeJW2w2NYfy0fMPC5dyJxQIABc5
rApV16bgwHvw+h9HgfoHCDhzG/u/c99+Szy0FQ2SMpz9jIIVHY92kezygP2RTmKZ
3xeqM+sWaf7HeJoR+HKG+Ts7ilf4RDqaTy6EL6LEDbExPxlIogrmYW396l5WBH8r
cHF3+O04BMLo0yfbzLdYBtnHHOon1HPj3fXlk3ex30frPGU3igywUFetJX4CKQN8
wG1jVqZOrTU7MKBKDwhEwNryiE6QL5w3j+gsTygPFd7HjfS7caHtc3/DmwZu8f2v
ELbV8C9U5Un8pyX0SFy4lMUFbFlpzbLxGIQiEOaGOzrbYnORJA5EkZRvb19sgd7A
ZycyJrjhpnniirS/0IhtpywaEIIZFSLq8ci8ktSfhJVzNoHGzXk5H6ABtaM5MZIC
Q6EZh8DDSpi3K3DO/otME2WTXF75Cgx3WTJKxhoReczZYCZIfVO9vgC5RRG0ktGi
LYUkhIgsY9B+dFeVzy/R/PxwYLZzd4MRxsCBcB2jiNdrCLbiJrWg12YzGgqDFh4y
+BUdNOfD1POTe9rL3RbBwyK4BfihXD8drkY2Jok0bILnE2qwfoMdnDaE+N7VbzKM
HoSRbUPcqUIYbXGjjIcDK0K2R/Qzf8NTNGfRqG9maL70x0ooDz6QwDJtVf+Gj7qr
jxVFLqfOYyX71eNR1+SieKh/Al0NG66hPhOVi3YDfuMJz/zv/iRhY7xVne9p80wq
w8Put4KtpgAOnK438IB9YVtmkMdJbLkvnKPJS9kLXj9xMO7ldYKKDWDDn9oi1XXC
kLlbBjmL0Dza/2tYysamDWovOM7NGPrOXRqRSLcIjDpKadnrJc6aqe+gjhtnqix2
KzCmnqFElw7Bsi12Kt8BMyK7fV5FViuk9imWu2CsTtHKDjzNlBQzt0dB8Xoo9Asr
xe+jc/R/lkZfDbENRE+3YQIxe7sG+/iTSZeXad/9GWuaTa/z1U50clHmxsOkjn74
82RQItMEOXA91eaHdCMhQOJTZIjNIwQldDNutTbwI+p7L9k2L0oW60Xl0O7R2T9K
/FLB93p4jLT9521bH6NDkzsZ+GU/TJjRbXWziAfAAeMO5V0Qao874FkwyTm7px/s
RVUOYd2P2JhQIUge+vuvtflEaxBaafo2/iJXLU2CaZbUMiIwrdnYmtlcXfHIeUV0
qycKTibFu7waS8VL+afqvPbcSoYfc0ML/k602xhhgkJY0qC3Zng48DDUk0scogNi
fHFjyN8RG1PkNGRgmWPhQYTzYFUzQE6WIdT0+6x7I/sxJhrmp43uwWxtEPFA7o5n
vHQQx2pzs/up9A75XJ71wW2uKHL2yBwo1tS9tE2EDLOGkYdFg4AOQ8wu5UV0Pb1A
OwCJTuOyMMk01CC7rujAq3VujM+CYJjMDYwWdHvEu3F+MnEAVQdU/Is0KWNGdJVv
CEj9YJHhw0ANBsuF29pPMcxtlHw3+WlpMlnR+ft/VhhUcmt4zSuNV/Hax8qey0yR
K3X4RCKYLvuGmNAbSHnMiovHIJ+Vridz2EULO2x79RiCvuOWGP2Ha6LGTEDgaBL8
yRkBk5sUowfImT0JbZa3hRKZtqvqc/E3ZwKwc4pMEp6tGnoS5JfmSTejPmYsori7
+36ZWjwGGmmo/vTYt44cJhCdpjsBPAXvZEW0wFvSs7grsTAiev11zMdqhKrsoCvC
RTgnkAUxGYptHyaojl8nYNy9bvN+W0WCtc1KsOmm71BNTOjQ7285XmZF/lNkgCFb
lBjQRu/omOm+GXtyIDicxCOIHfrOMriHJSndijdyomSHuaFP9n0HWT1kJpUYDDqH
WTmSF/AkloD2HaT+RJLmq+3sa8wKnFfQG3p8a9FvXqW5k98UQ2WlylsTwPFvnp8x
s5uRUFI66UvD/NAxgQDZPDBvPL6gYOgWcpImoLdcdU7xLBIkE+g/Lrq4/MO4GLZK
ri/DcLajrHzSCCv5F0g5DaNw/aUm8ABAnJr7415Lx2khwCAUyge+Tt4HJqOa+ZpO
l3pldyzpNaPL81k9rFzDPlR80E43LFENBPeZ2bqedwP9btKwakSPbV71NEINH+S9
gpxPoyHMB6uQFyT+TO0QRU/Fzt7trxfOZ/UqD2EugVisY2jyz4fhYbruNSMyG/Cf
WTzz5ccDY9+N9RRxpLOY8vpFiPAiAJDfCTurq88MqYrbRtuCA64YB5FT+U+wVu2i
2o/acVyYnm1f9ToIgRDbzVBwLZb912K/2mDTjzGWbTqfiJ8KUaP3LPfPy1f8OSKY
dU2LY+PeUWO/c1xN+bPp0jRLOOVrWxkz6oWufAjbsPzY0TAZZwaVQYetFuffvQkg
tpv1HwXU3qLj0nECRjjkXDhJD9Mi3NmxmiNDdmeFmP/gIxIcSfeRvTU6AVX/pVcO
VCOFP2xBmCvh5+58ofcXi9q/WSmJNUy25AXjS3okVhR3NaVDrbIPJGWxhJl90D8Y
WRvudlRHFcdwOaj6iVtiJoEjqNvwxcuElrWPAj3nLkGTtXe7Y6StAKMedQupsP+S
yMga5rAvbLga1x9zD6GbS07MDghmX0DOjN+u+cuWa9eZdrW9kuJQJBZBuIcRE+66
APifOiC532O3pAKDLxJKlEM93U1byKd03saRsweatIjvPd/Qd3TStLNxySnuhqMK
g/Jk9Eetyc2cnvWtlR5gmjNG6ZHifrNf/s3de21PRD7hzsm50LDt1kKpRxgmX5ib
PSp4PMbFxnLSqdIKULbp/FI2upA2qFawhGkz7S7bF7RoO2D+J9I8InpPWkjFs+Hg
EsleiIiM9KStIXWS4YaBdUrbKecnC94AY1QPpDiG5jzdKfkbD8RcriL7AKGdS68Z
eUgdZglNWp2SyH+tbXFC8IHrsfA0Ht16AEAhHEW5gG4kKkjQvTrMrXvjEH4ogi+L
rwksSQOwAL0t5enxS00japhEZJ8dhHWlXBifgM1uEFsI6WeSU5HMc88qeQK+eVbx
UtbAOSjbqDfqXzoZGaNnLHn2Y/oeo6uzB6sGNJjlNY+nB8I8vRFaRJ0gG3h+zViT
0B2Evz8Vi7LPLOecWytnK6N87ZJYvwD5U1WoqBQqKm1lb6zGNydas0lNW/M5inpC
TLIbw1gtKyxsrZliRxxk/+8Bi9qgPbV6PO544x5df//YpasuAZKPYWViUwGvWxTN
mbad1NKebzaju4U7BgsLBu8gzqmANGwn5swYJ7QCDwKoGWeK/rW8INI0B08TZ+wC
mwlDRi+tJFJGHkorUaytqAtBv4od+Ehr36IelWhsZFvJrlURBlFv/64urQjF4mka
kGrRkQMKNHoqQb5Us045Rh9gaoNIJyYeVJmEt/V0OTdmNzeVJEL8EL3VvM4ijNvo
haABtG0wNRksZC1emXwKDYEZqUi9fg3or/LnD77/wcyiowwuzkS8LrFWsCISLSRV
OpvhoP7EHrVYI/FPE7o4ddWpmdVxhpL2sbqb+5qAMFRORBrWe7u9xqzgwLy7xd7J
lobUC3jxjDnT2uutycx5p0yBB27uXLMCQ1r33gKucjWw317+sexxfFxZuZjNo6Z4
SUDi0rew30ZgyhgiRignWlFAGLkIL/DQoxAyXHZCZirYOOLsicgk90LAq64nfRgQ
QS0ofGzi7oriz+QPXfHpEMlWwyhEZG0VlMFsbq8BeAazxa1QuDTdqSUrk49pSMkw
+K9aL25WX/mf8CWvTl1ijmRwNGIbeHBP32pUjVUh4VfFhrKCKnBaSMZW2jDWahjD
RGrpEn5rVFIfePwUMxURr8jDlrlq2R2JiDUzCvCYcTKA7cReTfT2sXs5JswadZtX
AEuSEknWVIAGuc8T5nN57L7ReJF1I1tUAFG95pCDi+BtqTKUdwtJEFOQMZaqcI1s
7xIj3dJz9BG0Gh64l6QIPnfapyZgVzFKPb13Rfav+pfCA9cHKSPKP5MDcZ015UrI
UlDLY9l0d0eLQVGaz17gNd/kU0d1ukPhZsTeHCN5gUW+Pj2VvYwcQHUVqQw7ryKb
UkBsB4zc0sjSLRxuc49bM1m4EAFJLdBtHBWrcCds2ixQEncVO9TFDk/iFDKnApzH
yS4NJZ1zMsNDXtowYPc/D9/jfWKTw9Tu5DIFJVezkIgZX1+NmQ4RsQT/gHyja9rM
kjGDE5qmxRc5ED3SkF0aEN4KyTpXOmDg2VhQ1dgoyGoGoZ5gGapXx8BZ5YQSWyif
FEuSqBzgNcF+Hj9L/PPOoOgpLYzKxhlwzAEB3YWW2C/F+vUutL/TeH/2bT+JI8Tz
opeg6c8KfN63l/z9m0JVOB6qEPJmMIH3kUYtkXpZttvQ639QclABCoJMU3FW5nCk
/Bl4wy+BZwUXyllTePq53t2KnncXylpz1c217XRB9k0TBVRHNRKBJS18v8HZcV/J
sRRuVwLg4fOvmFNePyAS82b0TLA53K1KkeBUC25reZZwt+UVMPkHgnfsT/gMePkr
dmNO1wMcOwGEwj0JcnS3/uytfrvEzybZejIi1rbXiWemgo9Zl23Sd7tp6g/7XKAa
sMBL6uHYeXP0owM+hVwYNR/n7Yj2s6XGT5a1QkAKiqJ5so1qlEw8GH5UMDEiJjyQ
sLdYeZe9uZhd/ldHBBUh7mXHoNsodXdX35bjWuMC9Kdyo+ddSqrpJy202HRr11DW
272BnGIdNN8vfom/5P+Oh6HYlntM8kEn5FYrcPMyyl0PHeUJhd7HZfFgtf3idrcg
8UVrU1n2LhQHzksOJZ+8pxoNSFU+3VozRNQYX1yrKI6mHDTzYzkChK0p74VZp5wd
B3bbeymYO/9d2PsCqbT5uZBJ9baqL0l/TPpqP7tzo01e3Uwy3hrTaxk2DMQISnpY
ebHerghwu2zPKdjcNu5aeaOTy4m9O09MlELIvJY9SeLW7SKuMcrXVqycArYXPXcI
vhO6l4P/Fho7jqB2IbiE4eBWLZ+lMWb0E5je094wI9Ea3lYCPSwh7fWuFSokfkgn
JngI9JFfbcxVlWVfdNOWi+iaQiQFf1nPL8TFPib7OfqMSvvzrq1XiAw/MADVUe9l
WcWeC2VEEV/OXLqlqJFOvnMRUjXB6wAAew6ksF3weN0vtiGYyGnRco6GnUL0GqkZ
IoZ6d3Q9jTGvYvidZ7lFzdfFBzPzsCT+mBPM5UfRljRE2Sz26jGDW2dq98NZJl79
YqL+8bJmsvEczgu6O4xMoaQBn5kUfazjNZGuGFAlKmeZiioPCVz06LdMe2i/QSij
KgDbMcjN76KJislPkVJhR703cx+YCLZ4ZpubsFJ9gB9AunnxrJEF7T2UMZSLxa62
Lu74Kkxp2ercsEa0UHYEvb99hfsnSLGgOonVwn9pXJ8UW9VWZP4UyUSfZJZeDHlD
9mv5m68wq4mhxlGw2UJBrftQ83p4BbhGKQntlJLzaMAvxB9rQT04aR8VfP3Q+N/4
Q3WXj9hCttc8k6q3t1NhfTrTS4a/mojH3R0mshqby92fK9Dr2Ij/G4ZYt1T+tIGU
1a7s1iMta7IJ5WrgsqZUEUPyRgUuiW+QvP3IPodIzHcGRAvdm5MT/KLntj8nXp0k
AgMSJQJ3qPdhdud9Q26RCFdxkzwILQJklTGEXWT65TIznF/dUMYI0OUk8u3mS/BT
CKMCu67lN19YBf/V5SEcTbIJFcct0ZwyOneE9dG4NZaQ9WXUZSf8TYszEX1o4FCA
IhSMM8YhvPldn/jhCM56Te+hgoZXwMJH7sCLzq9ZpnAApB5P0IXUwHYJyHRO9pPQ
H2liyhiNJkF+YFEEk3TtzHa6snxH/QlSkbXzWCbLc2zHKRUoYhey53DoT1oPl8bu
Dno/yCAG2Nb14PMVCTeMOSGzBmp+ldrlGV4MtV72Zc9UzUR9MbL8rojE3slYkLGC
+NpEJgKcftbNnskya807hkX2gu8A73imh51+TFQ7PeIuKIwfVRRQ2UUtH24yJdpa
yp7XxWb6c3RDkOLprJ2t/BEnCHTyedseZSXevc06v9zz7wuGUWi4g2xWecodZgqp
g7TOSzEf59/CWT1XTe1fQ9mIOMCOHZZf+t3CQ7ukpR80pelP8t07115TJVLh7FO9
IO5nea3gz7wrhNNmcjZN1wYLEqETBP4rNtAwMJBMnfdidBxiqIoXc4So2DRCdc6J
nFw+h5ACGr8i7VdDu8SGvmmC8UHgxSR1xDtUL3mDAggkhjeemEQZltHbJMC6wPNZ
TR6IS/tDXzUEr/V5ekJ3jFFBGHKjb+QWM3XXPK/tNXzzEVi499VBszrfGV1enjtb
kMaLIf4B+f9AkR8z25yUdH1YNNGr3tzDF/BQbSwgUGPFAxq8QSQo8X6YeOc9o7ie
xd6YRVHXa10mhkUc9hZQOyZv79MN7BgnNir5iYOSVPhmZV52ZG989KcDfFuLGmeX
vJ/sEqrrYUg1yTaTIHVYo4t2oYhIHdCYdHr2MV9P+uG6AXVhiJ1SRLMTeKSiYgsU
2XcgVd2D5699pLb/NiB80FBJ9VHyRqcwT+O25IHfm5RG9JK+NuVxf2ufmg2jgcQn
ryUMmigG7vxyg1WBLwKrQYENsLHhTo+N76NKl3G5YQUtgeltZvMVLx/2wl6zR1Ic
5vsqvnMMGIMreCEAD9p8mYUda0lDyxRTfC1JMbVKOiM1mQvJp+CwCVJMhrbAqeNZ
yNaFOvkQIGwS8pR3DPN3jXzaYgWnZ3lPVgfXJ0zvKYdwBOQjoJ69Vk4N6xh+eHhl
tbsBJHBVhIUNTuvwekpUkxlXVk2PldmfdJWSHcRVwomYqubeEduuGbOSym8tmGl4
oSLSu4cs1meQHveTZ+/6s2PWaR4GEwcVn0Kr70y2BK1FqufNgF7rTQfvR5tYlDOz
1gz/kCzpQR4w/NdjUYIAkQbZT5E5XIKjsSHVf64J+fnmbCofn45AhBa5wRgATSg2
yxephDm9VkceCcgTCZyo3wB+vsyUwAxb6u+TNQ3mKyBaWmSWGwRmO8WgQ8+4anSm
T8QP/HcT2XHBymjMh46GiQuan4uwQQj9wRDj4MOgekGhNE3qp75yBP6/pt6z9amu
KJKjXlLKxcHgSUvCr5gxK7NOTA7DPfAREL8ddoESbWSBFBRtNFv2gtiiil752dwq
65U2sJ96il4+BASa8K+jDH2JKlcI+jLkKACldSbvZ0I89yUcY5qpqr29SdD2LSss
kp4e+derbiKdM4ls8Va2Rnv3wznQq2Loi4XVdVPper4a8G9fwKmHiuY4R97lljc+
yfhfBWQLpUoOhb9RHPKU3WrdCXgskyOcD5/jneFFcZG1WbK7WT5dQB0nXD7ioky/
8JMiytUNBfySPnjb5iFJHa/FD2QqeUr4WfY9MBJ0+ZBBed0YCAIHxqKqBx4uNhMG
od4umWqWK85fcgrO4bASROTQ6n1VUuWzMfheyR0ZXsxgivYmo2x1+WokaQcpdRkl
Lqh3Yil7nh8X8NygIxDXB6ddmxFtlhsLJxxjF3GpoIrEkcHLfBdd437xARgrHz2F
hvOqaN4Q6SSzm0A7oH9VQkOyFVexdCTUQ3EQ8qk3MSz8k+fCgCUc5LkbpG+RMwDJ
yAZNWbwjL/11prXa8+2omqKcVbexEa15xcR8kGPhxh3V/fOC9XkNU01ZYcwRo+f8
s1onRhb/Qckvk0EgesVO0RvFkUjN4xF4/Q/qoVHYqssV1wZjfytVlMfKg2iXtwhJ
m9G2EeRIEeQzo9nQ7xFX41yDTxh9O6MoRz9wtxjvtcVJQ3lJjX1drX8DRki6y/1v
Jzx/ZKCoK5+G/faKDek7K/5T8z3eCLAU8AJhcg19ef5O0avckKs3eulw5Wm1HoEe
npJJuF9jr3Kuw3SWBnuu9n3dppquVrRAkGJHlz72BZ2UypU3AIkZAq09Edw7c4tp
s3D27oe6t6OIowGModKz5u5e5P6NduYfmDSlkHjvTZIYHEMdum0xwYxW72g0CJSw
UYT7+GKm11THZ10uLKMQMiqj/i2wxeBzPYdaHVnVh5UOwwtVXIcD3eXIk2m0tzAy
iUyDhEw+F8wspF4F2iApUHkiQgMHdYmgLEUcApFSIz0GCOg3zIz9O9hqwmJcqBfs
WQkRGALM2i2vRNw/LmQUDA8wF4NIRO0BeV2zn1LlPYd7+QSLlbgJw1ygnz/HjVwP
JroRO//4IXK1DUGKO74IFt9tz8gCI28GUN+jC8G/zhBZYBO1CxPQhQvCjRPYqbuM
bJ3I6o3rj9llFAyMZfyVpdQIugZfBl+W/jsk3vpbEGkAx6ddTGlCHo9tiJcQkLKT
5KRSr8jgGmbqWL4zhF3mSkYcW+t+9Y7er82BSxi8DpOtmME7sxI9hNPY32l/G7r2
+CEg7mDqWm0lWYEvceTrxqf7q9GWkkArKG5/AxXLPR1I+CgKfpuZ+PlRgTthbp5S
WBGoF2FjMg4wpEcir4NGnlNVFwE61A+PhDtBJ97dkOvZptFOxuQ5cdOzNHIgpw05
KopjLh0iZQpvV3Dm5Tt2rcPaKb+LWmHZLhXMklH2g4KSEQ0yruGdpxwHwSpRge/H
kBdzLDYV0cnh6XTSX8bYmZkwwhDJ78GyAIln4lZ0/eUvVIsSFjdTUo5Y2N9zjD3Z
SwXq548fo0pMni8BqA9EiB/foko1xXG5SvstzmeEjlzgG1F3Ii05oXIiQk/ST2qK
HRMJ1oRs47tKUdSrWkzA/4U9kzuB3jN3yrXw+CbxbzQJ9BENmHg2Q29E4RLijPki
c9AL2mjoFlkeyArclC4Sh55Au2ck7LLms8Sc7mXPxdXhCgmIcHnLkOED/+FWL7dN
gKu8yjOgX0a8JkFUkCJl+/Vqr7/si4tEJ1h1cJQSw5kTwqDrtWk2ddMWxrbi8bvr
QrRzWQ6uJtac7Ud6BScc3XFLdpZr6mOUgqTpDEH8VCJ0yYmsw5d+9w0DkhOtlZXz
mXilBXKK6/0PDViFRm9+ZyJW23j7NgWPAQt94wtqPjv4QtyPwyo1a4wPXcLJBM0N
jL5RjvMlwhpJzqb+3F+MuKNTwhAU4M+TnT3wOOrPvp1d/xEdiPQHQz0SjbdC96yU
makltonuRjnX5HwMLz6amxDgXehr/TjyFwwRwLo8NBNkPzexrBk3fS2uEbXodkbG
eO/Hq9ckreE6yblADECmBQSySAh9/ITwjHN6ZB40SKf2amk9MGB8DgXRPVpi2m5O
64yLajqTzbz2n0OagzOlUCrbhoLQ0GtbZrrPFZoBzgF0/lP5bokmnLgsCOMh9XMp
JeKjXR/paomoSQ1+Y9/sK+F8/AQHiFGYfP/0FPCRzf5UZPCb/kt1lgGFPf7cTroE
RZ2rT3Vp36Ilj+YPUZXjqyBIU3H/Fm00osyHn5n96itUeT990D1lJzrcuYdugc72
OgZK7OwaLs5OR3Hz0lkqrZarpn8oke//YfLXbgwQxuYhbWWcQNvQtlBwKepJqLqk
iDcelg0t6IJ+yCmlJ3nadR1EbTsYrwt+hWmZn5lgmos3a+AeAqvli9Ywy6XpnqgG
1D3Eez0p340oS7v+udYs/BToPyamNdKKxV6gU2NLogneNl6ItZSRHDwjASVYxZKt
6CHpRU1/zVyapLrX6iRNwrK4s/K7smr7r7TX+FIkNR8VRs/yPyedIbXfHKAK/3yR
d58I8XMdqHoE011XZQuIrpRAmkoZS82edv3G29IgNSTLq2lHOAi+jXAMTO43e0No
hvEUdLsjNNkjLlov6sdJjHQMEkAjXoCDDC9deuVupRx7yHRv3+DMW23D2bsqpdpI
bnIAQy0KlRBqJeyybeVT+FsM1YvOBuVlTPJWZGO0Lnc3Sczq68HBrQTCBSL5xo69
So61VXLpnjw96erHZ68UggQ6phbA3Jm9OHvvAnv4UrT5dvmMq9IZrdFvVNJkrv8P
wyAO42CCzw4Jjn5zP2pviR6noepaJWTJx1K0WZQrZe6UDJ64xk+DHa4lORbhwn6j
2RTuSGqige7rc6qqv/hBc2YLPcRgnGuKtcWs1Nrk5t8ip9gaMjvyWBoDvQGjPCed
mypBCf/PEDMLDto3Fa0adrVvbBbkhEQ7vltfj7ZHy1gCWOA00rldA1nJrVjzJDcm
DzPTextZJR5/b27diB6pZEBQXqnpI1VJ/vXNAX90Yt1y6I1gUsOBBJZ7TgwfM+Ki
pk2CJ+b7CS4fGL38Yz5p8oYX9tpap9UFFrOcfD/KFRslK3XABAyrSDyNI3Ox5wPZ
gzFtltJJtduRdzJBS3fHKmtkFlswwf0WZGS4y+t6642ZBjWjU7CpLs43Cz6OtDDV
NBdpbEkrIFFHpeKW46ZTxicuJBD1jbfh9g/IyWkOFId8civVi39eP4owioF9TMJC
iEAUHIfvLbsf5/LB8W8FSFUi6ErtrKlOkT/2nZmx7fQPYsW16YLK7C+BLAU8NCQk
p5pxpemEQWCJqqxK4QhbOhgQCoxCNhmIGOdbR1wU3KiQBLrPoSvnz772vk+A7GLq
8OwEt52wk1/iQMzrIc1u+3Z3w0lQJ05n7HoldLEf8li5SOIazC0JL0f80rwNgbNn
H0M3XKMhi0gUlf7wTJzx9Vsgpro6xwS9yjZg475vigjbmhSz5GWVHRsJhiSUpqqD
AxqlMX1eyQOUeOvkuHVWA/Ro3eLQ/CfRAc5adZyGKShbdaMXUEPivaH2flD20KQG
YuktDXQNOFLSWoTz01adiydgPk1sNYYL4vISeY5XTe2BtvneIJrHineTiwtLthIO
cCOqElTxszThXubbnPoH0YeVGDZ7jN8EbEnEiGfghQg4ZZuZeTbNj1Q4hxYzsvay
onFDDR+wK6JM3vSLoNNXjABIFlvYBFL41hWA0JHCVxuGu4tuq05X5CCWuUpZHayK
4QABKCVy5baof7HUIUbkKLm3xRrErmpD8EQC0Y7Y78STOQC3z9AZWa+cSZ5xKN1U
BtWrLItzMjLjyj4w+1Rhxo4e8PTpcKTraGA1dX3rvKvSrqW7PksaPxk/dN6AF4ZY
QcQjcH4I0D5qeXVg0C/cF07mrxyAA1gC9ulP+ujB63blBotbTRfABBdmeEtb0NZS
H95B+sMN+XuAxchCjO8duQQUrz8nv3F/2aEtS7c9tUIXPZPiv5BPoQ0LGuW/cDEK
zq+VTDnfGNOJxJrI37eorT6ldOXj67Hy6ek5jG1wQf7x6roHmzNa/P3xngcYf0SP
aC51bRQM2iklQkknGDnm7koWh2E/NbU1YCxDzU6aSd9YtawykffIblOlbrGajDi8
5/nTeGnvqJe5MHFGtsNz+iPP+6ATVPwDKRuY0Bg8kQKonF9SxUgHzgrPdtewIss3
mBRCmAKNGuIB/i+Sdc4hjr2IYSGBmbEcu/q4bGDKG8IVhhuReXXhBQEbBI55Dc9D
erfke8/wriWPnjtjEx8YbT8GwZRcu2ody29EqZjwVW11AWNLmYAYCQRlx1xoitUF
l8cKCX7oloJubluYD4Rrn1DT6Gy2Gw5FNePqkQ9rHlbJVsxZPRlrWvCWAUY+yekX
Z3MsI4MU4P4E+jyRWRHOvXdKrUtq5Y92dAibqXHxo5ErokMnrU01tvnQHp7oK1Z6
Xmc1vfg0rNiE4ImUlGm8zcyoi3RSaDJ/+N2AVrkBcV/Omjyz6TPrQd9Fg4h2ljYV
nm5mqECq3/9Wem8HnuF/V7mQ1t5BK7BqHaia1MSbIGGakOtGkNDeRtytqKLVdxks
2dbepRWm/OSZ9z+qrmoA93jvmxmPcRGbmuMjth++YRdOFfb0FlbpVQit7RyLsebM
hi3PU2Z+3iMM9LtubBJcOQbIghkJmr3+qpSBL8mQsoLprIoCFjifXLyzlSOFPXs4
570MCThKl1sAC5Q2QqX40E2octcNOWSy2nf9novAb3Sfek3QlFACHb3y6qpGU5BG
zop31vluXAml6fQHCEWP/zcKDYN8IbcYqP6/tZY4BisnKkYsOjbJ024DBciR5CNp
2yZWf+8NCivyo2/XO6U5cAwGBIb6zHxIQcehKj1yxrfY+g1ER4JTogJAf7OJrQOw
6vjVs4zOfQ03//LMLrDpnRFmYqZTc7fc9KILIUkz+LKACN5v8NwlsU7E5ZDBxSlm
BVupsdQtQvAeiLR89dI/I11sedc7HWrNvyIe6awMX21UVNIv/5zW9npr5xrNpnVh
Mxl8GH7wbPkb9FV94Fpu/u7oBTQiqSzFepseFDeq/Aq7ebGPn2DxjICj4xgDur4i
iSGh0LBX1SDJdEQKhn1KBAm9ZlfmMjbYqd/u7c8hK4XRH7nZHVjqUiEHGumweEIZ
qFOWalqXTBoOjRxktNpo0ta1kewd6eJiDakoiQpxCK3jOKkuEuJ7gI6ErktD8IEi
Rcy/QdVK9T0+XjovI4Dp0jvef/vIcIarus/sDGRFYXaept2pEqXJkxM+vuwrZIo3
GA7wOyY/VYU6R42Mka6L8DpIXmBzXu3O+P7Ox++tLacdHJngtqpuJ+VLYNPoxQj7
wB/XXhmQTqyfcHPfjGsFNBM/yIfudIyCg0v0W7CRThMK4eVRv6+7Ql3s8aeHUJiQ
DjS8hqbltyA0aZlXXZSEa9J+QRgte4KsgAKU2+OPMDeHXkaq4PL4sQnM4QPXU1LH
hq7AjNsk3V3ePadytGvNe1g7EgfrNFCquggg0UGjpkVr+3nLLc0QKFYVHZhZnW8A
h8EAOIpf4g2Ge49P/G/925E+lABJA+xCRgmULIOR8/v/Xg82eivizVMklDn1PGEU
m/Z3DgTfe72JEZBD5kXs/ae8cBusTGiAv3vj+sVD2R8DaWEGBaqjp8WeCZOPF+7f
y8N05V3P+T4MHIVzPQBYzOCI7F+VxczW5V7r8DXG7DaUKl5YwADs0zElOGMsh2NZ
vg+Rw7Md+S7gum/qcnZyxKyQP4GcMvEbjZxFwIBTMDCm3PQ0h1EKw6wwLNty1dCp
wAq6MHVDtnVUSrsfpYKR0QlwbJkikQcN6j/E0MgfB1iAsnuDL66q4huffZt1Q+wu
I7BSXL0gcUo4ks9wl8Kk+WsezDRqM8sCNCKSlZE0sqZS2PoZXHcbB9P/8+Po0fXr
XvDdPyV19wr5WiV6OHqS+gIrVgPZLyFE5thE26NIf4VCY9f0wRj5H13MdG7SO+So
rzfEUEmZ/2i7wLvVnMQGME6w+/Q4GC2xbqI9Yz/X6DPlM8Flje0dHx2amt9h8znk
33wYqRAxJ/bJP6kUdstSgrdokc4UcNTEt1mk4Mr3BNXkKhWaNc2MJ/bCy5kb6HKi
4cVe0jUi03q0fQ0G1XAotkw/pkkjf8jgXDyCYAWkghkCuD/6VIYnBblvM+yKpMts
q2LxX2CaxOQvZli1gtCLsc1T7hSV5x0Rexo88U5jbHhfKZNiGhnvg2+brjURR0qc
1jgTDmK4gbqEvJnDpkCL2zyVCqL/Rl1Ez7ihCC0L44vtGF0rN/vR/0noOz1d+5VY
DnUzTPvvCfPKfrGQ5cr4H8UBe7eDeY11aMRHsK/7kbCzuGM2j8z51NS8x0FWmdCH
n4Jx+UO7je4bnLGtJ6s4qpPR0h0NvYNzoCYm6M3B7rn32QditiUTygXej2kX61uN
7335zUTETaskDJoMqEXVBMaAMZ4Ct0r0Z4RsaI9gfOYRVx5OjgfG/+w2o4iEGs0e
JQdpYeolqpiBzaUDPpXX0GWHudaMPqINjK4f1SId31i6zA98ihv9pKV64dcpGyLt
PFs9lmudm2Hj34Pz5pj5V/nZ+s2kn9biTuBQsegn7zN+L/BI5XbE5TBFU+8Jq5KU
9mpHvHnzJQ77KSRzTXLpe3c9lpO4h15vBeAVrJ/ZWmeLnO/2UDgeKyRyWKXrLv36
C0butL6Zms/NPvV6IjytY70CcbQJGe79qoVbfZswJ0AA5YMOgc3rl8JgAD28cq9o
28wCDhhdPutRc0Uc6m3GB7TigBkx4CPKSKosUe6GRY+Tuwexd/rjjOXOAqmXklnu
1vFatfANMxuqgx1JCQ7b+HrXXIwxEGFWtHPOr9Ob6UFXHTkQ+uJ+zoLPeytLIXan
B7AX5ySiqwgqayln8id+GxhMHyeM04szt3vZIWpL3zzm3TY0T1QKvE0lTWSJ7aan
ha8boC2kEmry3RL7eqA0Q8r57TrjgyGOA8XkbkkrJBnDKUGpy/cbzIeyCTpACmNM
wJ9w5d2TblhkGq0kbC4uPn2ytpYCuxKQQeweA6oUH0+6G8rwssvjTH2WsHd1Do7h
82wE5YooOhUv+Xwzx8+5ekWx/xYSH4DNSQqWP9bqs4H0PnKxTD3G5jROwQeunfrV
6dm+nmFrw+Us7DYm3nfTaE2to4ym2gyxNdY1r3lnflOWJbu1aKuefFTdE/K8ftiP
UTT+pcMGj6cSv9j5LWLYVgit51dSKWWRScqc8uknq37QZpXB86Ya97EvCKrbG9uK
7PgBMzB1pvLuefBuvYays6E5Kj8I04/UUmD6o77I1nOVefKaRphMUa5D2OOvCXXO
D982X2Fy67WDPDtI7jbuLSjkqtAltCpRZc7c+YlYfRw6Sc5K0JJ9Yr0S1mdiJKjj
mzwjTHxzaifa3FDoqU0PgyKPe2pCWQ7hu4P7OW9yPG3AmZ5FNZsdq+7NMy9KuaGw
3ILjZs5frS//C19hvMTHQeyJGfjmqor3c6ZMwEaVTAz/KD0MxJkJfo28SqFAMXaa
+Um2moGMbxS8ThdB2nVkUa322ZTxlKo4GN09100SlOyFLEG10BymrKjquAGpBibb
yZ2Ce3pb8004hMmUNHDTWRmUNKzQJw45xdZ/IOKaaD2+81OjY2nDT1Pj/9UGptGR
PgOnsvuYkIvnpaGMmsN6bpwv9jYFgZ9xkDmx/jvPsQE4MjwD4Idpigtn9Z87ARfY
6FeSyW/sZ9Kbitn31Oef6mnaajvpp37ltB84MPtiM4kgnHSB38jdGXclcWn9HrHb
qi0YbPpNNCPvul0Mk7033EaLQSPnm8sASGSt4vLiI7pqBd6JCz2V3jSoE4pFUWx9
ZW8nzi+mAg5YfnJXCWi/4GdSjPJ6xDyStMnl62yw4l0moD3kvo1wxd2InlA5DBb3
/aKS6yVMfHc1LnR1rm/7JhLr9ymPwsYgJ/3qBLf7UF6hPQG80kANOMh1KZFVcAII
yWsU24oIqRRJNHbYVknTv6WDkpmYgDomt2z03eeX7m2FMR9fnV6LxSVOEPDLe7xY
gDGnqd+kYjRBczVEcPDlXGfhuQKhmi6cyWznZ8xMhJJgvdWAcpzKDurF452j6WDM
e/ziwRO1gKifRDdYbvpZmFL7tYlbOd74+79QQnLruQFT28njcqp5KChRqDFilFOP
NuVzPSDx95JCLX9Jj7FwHzHfsONWleyaz3ZP+K9w42h3Bd89HkpxUGf99C2qVJH0
n16q0cSYDinOxJTFlP5Yw7GeKOh8JTgeBqBmzfqGXQJOIfr+NbHSP/7sLAHF1C9u
OP7Rjhyyn5NB5faiZOWolA86lzpagp0QpjQmEbivcjUksiEaP1MNs2ftOl0hVcEM
iz39bjjxLhP0/l11yp7w4fmGNSPW2QVrreDfdcrxcG/oEIsxjGfZ24NF92alvlV/
P4w7uCRBFimz3ZbM/O45EhTfmGsB7r6ApYqKPWrnxNwe1HeVyBJcjEqiMeq1SyRy
bc2BZxmZeBpLa4b3XY5YokBnN/+vRgZK+tFqq0jvTx/iaxxFokNHDZi0sziUmITm
i5HylULwfshWWbGlcDjQweXVwy5lZNuxeCpSAHePdF4b9gHDY6p70Aa4LoswPNBo
3GIGupHzSnCB5gLaXmGK9F0nhkUzAIURsWuGERfC1bteYKYSLNUhtt08eoD3wRi6
jo/8KjN+7OQEbMKcQHf0JglgKyCQamPJEIRW2EGnLDkOUTOyTLT7EgbxL1Qyi3Bq
u943q2yaikGeQSn6EWPM80d80Sez+aeCI4pxYAV/t3D3qTkCwVuQatcZG8r8be8r
SNTfg0/6/TzGoC8ZXvMq8yVf00eYG9amsV6YwjaEpNtg2DnfDgajTXn9HEFctTUv
2rDxDgv9fTsMPBeXYjq1DnwQk/Xo8xCDaQ2ALAOhW4MuGEedFjrjaIDtn2E20KCR
2SRZ6NkWBK4xVCgy+rZ7EoXZ5KTjwtRw7cHYzJPJSlMsYw3GRGFTWmNOz05y83BR
z0OngWt68Xmh3hxBoPe9aocRAG3skP5wmhAeVjhqCb29WPVGCx6NTq/zL+9cjIW8
MkbwswG4dMilIzOltutE5A+qkZNb2A1sSseYZq7hU3Vj1BudV0ShqVGQl9gAS7fW
WjgZ9MKxNKJSoT2c5g3wX/cwL7ZcRYrjxCjKAQnvGpYNUxRsenlWqLVme5L7jyJD
vzWRMqJTOPFqsb/g9qefPKzQeX6r8306yBoRBNsXHmg/MmT+BiFKiBvZmLt6iKmG
tM1FYRYwF1uL40m5WAQj69O97zDzkKUT7jcjLRlXnYD0m6DonCw0cNwGeK7PbHYm
bYmPQPk+FYO8as9ByIA0oQ9YxVEMOLFpI7i6U56brM+A2PHEkHU9jGETAyzMlhR8
LDUt5GwPDyHGGlPkbAhpcXCyV4R7OkxAX+V1YY7pknScYukkuZL4BDYSSbWTq2ba
Qcho3JHz3Wmt0GTifkqcHC9NvNLVmaOXoLRRiBRkI5ZINB+Rmq/0XYgOAD/59br8
MmBhhBXnp9toWThs3APfaYv6rZMBY8LUek6MqFO15BDmJFoSJEUmM4xziVZ067Wa
AkX3tJYBYI9YyXt+jRMFGb2moFUTe21otcFxINuET3kY2Ugl7NR5bet799d+JrkL
b5a0zLOT9HgJWFJd8OBxIxKqYiMn69ulbbiB9SHdpvqSvLyciacu0VniabNMEHlh
B7rjVi4kVcbJ4BfDHTN3eM5Z0yoiTA2EtWKZyb/W+k9miHshZ6a1LMTebBB3JoTH
B1ayrqL880NtocKp+5HAQDDTCLOtj3Ah8DAFIacUhTe+ud8L52lnwarmRVTzQNbm
BTgMz0uaHLcZ4+0jkd4zlYKD0cl+v4Xy1hjj9ZM8Eujwa9pFF+qSUvZ/IUvOWAYK
6y1qcve+DrFILFE6DQzppoWv8Awl8MjFsh12XloA1G4ehgAy8bQXytSyB6urNEDu
YtSYaIq726wVHP8rDNMo8SVH2lZ1V7MVHlxV3fP2VHdtpYeCbX+8zN1itCmWJmiU
ucSGwKBEXsATHozQJieGoMXzFhmSheLMJeDgp3DT8loBdC4GoFFpfu+CfD0PcmAj
3OndSWWOCuFOElAn0Ki/Q5/PizgVaI2Gb7JZMKMTpM8Y7S3JFzKUe7dy3vvhfFBQ
hP7b/dgeGoUd9fv1fUk/HX4UzM2aj4mDY28wQoPMqmIDlOFWHLc1n6S5+hrU5uS3
wg/CGzaIzTEKJzSgHiyTMShY8ifJQGT0BReUMTcEPe5bhF24sbaN7kERrYHtJ/Lm
uYcYobeIa/TQi6RiOX9l7XD26YVJIqhsH2AkwcDCUedlj5cXCJT12JEtan99TiGt
+9vODXwyHSzTYeTATUSSPgspxmqWkvmR3RLIJh1J+9bAtdA3yHp3X0FhuZ47c6wo
fIfV0pvmkCS+wzxlfJzkRpPvsUzawNoDfc1fy6UFnWkrAUCCULbFdWtL3JLDyksW
8Sp4INzWb2mJ3JQNZr9N/So50mbGQbWdQFf53j4CWYT4aO93yKfYoyxvN5n+9CVY
Jaeqp35hRapnoOA/qJ6tSasD+3F6z7wyEIFN0XBmTIVeVCMU7p3yDcbZ9nYBYkMU
m87ie+q6eImJJKAGJ1danb9xHpi62xcmVc8aNd+RyldUGa8HRjCZ+QMhZLL728Kg
U4BmPVhB6LVNtmFlAXEhggr2mhoiJle7VXeCpCuygNZwAmnMZkGoAKM1Uj4pdLJx
8p1cHP5ElWZeT+S0XdsYafn7a0NhltLGSvuXCI9CVmrt6JXhf7GlvY95W1q3ozv/
udkr7GQL58kwSCbwSB3NCb5k2sFWjg2lhinH4vSvkxChWp0/U0Wk5zdH3hVXo0V/
7U0w9qTg+qqVfObVTrVxzWdwiCjEzsl0FBe5fpD2WfRh2wo5uHoJFFdQXFYgNv3S
1eeZxua0XbJcKBrkhhGUUA32KxDDFQOrUcjh2kgB+/N0QiM/V9eq9usmgg9rhNR9
8LyCheMvdUD07CkXdfb53t74GqoHNtIalqMYr4lo2nmWFyWGj3yAE35I3HLdCB5H
VPCVYyZePfZ8dbX4zlNqJuZg7sOnKq4cEsT3pSsTloFNrYkBTAN9h++XgyBnrlHq
hpky1LFVhOl2iKXaGZYSD1RknnV+7RWH3KucAc8BfFvwHMNjyVPwWe4heWdsKn3m
oTWXTexNQnpWUVuFWDB7TPkrqN43Web1hLfvjVDebIzsYbho77lk6QMiYte30RpN
80wzwWO4t3NUndCtuOcD/ZiEyIYMh/gUIBSXZ7VdA9ZwG1/d4PrA7DrwYkUA85Uy
4TASjN3qKWulgyAO9XPxe8aM1Q/uvs9d/sGD54WgPaf8DSzjB/eb/1JyYrKV/6oU
VtjitfK0Hg2Ou0Xuacw/wjtIC+vvtIy3N5PieArGG2QgSWavpVP7BZ0tZjqu1WR4
759bOE2jgA6ptQcYqv85h2LsBnvfsV0C1g4TNof0M75MSWrCcy8fDsfBtoK3bt5S
XNYuG5VY4OOmmf+Sqskqcf5uLeXwT9tH0d3AnSshUJVUgc0tYRBtg4SrV5OJGEn6
yqDqlJJQ95gSyYak5yFqTW3KoWbpP0wujszngM7NSQL2/C6qwONlDH3IaAXmar3j
2EB3g9gmiKk679VltPGaIkJ2eXVif4o18BHEqT/wuNCZFXrFHhS/uU7mPKwL4QPA
oOWR/wyqWwzBvSZ3oOwIqMK9YDaKKgVfOq0pnuPCZ91KuN+qfZKH2KmWzcES/GUa
XBGA1T2etxa8u57xAkqF7TmApVGSTudrwuuF1L2uk9M7reNCbA5tkkMq3z57Ozxc
XBMV8w1A3NQ7baTT+bjLdCemyM7DSXpdKbWDXkGC4Y3sZIBAEZQuOMTVHxxcD5tN
uT1exakYQMplFKO8G7f+bNlUB6fOvpsiIKGRjDn8TqZQ9WBk3gIj/oOJkYlkUI2t
3KeV5omTfLIVMiKvyW627r2wrOcIvmGADjr5rn195b6TmyfYxhihAPz8plgP/008
3eGRYo4siATxwS+qb4EBQ3d5Sz+WEXlBnWqsclO8BHca9Tg+Z8r5xE6DinxFk+hQ
K8hkthbNeQkFClzlrssYad3pSp1mzP91Q2wwCPmLBAVICv+eIrrD49G33/cJNTij
8+OzJLld1oyjB1Qkgm6KsXfR/LtswTNw6XspNt2gp1dT1f+kbygnxjRGkk2wNl+Z
ue8UFaD2b2qKtqFYz4XI1M22AH+FtnJKITlPFzdGCkNiCtnpc/2xKH4SMq8CQeIy
IzsYgkh+vVbhMcz+9UEJ3PsaIlX1q/XbWg0w4H6Jq9z6zwEej077/esHzdysjVZM
IQPMJIK/H0etudwCKoNnRefvh1QQTqfPwn+WrZQGByktWgjSTlsaTFISihf+0G2X
ZJ2kBhupNVUeKFRSfM6bnYUXqAxCm4/qy2yzYlplfBuOOM/GijebDe44DB8vzP9i
XPwduDGKj1lUuL1vz+YEPHKvu/sGqEnmRc5XFNy14K4NZTJiRrn7KpfXZGNX2z4E
HVGl1y1aXVcahsMzvURO3cgKwmogf3P3jIt20hFR+LKBYPbsyYIT9VM1qthhYUye
O+i5sNufGvYhbeFPnH//frkqF/EVrgpIGT9ZZvYqa77pQ+GDHxQWj//jG1mUkvNH
UX7rFMzVpfk3hi3rxYde/5SHE+Id2M9puCzD2wnevJWPmpGXZmrL44hhyTelUMLX
2zdVGNj0hAMe7oEHiyBL9nUyQMId0AdmpPVyi4hqgfl/otlfNKlt1+p8RLwNT0ii
2YyO9PAjTJvn2iISDbLnOjT4ljUAakuZsDwh4WS5Y+nzNNN4C9zrMhoGIC2zUNrQ
/irto9hUykXg0Noz+/vqW6KBvMBdY5774QMb7ghWRL2HqxSQN1lYniTTfyADmGjJ
Z8AEloZAKqBbcRKkdfB02vOxB+spr503fAENVmD7j0JMY+08+nAuc8F8hwd8JRDq
mWLN4qYLxTZ7Ek8GfJmsMhsr3oOUmFooAoQhJ9LHDRL/FHvjhx8Xi8N9mOCcpNt8
Qvc7u19s1+5REahtK94HQyXt9RrbNKzuLNF32yFxkupX4afCgd1FuVwv+StdIgoZ
dZthmFpVD+xcHTqQYm8txOQspHxDQmsEyJPxHJCGvQC/dEn5j2JQc+pjmNnqad17
DNgWeyQ3diIXc1YV9W/riEcamf3K1rigK6xgwmkA3IL2aGmXOlmOWIKq6vZamuZx
fArbHbxS3WLTGgvv9Hm1b16x+Ov4MlSNQ2sIXmuX5ff/+i6LBusOVRwj1kY2/TLv
ApPU2+R6/4BJLbZXgEwQJmD8VsSLN+soF4utJqvu+GRyN80KB/uqN+xhJHXRAX0F
CvMfXpZLMJU2MbqkDPcTVAP8ptY7Ddyy75tIREMCGusvtumqLRy5454cfZFuTCuT
c0M8sSfWVTI3bQftphs3oConXSC4aUpwY1sUOEduWrvXcNCO+reZ2YgsEc7dFOwk
CuKRUEr+LKWwyiqfwJHT9Vp67ix1mMbaM7Bs4jffQcv9NOV60kzB6BVMNtiuiJ7w
vw3wx29V7b855NVfuU38XYXIKMKK+KKzHfZD1ySyvX1UbpbTMLdydT02kEYsLoNu
h3wD//O59nqwW2ttbH+AMHj1eeZ64fVkAQnVqhaqSCwelPWln8Unfj9zpKQ7ECzZ
am1eZTh8UcJoQ1RTjmoJF0jQwB4G3/uGUbJl1vLUQ5rSHwzr0eQ1ew9Ac+U9KE2f
rzAizMJTRksccSLIDICAfgM2c8XZq24dvOjdIlZL9GjjF+O0oNuitmIpS2FHjiM7
DlH546r3y2b1u7hkK2c2SfF3StR9lS6aOKOCmgT6o/Y0QXRmVQ+ullf/ey27cRAv
p9muW5eN/Jj5OzkH/d8J6SjYf0E8LkKe0MmDPeTRoHghqPp7CrSksk6DXe3gbsJ6
mLvM1BRyguDknVp8RFJXlcIzXDJScwelW9JJAOIGfBCpSkJ0vejpMid8xkBwrAqL
06Esi+4Dvlh0LEO2OKcVGdu6DYJAD/ACAPm0qMuvYcZklbL0F79B/IEULwj4jS40
LDNXhtA+yH5f3u6gQzxHwPoIV9erP/ioi8/WiNMdK5jwf3yqI4fYUIxwa4h31Z01
MwGpa/rwM+MqFs9LtcSdUJeX5ypxGh9uV6WFLQrvhxIYrdweLQ6OsxlCKy3bmKZb
2BZkn3yJakDJjoG+UWlfP4btkjS402KyzbfOc8aOnTPnP/zLtZxnEodIhcjf8gNN
gBLVqxoStFItyFK62wH45PZDa5CWuNZja+pNIlENbidjU2cQED7ONIxjjxJScCw5
KhkjYncZHEW2EXI8tI0pmlK9VokU3jjvkf2dtTmRkE03Kle+tAKHIGwXnwrvFU2P
OrNxveuLvr0o/FxI1ZU27v0zVjRkyUVpN8CFptl1sGrZJdEOTGzhzGANDGmabxsU
X4WoQGPCu2O2urergbl1gwkKxhsuTzjjRHMIBT+aKmvsqbcFaZLb5gK3+G/rjuST
n3Rd7mKLH6N6fWOmF3eOs6J/9aL/QFHDY6DHjjRvgn5Kyr/iC17NqD7bgfUHReIJ
uDu4H75eCSnPSRTMLsccTtQBQJwybJFtBzOkxDuaCtQBDZuTrnoCOdPzEvmE5mDu
KUdlU+tDYIVyYlJi2fFdgQlfY1EEyVcIBBZOvZDWvI2z7hCvQVcVqVSjZwTAfOLS
I4UChrj2Bc+L+Y99i91JZSXpo4izGAHhRRstTkLQ5vtOLqAl+PbGLUc63nxmpF2P
Fsx5OaLlzlUQNB3sqhX9PClmCZ2J9Z35utNGhJX7VvXeze2/93cCmWilIbhPRfBC
+4W6AWSBbgEQzRWG1lebVmPDczEaoic0drn3CjO+HaWTwXpVxllY6xoHx3G3PmKb
Zseov+5eWSraNOhuxr3gGCu0eRbLtZ/d7BDYNUxs7MXiuRr/zmaibbdrApUihSBp
hx7zevEYZdU2n5QPUCeMFEgqcMy2VOrAuPoHEvh/ppb+qHNzF04g74rdkz/tzDb7
mGfRvBgH0nBcVqm68/90HDRBu/f0TLHWku7p0VLL41GE5OFq1dXnBsKMvVFa25BP
e3KbICGooKt0TnRmVSeoa1j1xD4tyHkNKQrfkH5Nct1kbkGBOUP3oXOvRhLXu8zi
Evd6azCkbkncgS0zw9yWJwltA8LVHpFaYZHdj1WAI9u6CTuEWlCEihf10g/4DFak
TZhTJ4dtEZ5u8wi/il1jwFufRXa7uteekZGC3p39PzPshNnzUe5XqyPqiTyCQYWV
11uuUOZlkJwdJZhLlJJHbkCgpqjEV7A9EgIHXTx0a69IHN+JGA+mAck0T+VEH0k1
2oihM620DyviCcB406+Y/jre+83ljmeL+P19fYHyU1j9wA0Ns1Fcx9LqmznDBts7
f6d13Y2Q8ZE60+1DVmRvR1x6omipPt3aAzAJZZt3LLkqhpPzMQLXwIO16uzepJBy
to6wWYzuXlU3XewSHitLigiPKSFiUzL0o/gQI0+yK/+BZzahlQdXl0WEFuXnFRu4
HptAHnXNdk2RZ+Lmv8oyH7DzBJNKe9W0bIuzHbIupG0ZMkWlyLvp6NL1P3BpN0hx
dEVfVJyKogjF6W7DX4qpLTFcgH+CN4BbDyw8L/mBO+yjDWlqPVW6/HT1iLYteD2Q
/O/5zysmJPEqyplWIYJb7JoOqKmJd3CZzzmfwTlqNxxXFO2FEnHLbKJ1ERq8WROb
+DiX1tEbhzju22KCdYA4Y4FQWQGVyPLTD9xbApjtPyRlzRnvGL3LAsHXUJz0t+yn
LN6cm+Q9C3AQRYqd0FHnX/Eavriwrign8qLonH+lrt883gq4fBNmiYYgKXumD6Yc
ZAOuWffUMFMzhUJ07IYzc4c7kfvmkgBxX8fG6BgL+TEeRFw/FaeOpCcrw5IHND71
rfxpR4LMBhC5qA5buqNsnxxmuyWHxth0B5gx5UK7mkeNLOpJXx9CEKHg7mSMGA0w
xYIecYNPGags9ido6BnMb7FURHi+4mKv8G9FFveC9j4T7C1YiwEV15Cskh99xtDC
59VWoS+4nbZ6Z4JDTTZ8MurCu8lLIsQrE33QKK4uQ2vRtwLu17nEO3EmMv8z5Pfn
b5jiaTYKLxlc4z8WkoWJNuTXTSxcrrBOT/xcLiCkll8wafoJgqs7eZrYqoidPWJk
dgj3+oHFOE51u5+RQtH0unuPk9GnakTD1zRKzovzt6M/TwBZblEPgitdkBmOaylZ
4e5qycJtnk8DK90Zz+V+eOuAm+9GBNe2WbtaE0eCRhr5XqFUyhgpqeT32NLVzzgF
LMt5M95zz7WlmHrElu/yPfci9Oqh1dku7fnmVcb05NI6d7jX72ateq2W9eNa3Wlw
ErfHan/13FiqtTyAI8AOJYSPdkW++ncQ7Up57YVmNV5wPoaZCxXf59JQvN9caaAx
XTDvcwosaQ1G1w4et2FQOjelxpRuh/evB9iaE3bag01fNG4RSf4bw7uFI11LdeWC
x+bqYjB9Uajs6rZmLc4PY1OKtPbQ+3X5eWSFhbEa2/2JU2M5cyuupJViPgnWyyA/
ms1Altaql7oBuIAm4hIVoKUYfcVE2HThwLEEOYmR66VqMxpvRiFNBbupv5fXM67Q
hLUD/WDSF51kGBbJdMDWOuPrbXII71XXFifUDRiQPqklRWVMqmR3qfy0mGDoVUJ8
PI1MjTvl/lN4wGttraqLzjvkBTZuZK8eYQhM0yY3gmY0U/menBHUv+aroKOzXB5d
rtLASCzltqWHygceNUKP3Kl3kcieYooE7iNXl68EVHBiJXFUrNzJkFEb8+14qSoj
C6t0gtlndRLW8K85YrSyG/pUKjfSS60q5S5flZRuIIdqoEfNV9n9HcC+wa2u/Tts
zpZCdTmQ+q1pwaYXFjN0gjRHWthsrYOZ8TbpSNdlbbBypaqoIvIlHrfH2J05YB4D
5j70XZu1rntmshXDyuXemH2/LSUwNtaDfXC9Pr+xdBoD5mEY5mLpvDCGZXnMis+R
C2lCF8t0oxJ8z06qcCQQCkRMN2PuCM4vLAy9aKj0UfnvGGVkQu/uv5emzsIzyfxD
OKrmzH2D8/NulLPhnAf0mh9RKuUZ5NmNYjuhHIF28ixhq0V+pyWQr1AJAqPOOc9C
A7g5i0v8+jWUXBfiNFTSbQ8ct7grLV3FpjYV1rFr6DnuvMcz49hTR+eZIhv1AHUm
dIwPSzThbx+G6fA9Onz/41AFUcbsrA+Dk664O9//373A3fF9zTaalv+GSBjRaj2/
rRyrMzLGi6N1eCzkm6O0GVUtfM2T5sEca3C9WJxYwmmsP7CRHVKOivCjNsL67lFI
EnRoSgHy2qXVadf3orAM82xYOEo9FsjNUPq4MY4CbYJGp4d3ZI/g/MmzNl8iqMaZ
2/QE6vTdFHVTN9Aforz90qvVpxivEobG/iCljwj2zDO6F+BAc17H7iUbpSKbokJK
Ryi7of9m5tDGTWrrzbaqiaG3d61hR0dBHRz/gBOWPyI0te9qUDms4UnwFBJH3HGV
5lX3aDcGy5CQ1v/pSgsxp0qCYwwIMG3tnaIdNXxLeAIfL+9aDjMXG4su1mYE66yy
N/T8TKnL6SenhBI181YfOk5Z5ImdSvWuJwmyMV33ySbnnw3Mx6OPGhknqeo8UbRA
WIbuBSoYsveEsDa5W9hhpy1B+lPww9onNTyP3F+8X1jlr4F6gXKP/K4aoff9GjL9
rVW6uJDAZbjFnKdaaxGMXr4LtBc9oI3HgyIEBfXafTsziANWFORVOivA8e0mhC+B
eDeBwKfiguRKRfLnLG1p1ajFB2ZPGI7d6FPd/XyEqoE/UwdlCHp2dM6jMR8rl+Zy
TUa8Diq6ummMQvMQYIibLFuqfcijMb3knntCBeYpOZHMGbBykRqLDhqZe5BbzoFT
ngYUEntpqIAHRuYDDO7m/TUlrEyZKakWsT8R++v2eDMGWhgiNLIdqBfIKi00c6w0
srnTshZ14akEmsF1Rs7L0uMTDFsXtDn648CBVGMGxlxeerPF2+qYV5wzklFAz0AC
1Mokg6Wv4pZngIURZnNNPQLVn/+vFlBcV6CRgw1AdhmuFtvfG0uUiJ4Q7zeK2eR0
JIRxZ4aEymacEh4nFmv2OpNYAePFpP8JXnCcFn1DH/fWVS46Hr7+EQ5oN31yCFhP
tj3GxJZok4ftI0ohOTf576fkFOz+eNWd+OtpqeZZ0CxaC7TsjQycoTf+bSzzti3w
39uoBaTGLFnZBeUKQGdPl6CaURYYciT2pRK4yY8ajsvow2Aj/mhEerHkMaUuzJO9
W04HwXthK/DOq25fqRdrHq0Jylbarxd/Lj1zElemCk7R+rqcIIxPKpJsG6q9KCt9
//hQtDZ7fBofgISHE0eNSkTRQXnCwI/FjP/Gsy+WWjkBtonngcGNRmACC2l36VKk
H+LGHeNjQ0VGNHsB6R6/gU67S2EX9BTGNkchD9bDCWdPGLN9OT1IztZCjA0xJanH
WlIPCiE3XtysQreQiINp4JNARxymqRLESE6PynmpK3cxpTsnAlnX8Uq/tgQkPOZx
SQdOLrJ0+hh+P4nNZfVrGLOUHIFejvk5K/pbn4dsh7sPLgx+CgfZ1qkr1p2U+jOr
arJJ3jam8/w3VDB/12sW0MHzK0MUEafZVHz3aN+Ua3GPbHAaioTfpslYybUI4LxZ
eGcRPOdK9/XOC9b2yJlnutoKzdehGgykXtje8sXYk6JRj4A7MSERwmtkfp9evnqH
jC+DQxCuOlrpG4U1viMNQ6YyZl5Ed734MH6xHZpKfoJUpOvWlJsBANUSPZTTvnSF
KSffQ/G41f5MXXveek0UdfOtRXfgXtl+leonu2on5Cn1Q3mZKlffhzVHaRurVka/
Y2rH5s9OMoUoG8Iic0xv8EV7v9zvsU2yT0BXOIMdJgq0pgDfHViuLCwAdsMGrlhP
94CAefR8BOyBecbnoOQ0iahekU4ygVSwNNOo+U9wJNO4xgKk0ri0s/TPKBAFnJJg
BG9UKzkwnGGXOqho7HuaxqYAdPXhDS3GM+GcqqdOrrUE4jPywM+eRZZyyJi6BNkm
NCrKPXABOWm+70eMbhIMFNQiYF9t/jMibOftr9EPfGpp04kI08P4xhmcIBWPjDT1
nBfmNQqEN4/9RG2UI+ERXdiaNuh/ifylp5eUxNAK9/oGLBwU+OckeFzra+eeVv7H
gqYfYDFItYOskTW7psk9r8vpCtLJ6TNIfY4nW5NKXatF+s7YtEWQfOJXnJtsK++y
3xjMHUXPSbvxWcaXkbNrdwuLf7zFvS2vuJpfe083rzcmXeDhqcihY13BXebEcq+S
ZEsVkd0gww32k5W6JzbVEYQkMD8KFz6kmG4Vk1hVoI12oHQxQspamxp0ugtoLWkw
LayA3ch/cXvgG31t1PWSvEW/7mXqDE3otlOuJR0EoJwVJdiLubgW20loAxjMyyOR
IXAP6LTL4dVHG9mb/CJs9HfvyNjgbw6RnxopVJH6u1aO3R16lkpbxtZPGwg0EWnc
oRgBXWN1qFpXim/NVoyznCy51h4bvnPMHhP46FJe+BD9c8dmIrrckKzLdYDxUWFT
iv6rgITUCVkS2fHWNzoY5XtrsJ2myXsF03HL4krHXDijvKo3+uDgn7k0Hi4GDPR5
XhweA0JtHHQMbLyTM1OGE6lkA7ZQuYV+VXRKxnIrra19u7XOK02qzB02o8FtVChU
kNosJR/f6MUtsqHoTps9+Z+PzFvxeR40i5+hCwgZHWVIqAqmbafAbF4PA937VE+k
8afSibqLihk2TbTVceJ8AWOj8GG0w0qDMyAjQPllLjFM2sGe79Sk8O+7VlcP6Q11
9OIUTPaJDlrnEtyQJ5nKCcDeEhJ08Mgwxl4F+JCRkouRU9wVgf3Pfd8oZPeqDAvG
FqU21a541LVnULdTKC3RHWGrC9GLJ5HbQSLTVH9vtH3vIqxtHr/yTiotU1KT/uU0
hN0BTLf3vFuNbXN/+29epJqzJbJLhyu78g3Ta+YfYAR91g22tYqeFL4b7qXsZxfG
KwrLjl8bhe16TmNwGxTKVBJgIQeHyxiINjlc/154xRtbAbBGSB0iP+aylaHwvpyI
dFExvwZPmjXCIysIIVWmRw+NLZmQ/UDvVYc/ST6gKFxPSPhvoroyloGbySQTehm3
lrEGB3hPm9I6JsTSV+xnlIBU8Y6GPghzw2Ifs7s5RWLLGDhR2KJta3qv7qONmJPu
BzfXGbXtVfQMt/Sl94FzlsgY1dUlBqftRdxBZs1882NonaOe/4GEZQpsp80jto2v
IDeX7PveGohvqco8bJBtLAsBFnlJTc64DjTAEcBfkU6wH3ccljcEwFrvHmw4IKQq
rXNROhdJlHo0RQA4CNyCJESnbAACFl/Gjm0IDO+V8QrJe/MT/Waly7aUbZFSbQjz
IE+M3bqme4JK3CwlJQLmwTU6Lpb/awT/USCOeVCGyf0uGO9qgvCYrKnX0L/R70uj
f7I2qqSXubJnmDo2HNCqlDOjbs8h1I6ek3pwEbsYYW5OSs09wol8WmVHuLsli7nC
0u/ZiQuAtV6RMs3RlPObSC+DDx1vepYOeQVDpdYvIGrjIlA7URB5FiwD9dXPn8hN
Of4+mTdv16/UMeTtalkyzk82hLWh3aiV7gdDWnOaWdBGZ5hz/I4dbhp6nLxulYdX
4y6PdNB+IQKGyW65eOuCixnRj2OCL4KNX+ItYFJZtNZPe0xITAelQ7rPBvgEHki8
CPgfT907q4uQEjn65v4FXvQRIC0g39NiPoZIi/EWSi2zIDY49SePNqbyOt4c2JwW
2IjdQISRrkFO9iJBJkeyjRHVTqY8D9gMNFwEYrNzcgUAz056cCpmVZ0oAk7OCVpU
rZDImcTx8hs1FYOk7giCY/FtXZbhQ/W44uN6Q+mAJdLTU44rIbu5+2pffceQ5S49
RGQVuVdh5RgN8ihi8X6SoBjJEWwcoOpIhL+vWm+4dh1kS5bGUTkLHDqb4+nDhBaL
E17XaY+hm/M5f9tjUJ6oXfxR68hMi2c9mWUwQhY3a0fVNCh/puxKSlJrc1tEPWU8
qg2N0pBepKD/MJDKwtbuY9v7VAge66COTFhfytzMZDH0/ZV9PND1p6DxLagYrfrL
2NMfWSuRtAU42Bsz/ErAxGXOBaTfUmy8GDVGUowE0i383u6tX4p/EfBWX9MvJq0t
93wLrNAiTRnmqVa7ONqRITHvTjLeCygIhNwBSf946WGsN+U7CIPfSCObAVz2mQIg
Ka8aYy69LTRJpfrTtDxRBOTYMlqjQWjw8PPYSnQZ04fWBM9T7u6Ccw8r4gJaFbXJ
p+JX30b3i4kdCQVaNHCWUUZYpjwWSEgpQ/VgVn2zTo3LlvG+/f9NibyOt/1j1dSK
SAy4GPClnQks2u57mU6NWtzfDci01GmWIcw1Q6bOJbhOLV4+zQfCWqT7zydR5Eet
dqy2MDfgz39klGkUrC+EoDBJtup/ItdHOVrbmqJcOWamWe6qnf1nZMuCX6t0Ts02
SlGAd0fVpNeY/5jTP2Mu4WGTZPY0Miph5hcC7ktJA9nCuUpPKpX0aj/ssE29ThFr
2taRuYK5uxcCPC3LhNJ2nknQTxSBjhu16HsdRVoYMnlwZLFFgFrc6Mm/RX7gbuFH
Ukbo6yPm7VHKYTN/E8M04DQxoFqGSeUJTpebXt7oBam1mtVcZ2Yg5XldNya/ckkn
F2Zc5NlmItw9lAcUPRg+HVrP8P4pRo1W3Zw3QOi3DEPuL+XsyBfwdAQ5SWFpnMbN
iNvEki8Tu3+JhXpV6VALkyxMybDGQMUN7QiCfeneu0qtlisox2WPerg7nBqDkqR5
3cCOk/IxB9OYM1bnKY7VJh7oP9w5UOS5aiKQk12uDmUFexje/0I/I+bvLRJLyhf1
xgUS2X5dyeTsr9/t1fOFrmR1ILPY96hWndqmExxOCSJlCv6fed94ejH/htiQH/Vi
Urjgw8HW6D/lnrUDKZSiJ1e4ft9hch6EneiP1iOt0884dtp1S29SNc0LcRsYmK8v
xsOu+pK6DrUlL7j5CETBdmf4u0zA0lEKvK0+pplPwUUDnthwBLfytScbPlXWKLC8
HLarsuxI0Ra8Hz+R50/VLINdfl7qgymjsiz3PsPdyzBK/UuoQ4luSwlhr34oZ7ft
xPbkZ9nrOHtfeOkor1GoRk43fdaAinv+I36SBd7c5j4WrBblG4fe+yL5IlcbiuZb
KC3QIrfVrYgcpjWWQgCsVNT6Q1NQ0kgD5ToHsQlapF5Wro5G4XH0wL40eRpyPErk
3Qbfu0eqfBxiLfvJB9T4zmcLO+aBRGL6p4X0b+LVl6zc3yLx/gNxykkwtrzsgmjC
/31vgAxBKGLC5teK27lVCz6q9TXQnHdo8KB4H550/4ZIi1DZGA8gr9MmY/5DCXes
E8yCMd6pzmYomGlCmGj9FMQl1uztDb8Ozd99VvURsG96Q5cOMnctSpUIoPwqgdBJ
sw+SZVo1XXVnxJas5ReUpCkjnJeBJw2p19qzUNLceNqvx8ydynQp8hpdmBIOYEKX
Z2N5wjFVGya5H8UoPrbOD9RNQVjJjnWpuG/9MlJmT7X0Yl2FsQyX3fL2HUjteiAA
SC3C7F1zs+1Bp9TFGePOESqu0mq11JNDHdoOCZVnaa2XDlGOO6lwtqHfBXBl9Pg0
fEFBPzyOM7kjk7hdgxHB1fQGrQxMO0vUzyNGhMOAXVD6YeEmULa0TrTPYt+Q9Sn9
UIwt1JxsEUHmLlF9S4J+ANHVXoC5pQGjoAs1ddKPTQLC973IPN29BvBN0rDUG5Zk
ND222ULj3fPTTPKMqHak+K/sr846LCby5KH9nIas6VvqA/Xn8gWuGm41uO6MAEIC
vkR6JAy4Nndna5V5Bcu1390RyLGcXhDM08xrOzEu4bKhtZu6R0rrUKE8l13YzxrT
z6WOjNnR7EGguio/dgXzW6iSKXb9PoT0Zxgca4rl1FBTife4fBF5LipKsaFG97yS
9JmhocGC+9PzP52h3iY3VQ7lpihrJJ5lfRW4G9TGy1yz2fM+KhNpnv2wlfo097NC
OnhWKbo3sjAiB5QY/00Qr8M9El6yESqNUyNBTKQ6pHggQPJrAYz2fTTPQs4ViZ3u
k9Jj9C0ga5e683iJKQHcZNd0WHUdSHljUHeuH0iBWp8mm93kyRxyrP/Q5Pt8ULjg
PZHrDCHZmsrl30i4SOrvsJceHg+6THQsVvpRha7RhLvwhgbBjzG4BdCruk1xI5pm
mC6W820kjHpWombe6FZwQRkm/Jhy13o6Yx3M8PuRxGEKP+DNPgygAGnFFw3xXteC
pEmI4BXq+FxSp4LzQCTHuTrkGbGweVBYc7vukQoVXZl5NW+Fk3Iy5kIAUQr61lug
7UzbKBhYYSJdoPt0uRrBKhSkUt/5k0/Zj8lAwV4kZbmZsvMyfHfW6T7yJoOEYwjL
uVtodu0m175VsO1gDvUblzizyDMwoaOeEqAS9kX1rwJIjv5aoKPzmT8FW7mpiLwB
KqQN42oKLU/AQTSFnzrmuGpR57lX7GLSRvXQmXYvNtjuevH6Tjc2zB3DkUW114K1
6YqnPQ0OnpZMwcKNXV2bAjbGsEOAdaKHKa3ZnUQ+pMhiSKl8I5RaS38KEkOfUKxD
8rZsSKs8ORjVCMJYB2IPrVW1wkoXOf1y4n5u1kNB+EovsEmJ+CuAfau41qA+FyN8
Z1F6Xt2iTbO3fMW50O4gVb808Nd3F0sGkC9ylhU2GNHqCsY4q1SFD/Gz7piuNWMr
L7uf0V93jy1oMZA3YmqgpfTt1HyXgYbkc501IuZ/P8WaYSp1IYDG1q+LcvsDohlL
c/Jw6Cmx2eMbormrMlp/4NnPUEwMvETpLMXfCPHsnOlOaXw9JlURUbXkaJacWZzE
xauJe7Kggew7f9/Kg9M8flQjaWhpb/4CtPhZYSDMDRlrzlmIwbt1eQbzS1Ercqy8
3HAoYrpPW0vczDPMYxtozXwtO+hN2/EuV1RVJw6tegdFrw16daMaI31KRqx28Z5v
r45JCx57I5N9mKjv+KjDm5+Uq2qqyFfsS6o2mZQaZcxrpCK0aAAj3uS2hH7g6MRd
8y4OB4A4suhNEYBEqHOOJJ6KwJ2hQx+LL3qMT3lKqtV3beicjBIMgxtbijAYX+cS
V7h7f14JxeKVqKej4tHtIoXXZQhbW21IE0tgXZJCIz9aHW7+LH+1q/XeerNKbQrh
UKuAaBP2JUT2KK9BsLdIgcq5k92KLYQ5CL7XLnC/Ha28QEevsL+rczTFS+yVliwd
cctl1qjaOxrFUTFgXcMkzswWTNXT2QsbZsoI6t/ID7zvT7L2KVnfXu8mT1Jrod08
821rq67bgMJCEA3sLPDl7C4fVA3uYZ1/z/bQjlRYK8L1wmu9sdKIT0gMDxGM6oYa
qKjGGTLF79NXnHcqgrAk2BqJ591pqhv5gRJAC9c6FbRC9nMf+CI2Crzro0ijnA57
6ndy62Ab4J1E3KyksjOE5tlINeyiTN43oHQ3wtv0uJK+pT3INookzeKYcIi91gvx
+McrI8rmp54ScQwjZwU2T7p7c2Zs/0Y44SaJ0nBl/TxVPM3dwNvltZUcEEGRIWMb
eGIUkfEu7FfuyMhJjphKuGCXaTUSRLnW6tV1F4mmc0VTnv7k8uOZNE7QV4vHPybt
HKsgtlMiC3UueQvHH/GXslGtCw4KU1z+myJhpI9zTC/mrdkgR12ZwLCwCDRXFekq
rM+1R1tA8yh2raP19jjCceTZPsnjBO3OqTO/+v/GUhozNS6wfUA6lLiScAol17Qe
J7SCJtft3u+9y+IWKcRd9K+a8ZQOzvPoA7YoPXHB+O4MiOfK39XVRuBdzFWGzDWU
oO1PLFasz4i/uWyZIjUMROe96cWZ7vGvx/WzUzZD1fbo9rof8JjIhVerDagmlQv/
e7vYfwX7hvuh7nVzmdzdjgmi0DMddsck6jin6D6+INv2ymdmoCjVJPL+J9gNpBFf
z02MyKfO/elhXJGoVLPNy2TMUc0x7EfpIzqUvubb5/hbnsWrRd2knbDcxkuxQXph
JyB4xK0pgCNys14CwWe6xBin8x1JYARMzQymeRnYWJJZCbJSlul+vVSa9RyRdYzD
waSATNWCwaGaTMOTnVXqHgsaGFEL9TzMLApMCitYKK00wrbaDPyazz3ZrP74jtse
RvF1lsADkqvewy97HgcZAVX0i8DhrvbOL7WnsVYwT305+p5M2zF1dpBa9FVug2ey
wVLvYd2N2HuY5FHH/DmIwbjON0O2XxLaM/UVCAQGdgPlyvZ5hopbObu8F3tcNwkI
xRsqQ0jxUVdtpXmVbhwTdCWNTonsUDNjeHqzPHDLsAOn43tqzNE/CGGyZIF3g0Vi
A+sE/Jj73fO23gw2/4DZcJ8Lnn87NtT8AkUGruv2mxKFDQcDgJTq062TLThVU2yp
lcQS9m/RGNmiZvwCChYu+oOYtJiJeuGBsS7VjyJRfW0dqNbwij/ORLJW1gi5UxK2
Y5Rn+AT2hgA7PnvlvwoVsja8w/OS69XDhyx9IAyHoIn7Shs4imVWi2cxV/UOQ6/N
c1o1iUgdEdv5Eie2frkppEtT9Rc31Mz4jtNyDzjebHTuPmlHMmICipQzwrfObT0H
AyxKmQR4RGsveE4fxC5vWR0rwaVd08DvbE2wJjFcSt3tFJFtxVYHCVjtFyyK0L+f
NeAnkJiXvL1xkzUs/CzUcnLP+CFwigrh+v3QWcZeDoVf+6Qdr0kR7Im0H2sAH9Eu
QyLwt/GLVNQ3K6L4nvhToGJOd0rMuzOpNVsD457NyQU0fFuIl+jIBI+mM2hVJt1j
DI3eXXrKCcUXHhuXZNNx0dGCh7OyBLC1mUd4OEpNwXTyQQN+iToYp17VhRxs3Fi6
iwTgVmZzFmXfTmHj1IVZpzP3H1IKAfqHFaHC2S65hgTVojtMtj2OLJK/4s9fhaFZ
eiOV4C/W9awOBGd6vroQV2J6LxQsVSS3aI/UWndW7q/Mcjyylx1wREIM7VNIf24+
I4F2K2LtBRS0uQMAHIA5Ykd8X7U/FRuDJGUkTBZgCJKx41EiWZCJQ1z0hR78kR+B
4tuWMMK9JB/wxcIUtSUOWxt4ZF39TBn8TszEgJEnSqyh/xt8n2by0H++Zl65vuAS
wAH/EJfjE+x9UkeZ16hHeI2U0rerinbwFH3U8DnV7UGaVuwo46U48tVjE1UON2jN
MV7iOEyFxKSdXMaHMvvAi7W/9deNHX7SbbcMFZhseUBilusXerogMH5bRxczFBRg
cFHiGleCtlPmBWZbFFwc7ApW2RMqXofxncG4b1Vi8oj9tkat1yv6+zVVPaa9roEb
ut/aOuVu9f7b51pXRADoZbf/C0Or9U4mqhKvB5clfcWh0km+DzRygxea1P5Whx2O
IoQc3oM67dLuI7RTg0d5v1qYiSE91ZI99k/qq87AziHALHLXTZhPVZy3+cblN4pt
Bgz8D/tUl4j33cKcUi0Sbe3ANXXrgF82dCHqHhQqt1oVdduYGWOCDFiNSZ1DNBKx
sbiFWLngL7kLk+wjvEKSL7IP6q1821sUpiDRolkXfSsVIWpCichI5u9lqEkUuvcU
qSdGEH3/KaS2RcZBq1FcdZl1FI7I0/seuKkeyE/5SmBMk5VSG5hwjekM4pt98HKz
62M1ChYrQrXgksqtqJrf087yPZZemzOLhbSiGCgGN5KHbTdQOAvF+wbB79IHWhJa
Wrq4PwoEMRibqugNcxyEYAqZ/GF8umbvUG+Iy32E8EIyEiaq1EabF6elzZluTtSe
oCgN7GGSMLm/TW/t7LzTxuqiF5JI9OG/OPPlPuFKXHrwgqeY4lp5ZhhUwtGAXQ6x
6FdOSvSAoBz04sra5nZ0R6/6fIRglGkFTXNGSouKZDX7kXVEdJF2YW8vu5QjcKJu
6zpvg9SAdfoKnosZ6Ir8tG3gXuNMkRJDoQuzmdY+88EEGTaXAaRBPocuszq1IS/4
voZXJSKuDvpsMYdQD9RCvEbCwmTKG6Q0Ss4VEytc+QOavFWiwfY8V/lyLySZb9fT
G8YCs479ELhIkEJjsAtjAFtOTD1NxYy/Cy3VIo4lVkLENXVMWzI8iu6XklJvfSbo
1kPo+/RAUgDwr+oIcjkQ+i6dQ/EK7wjj/OAt7Yjge8flrDnQilQ3Ac/s6ybf5cpL
UekvaEBbhIvmBL7yL0mJZ+oVee/VLWUrOLjT9JOZAPEc3BwOmvU0u7rhu+vsPzal
Gd9yce5xM/Bl6f/BTIQUUb66gG6nbm9e2HdJefYby70+XnEjZxRVhDzNt1cNSB0v
gt1vw8261v2/+Or3l6eH3eNkeE9Bd99lH3q58+uWOneSUD6eT5tgkuJk41aiKhuE
tkXZ5Z/hw4b9PAg9t5dI8IOEQo5CcB64yp2ctGoCDgzcTlpnWyUee1nSs4xg/THS
b96wWQM7i6kRDlnIIWiRYEdRA9zt6UXFWzN+C3Yk63+3rwBWUfh9DzvdEdRIQRbI
6s/KxL7kj4XrT8ApEbHbyrka12EbR76jgqy6lfv+G/SDprdxaUJeMO5FSBsctESt
8qMgvPT91UOiwEZNIM3kXQ/yGpKth6q4wIiIRb0z31SZQ4CUVUk4pLKDUVtsvW3Y
fRoI5vawdgLLBwsYa7gf0f/J3pYiFHpqIh0ZrFVFdomkor7sZo5/0ARNU0IuqnO0
7WjqAAdPamuG3HWVexyN2y9nYXpMyaRUmd3g011UhdN/SVCHXzc82q+PBgkxKc+H
DdCi4ur6ldmHOnZYomqIaAsWwzByJwRLepGEsIo6rr2aPv0OCGl/+LU0FLXVulBs
0s4q8Tn3C/sZoqLHXhDcviQtcRGvhYN1n3JrDQCcpvUwRy3LJAz+uQBxtqNax7tY
OhM6MzLVYa6JoTydSKaBCOH4x+njg6brtCqDK9J2eJlAFdlWeXEsNg3JdsCNClfv
5AP9qPMmF3yov+6PEMVRr6twuWxI7u0yql2gPsRQTDJKATmhjl7L3eIskWCvpqSY
UXnv4rMOpemzuqaKs/zg5sZtnZN84K8Md9Y+BTV3+W99kg8LU/rh6OD+4ChxROv2
JRjnFbVgK6A+XxU30d8ng91WFNuGQKgVp6VPfAMQgAOTE/BbomZHATb6ttzwjPEq
L72NZ49LaWC2zJjyhqCnET0D1Pxy0Hjp2al7adx4lYXcT9pxmO+tGewnnV515DNS
Y9WbEV3gYGTSCDgdKCBKiRTMexOFq+NHx0cq6RDBrqUfl1RLvxk1NEAIGVn4ryq0
irF5crojOrUBN1uKISWE/GZqVpYdISjL3zPmnD8JlFowIgkBqSDCjO+0T5CFb/W4
euhN/IY/PIcZJyAoiubN4uTG88fsUJpBqAkJOyVElFviC/hv+hTCEaxEPgUjR/uM
W2hqk3VnwhkRyZW+JCmq+XHYMhAbSc8gqoeOM/U5wqpd0F9Y1eYdA0usnZolqH1B
5LDMWrUOeUoQMbYr3D7dyEP87zvg2PreHClUwi7rYjDJ8d6KISP6FanluX2/khmL
zO3PSBOelvz0Xj5F9dls1A2qLTH8pT7ZBBAprc6Jij8tMRNW4i7xJGG8/E7aSlJ8
3WIo7bRn//dH04VmCO3iwPBv6V6Ua9H2ulrvV3yxHZ3dB030iqzl8HLYzEKxPE0Y
cOb4f50vnrHYclXjpjbQzQ/laxsJZLQeqp7+R09mzdh6sIsfq/2Xeeczb9gf0Ld6
FmF6vQELhOIxKRioPJbuw+DDkhE6Rsm7SQyfBeFiTOIHIFB0OwCYwW/Yzx0okDUb
FwE+IUCNWNiccYOgcIlf8TNxgMUjS+2ixa9NRnvf7QJtaceq7ZrEG0wg+Zu8nbpv
vp0ASRqbxa2FjuUlx3VO8grr+a1x8G8cwkYWERV1gRxqXBI+g9ngMxTnP+/Ko8E8
/Pgrz+t8PdiM08Tk3HqbaTdD/tYUvYiUaNIy/irzOVaEIBFLHNASWprsPRnU5jyR
gR6UpKqy/qOadCJ76MlF4WiRyCwmBYUDgNMsqxC+eh3ywlbLDMbh9sEbeHj+gmrf
RWJJJXXlbK5nCE2xubjQC4UCjHvmp5yy2ZC/rzkA8wCjiqFFFKmVSi+0dpsF9oa2
9gKw89my7NlvbOGs3MM0BTbzxNJy11lvZJ8Mr47xdi3s+Muw+oPxNNfTM/GOvlgQ
P/FOS2CpW5H0YdRzjC7tfLcHBZRTSSUx98NMu87Z1rfVL5u6Mu99l+QTweaZrIKo
8YPhWx80E7C1UrYQEPtQaYXseC5wVli1WNwYmdDXykWENFcsJ8K2wiR2m65Y08Z2
bj0esKQIGzDClSsp80QkVAAgKMtRqE5XxWt16PGXfa64Qnu6pmG5y508O6gZhXOs
2t+Xx4iUEL86AsYT8+iTaGLjWSOkOzdckE3TTcJpqU12n1KkTwPaLzj9vYP/3oPd
rCpyRvJUQmhOCEQqGZ+BD6zhbQajDTHMJScHPsiDXF1sg5vSNCT1XAgDyM3DWROK
U3aFENXW+LxdGeDCPolblXUHlWmxzZEsh8rSLF4XAI3XEbtx4yzXIyKP+sh8KlCh
0P8zvWRGS6THdwOoziqvf26vE+gt2HRnPK9Vv+qtCyntygpS/4/rc01ROTvj3VPu
CI36fyCqfADsWFSRoqluopaZoQttpixNizce1YBmu28jGfMOqG/IpWHryAMmc1Px
VYzEzM80RTia3D4Uxg8QfwsLVcJZHN/otmoazNeLv4uPolTxRbtUCwsbyI0Lj9bg
8Bs/fEa1lKx+1gPgRxFN1o4kbIc63t2wL+wpXkroOnyJwmF3fc7VNq2BUW7Fg+jn
/6l6DDRDM5H6lNkR+IcDnGg4t3M414QzSYVFxRfyzNMS/zXfVq3XohD/DRy2H7T0
bMH243UG6pQj/4oCBNfgtHzJTORKRgppOUt/zLyu4bpNIj4kD59OvtrMFTLtgoYY
DyQuTgD3lLZtdeez1F9NepE+cHGjdarSqUdfUUDGDCfum7X4kOZIBz2a+pWroW/D
2EJqbEqw43KQ+Pq/5Ual8liQ3UMFsa+4NTGjz9xjV7LOglCpNNgxwYXPV95zyeiJ
zxKcniCF9GZ0emQotaJk6z8BFWGUcIFNHAxLUyOD+LVohhAR7xs6wlSIiQF7xVi0
ShNL36n9wxBuQsddA2cOfUQZCjjBoYeBYcJ0APKILI3JSOviSNklv2Xx8ddL6BS7
12EwOqJosSw6F2c7dNHjHbtc55PBoh5Ah4dZ4SFbGbXJHu+iIt9zUgzCbes1YPzt
4lMtJ+kotDwB3SBD8LEoeqdSDxC8jThYmA3VPPeomVN4+5UIiMfwTp9F3vKiMfUs
7e1T5dus4W/s45O0TSZcjEEu7kUxM3UgXQDsujtETThUL8PfBgrUhvODtmjmvo4y
XS0yhqlFGz0QrJ8DLcoxcZM2UVJfXY5wFQfFXNLNSouXyVJ2BO3MX8B0NBL6V79c
/+VqoiA4/sfL2MVa/lkhqY7Bt9gfO4lQLBcghvNVbes/cyUMSQZfjTTLiX0rcGzJ
SJFKqrd2wotI6lQRS5Gu2Eax5VMGD94GoRFr4TZI0XjxRE8M7SRQElNOTh11T1HW
BUqp3zGPp+IePY3pWbUBXDjeiqFO50rx+uKQ1xiDUZYP2h6jhAcKcTUaoZm+9EBx
W/4zcNWFUGXZCw68U1ceEd87bj3Et+s5RXF22zy746V1mkDvqWMzEV1KQ5INAryn
pV6dlEO9shF/sOBgW9aueVyZ2xdE32HcnwNkZ3sCjjwWy0j4tRywHGMu24di1ImI
yOQnnlyg+P9e+ACPHHfhuSa0EUxoVZZgJ82Sdp4iX+lvwqyE5tTjcZ1y+clh7uZD
X4OkGFTFAPdqkEqDVzA1/BsXSDJb3YGUjz2T7Ewu8D7DUzu/7TKq+UCKK3C3Bir9
TIkPLQhtuTGsPewH0tzts54XP0tPeG0SVXnPuZKz1PdENTnOyVGB8LJqoNBoIkBf
rJE9uXm7RO9Gjk6EQuObhClgARQgfccrJGOuzQjJueWOwtjvdASKwhRD9kT3u+wX
NgKkFgk1Uv2UfDUbXIn/nEpdI0Mtce4cdw1Tv+uwY0+wTdgSZ9MZw1ZPXP5udbTQ
Hjf6D5fVC/3CloBAP/7ey+JVHfNUQTuuCCsdFH514MOdIF5oisd3npzkEn/gBOaD
lExDxfrwreolMdLLCTcSyX0AJvuTuMc8gF6ymdcS+X6xuiJoUISnNnFQCDawjJBf
HdGJNodz4YRcahy6Tm+0yswGF16RDxx9DXYa5huDuna8bgih+91qpW/NkDzx6eQZ
WMnlmpezoDVWT8buUMAzeaLJWdJNJn01W0lixh0P6sRmsYfpWpVZo2rWiPwfH0ip
1+Uz5fAnDjX/sIMw+kg9B6c5nYXPcnKREcMHR2ElUjEPRRKqQwDEK2LUQWx6Bypm
luUQzSHXKuZx4odNMDmozv4XVbnXVXmgNenIFOKufJt0bLqYvbJizlYN2hCL+S1k
OvOvdjDQBVpIbICju0Qf7JzUoOn0h9LmDsPaAVaIHAcI7m7lsT0x6ayT70oqr6EA
z0nO9ie2OvyiHusLypaNw3ggADnHbWPXQ9O+yEZiwlJCjGHCrpFdWeOlDioQgk09
Mt8WueZkMSS/pj6pESbg3PbQ5yvNMkpA3/M3QOVjQoBSF3IyGYY2ATbaiY8WsdRV
2CPJcVIGqVKHNjV4QQm2abIsicMyKEho93jxA1Q27KGjdIlNyRnopAc2kVtRVdn7
CErs0vedTFR/Lv+2hD0XscFbE3eqL//H1yeELfQ9aTkAvcmrlIl6X4uHFOordbLu
Za8bmRS6Y6Uivy7aJ1ZKQqrNGTznZlPnlNLQ2M+u9XZ2Fkv8OFptZV87CIUYLsBj
cxtaomvisaT5RgDzy/Hw3lXbBcfbHvcLec6uIofgRTB7le4aUQLz4R4u70L+IlLy
MwxWb8dEMla4+V/oTr8tQ0benQHm73CNGHUTp0/c9AwNDOpPEe6wsUKV5WyFKFB1
lPqi/UrLY1a04L9Ym0nP6ujFPbGlTYoibYYdUJhpxzHUnwiJwA5txWSZitDXoGWV
bgEBK/+SsS0SuBy2lMAoMQUsJvF6oHXOjeDRq7a3slykN0+z8mIrZQqKtv62LuS+
1S4oAJs5n8z3mQQggeLHsbZiBecUf6ElAn3fvJE0gNc+J5J0C5w/UZndbOvEZe0d
S4sP4gnGrXhwqcIolb2q6PvL+OpATl3vh8avS9BaAvkVBWijhaBuFvpRakYhbgn8
HY0bkckUMcT+IQuJMEn/Ane5WNGbFiDvj/uWJkWvz+l1nR6sQEU7JOd1OcAHlZP6
3WRz4wLoKlVlqlmjugD8cfngWG/z9mipJdMlwOOSKpWpnPyTEGdFqriSFUrvDF0J
aOvaxEShyXTbCFl4Ut8E8yvOG0op19V6ZPhNUsxtWt3G6RZBDaoQMgHzKLwzhV2S
TnJvJICexXx5wuEEzUkP4rrMxVhr3KrK8XLj4fgrlfYWGqScE9PHCHZpOBL8q1d/
1sItvpnN6ksIk5cHpXXkL/+YuIpVHXZGXMhT9LCU4isxv6ToNTRAvVSAeWioGrhg
QrgjJQRe6pY9jm40zs92a0oedydLpjwOfD4HTjkypyMnC70J6lIdr9kesHBhFIfq
QUXrI204fJ/RGonJkZh0p/iXxyD+4yJcaDT1IRT+59mdxorwm94QR2ACpInp9K+4
aFmpK2nFw1DUvp05UGN1jk0D2kbg1Y6/bu2QTgq5zrz/GhsLObpG7EX5llLtYhr6
289CpbtLomo63+SJIML7+NjHoZ/ER6rv4qhbrUY71aHu/Fet0wSvqHiv9aG74J0p
bw9VIY5QhIEeYxu8iCdOXT9LF/Q4eTdJ1OQwv0O71BJvh1cGpFWZQ627H923bpXO
TsjSBJrLgVutznFDuUokGJ5zG8BR8WgDN+65ZKgdWS6wM2LTybxvN8jYefvAuUTy
VIZ2T0lMgaDvLs+nThEyC/deeFnSVcA/2tP2ZoDYjPlgrlhW+t3l6/852wfzmFuq
PgkhypuLIz7yQ1/ejEBWqDs/OR3hdIXU4YX4us8xv+kYyqQ9gn2N1i9GzFpMVpuY
uMgjwDmnJnzOF1zWPuXcD0rLQ9wt89reqdVJF5ab1nL5BAX3QAlhcWvcfQEDgBRz
qLhPqlQKDSfoZI4dCw/kCKUb5hGdUntnmFootOca9dY82JJ1TioFau/csappUkgK
xz8/XqY8EamVd+hVLq6MriJKQaUyBrle7FIGJG4bD55VekktX8kjirZi9+2FYLFC
G64tu7pvbmPO0OMPEAkvl/ZztfGj+denzhBnhLiJD7qlb7yLuEG8XLt5LGS8aHbM
7IoliMdRWukoTfX/biNM87S6fYklx8PIXdR3QM82oP0TyBSv+KSkQF/UXk+TfwBW
d+sqdpu2j+e7RYwqsilok/iMKhqifwdI3b/WrZybtfsROIEFqVY4ujMfe2zN33J/
bjUus2GP3EDykcxUTah8hCWrwcJcqC74qHo5Vcg5c1Ebvtf4nHsX4ENJy8Y08tdm
V2YzgqXzbEvgVPGcbGOajhZL/81syx8kEqO/rMDCk9RWK9I4cG5ypZ/mmE+orNwK
LEqlrDtWMUXU6n3LiyRbqDSWzxCuYhRs1sM2uo7l7srr8azJ4z4dlJRkhjtHt0Qx
SHvjkFUbmxLCusMX8mV4qvU53VeB67vWKlcmGhzvGzALsTGHa1XNzvd8gEbwyQll
80pfrs519ZjayBaABBvsOIpHVMUTXaP3mqmoESGz1t6AtpBD0ekE2KY6ohLguWwE
LlANDv6hS5MjYzNTEL//OQ7qSiAa6Fgsa3fv/qBM44YQdnd5PYqo+HXcWpcLdTB8
XeCFB7jyRNAbYiWzk6Ua38aRcqz9q9MvCTzVuxFd8/wsTzspjdKl473FbIKumeN2
ug86K1a+F/DvwmiZhSY8csHO62aUMxoXy8fZBEuXOEEZZKgO9iYJyGjF92NiOTn3
EBCz1zBZvnqgZCVfuRgT96610VSjqe7NSrEQUbZRpcejKOd0Za3Ws4nrBcKsdDbS
giBSOTJbFuUy8bUgyOKPPPmSS6rIes+V8Evv1NOd3huEZtXQ4f6cBRJJisIs5JxW
+J9CmWmv1oaItjK/Wf3f83hCCFzip0CksUFZkgN33PV6bM397bXQm/SWTcerA87w
GW+1nOPFvzAYKl6hY6xE7nyzqfTY6PyuVOAWFSiC15pfXO5hmyAGLPUX6SbTfOEi
GByi6qYn1SAasP7ZaI8PvZP1WcB8vVTXiv1AxFPktaSWs6NCYLmEFanBpFo70J5m
Zs+SYyQR0vvFkfJUIzlipy4SwMFPT5b6o6tCdNSajXEJF8t5g6JT/ITHzbt1hDdP
aee0kaB5tJws4LGgnnvz9DqV1TFDmtbrTxdESAsiEG8AtuNGbpQ2IGsC2gaapbjI
e9kPygt6hTURdKslnD1aC+Rfi0ostOTOBRikouV2V+FraygdwBkhTxgV4BiVmNSe
vv/S5qVhOMAzZn0GklS8xVvZqvExl5324mAHO1Nd17CBRB6CXwjh1SqR+CFtTf1K
7M+0PXHI4ubBcFcdB30nD3FLi88VysvK1MRrLrq/fXIYN/iaVlgZoq2EwpOKeUyP
xQByg8Itj3FPQNyv7Zqj18cXbMDguzUoy/zqk6RiYw8B4RbINTvdPnf4PE6DTZ1W
2Eu6HFDrGEkh/l6SxMJSF75deAOZ+lxXn1ddZXuimniQZt6NR2pEmdeo9YCRIBae
Tr7iF0lfyy64TP1xH6gH1zEG79uIrUTcO4u11xxViek074s2UTrcMFuP7oMsiGFl
o21ygIrBaMNdO+UDyP5b7qKRtYQIrfK/1QKBoSK34uKIiG0NFgZr+h7skiI9eQs9
58HaBozq8KwgwkNJBgpnNrJdYc1KCZEGtGSX0yIT2U1gobzQ7nz1qULoEWTcY429
3ixD0zfVGuYHM4wOPtZ2/RMXgvTJ3KK0OporH3nWmUE5urtiY2fXyyKfHZ9Wd1gN
m73z9dtqCZWYu3oT91RCmsUXSo9MAjfQgb1tHKL/R4RGvqAHZRjcvJonwXDCEdXN
N7XYknfnojUOgdCAEW008trZM9ReMloN7ucVINKAlldCPC8/j4MHGT+voIzE3G4L
oNdQt2kTiGAPWQN3oRKO4i11FRYIgIKll0wgZCbQvKNHqBCaDiO60+HxcNMmg4uu
qz+PdYOZwl8T/bWN21298TsykHsF+STqlHZ6gb72fB3ionI6eMg2vZcgc6lhNFOL
HuxdX/ZK0qqeK1L+tjCQvTjfvUyBbm7XaYYEmIih4BHOK1U58xM98S8rP6Ago82H
C7f36AUSoZ1o+8ebXKFvI44jeLVOQWoUUmZ8h4xiao91t1xDq/o25aOtr1FT044h
dNzVH1PS9X4JSGZDQG+KEVoOOp9q6hCOFtH2GjdzJ9xbn1DRW1nbT3nNyYMYNjcB
RKcVIo9yV5bR8MmteyVxqDGnvdLZNU0CkTN6dWLf7/BUMWlXWd+tKMDguAIrqu8a
d+qVpGHXxXrxdTVAuomahwPW47yzlxT6qaK511m+5gXOLPYBSjwukvryjcQrI3Fq
6fl8lu7yvMPwz4wQ/fUsSu3G8m5Ea0LEGKGpMorvHlZFpDHu8FCYMErSca/ned/p
UyXtEVEPBmEcI/TNb1+HXvPCFAk8KbOf8rv6wby2guR1+wDoqbwM+5ka7kW53h84
MANX8ESzB0zuOK0sbIwYjq2PBCCkXXN8UDZK7FGHpLksjm8SK00TNqnwBWENXcfT
fmw4L3cB8pKDxYN3HAQl1fu8xZFzOtZD8CDfS17qWgGYeCnskCURsf+X8JUN05yO
TOpSzZ2BiLGudZILwZmK/Hx9y99qdkT/uCMKNoZaWOvXhtsK+7tI+oSg4moiyTns
dAkRiZ9kX3x7FNpLoIaZ9VL1hRvuiCfPMkEspnHCR2bR02Y3HboENE+X/S/XBNLN
rS9PjZbNxDtGSJ7jwsAwAfS6hSN5MSGvEejpIaH4Gq8c8TjLtjaBhoDd/8CJcgsU
8HpJGWfN72Rq4hqI4jH7mHnD+WNGNXpGS0ZPhfCAITteIqPqqO7zGJvlG3Se0O2T
eEZ6ncc1sUs4myyKwxO0vFnbzCXbHOT03+7/EbKBMIF+pd9EVmI4lQS8X+ZG7kol
kR6DC454QDFC933Jb38owj22iuqcomFLcdagBVWYTeGnit05wWTRbF9QxV84IjQx
6cYktgqnNnrXKxZgZtuImjnNbctcAgN9PeOyXiaaUN0F2ROUK1ajxU/tXiZSKYVO
n7r2ldmu4pP2gXwlt1utMJ84MfNg6gNZXqyPWz0VjOhtdBKkEG6zTfirAJZj65R5
yg7j9cShKy7PCM2FfaNm56P77Dtc+8NUmriL7FrbTcIfq2FMquePn6PdSe+jjARU
pON8L6D0e89Uwn7uP9R201JXRcabIOcfP1SnejIGfHUsPoJ8SF0r0V9bgN/NmwFg
QYAoVTtP/wAOe7Him/3MksW8rtc6VGz7E2vPT9ZecydCkarAdzDTc5+KHYA/cWAY
Dmwy1lKeW3FG2sybG9aU+NOqVGBYTG8FOHQcPBOwVA4QhiQdfwrILHYSv4QY+HCt
sSjVzB1OvqdUp9Tm9PqXY+BihwotdJIERReKW12TfbKF/l2OStEe3GqQ23LdMSLP
GLsabBltaIV5m/Z7R6v0SS1Hh9ESCnZKMipDq+QE7BQpLrOWXvu8sjL25TG16q01
Oyspq/WitXUaVywKtCQWauXGAYlQOOJFeLFmvyaYwu9EcwKeEUWN8ovL45ZfRhNP
TW2Ne0H1zIr6VSHDunLk1UQ/6JrVZKoFsD+Gh9B8qk2AWdsMNjUZqyoBcx8KCcHo
2wEnU3V3b366BEU31fWaIFfABWIWc5HeHmF1JANQ9Rzbu1+yGc/V9pCmaDY+x1r8
XTisTIHVhJ0y8uUr6elq70flB2WpxirF7IMrFowTQXlbQ90nTNxpZNmVU9TgvIFk
Yp0eTiYaqB2z/WJTHZ3D9Y9BOsm6LheaYyStX1CwXb8VHsI+IHpnI18M5x6FbCYG
qEiTwrAR5/yNCUJOp5AO3LwYvjsdeAi+v4VoWvyQTWPvFvQiZ4YXwLPZ0bGRwApV
mhEFgSRQlS+hNkIuSt6Zzga6LwUYx6KGoVbFQe3f8Q9XNo3JP27yC2yg+9LGS1vw
kO9WTBbtn1vlvGwUri/gycQbeHFH7bRN8kaTfvGa9Kg0ytrZxOLySQZtXO06Rtgx
lfKDZuNphiZhSLJEisTJUkkrQkQ2kbmlDDWZySXcgQpkcny/Qa0dVmlcaPyUrnrC
ypbQghRTaR7JpypE7hdZpcya5YFLIFheyYEC1s7ktYeeviqmyk/n5/JOP6qvjCxi
WMW8Iaf5+wQKnUONMTGmPFj553/aZc7V06s3HCbuCUx4VxUvzNyH7z/WXWRovFvN
8uPbsclv0+h3/otNMuMO/4h6VSC+cER1fuIFyKMIrXvKOUC2C/JQVOSWIjlF8hHb
ybk6gre2fpIXjMwzamG4u5GIJ6y0anlfu4eAPlSWKrBTVvsnuxL/HRIIRvbty8k2
JN81RzgvRVrUzAA81IorWcayLx0nQ0tc1GA/A/xWenjg3M0S5+C/HGvseQxaVetD
d1V9O0t7gD0U9qMdjoaL7vIeoJdQDSWbUnZAUEpJEpg26xaucFU8YdQKKt5JRciM
tQoASX78z80aDMpukslFPoj7xkMccGTvNQguPg2Pkrb6IyX9Ul4ZvHwo6Ys3Q34k
KT2Wlzdo+XssEqXsMXcnDuo3iVf6/gsA4Jes4GFeUjD3vUhivR4dqVfc5wwkWw6p
CkHDV61e9FuzEH85C3QmeKDUgf17VZHLQbM5ehEdEAVAY+YQ0vCQYHbi1fPzTkQT
W35UUBuom4Az2z6WljmU4mp0AdkeqBr1D2CRo9tGDRyssHWsW/GmEmfSoW6dAVkx
I2lx8Y0IY9QKTLeyT6AvVJ49fApy8Jg4P5Xlw4OdlHMrT5WRDXjBIQGdraCOCfnK
yex5Zq4kNezsUIVKhW+qL4BJPZBRPOnexfQk8NfYYQo3ylb/7UkvtY9ee8DonjG5
yThLT4aNn7Gmi9P6zMSMDqlohFEQnavaPKgYVzB/epEkUIvXsycU/cqgY/pb8rzb
AH1KFpANxRuRNO6UzuYVs2SPwHnVrWOQ3kksC9284gfYVJ5ft1RPg1rb5pww0BOA
filylg8+8XfT4SN3sttMvownRTRTztC4+4lOaneGdPbpJo5NzTbQ+q6sVWmf+Hmo
ZMHHJDW31B48J0Tmr9MIV0VnXVw57vLTIQSqCfWh3WBvMyLdrXBuIkZom60JZmRN
N8C+/7SETTvRXP8W1r9NcsjZloe3p37Q+7Roooz8lb3Rv6h46VpcF6GBJwHs1H6p
u0SZh3GW8CC6M/eO79xrG94607PCJA2AwstUjxPUymM/Qbu1ChXCcfDg4TepC3iR
UaGEDkYOLuqYk+N8+70so5zURmDOHEEjK/ASJFvCasBjskwQVasKdw84oRQphpYN
18Wm4LRaok/k8k41cBZpG2hwCtjm/22rGbPcqNgHqOWa0N+m+gkVzs/DjKzZkLxX
0b/xZKgGzNmhKCwNtFvfw9W0e0n4CJsiMAC/nmKDXjyOJ+k59r0JxtQa98vuKgAX
UxheW0xjwnXirBqXVPPTNA9BI8e5Ej1EyqaD5jFvFDO0JMlRHAIZ/jc9lTzr0LDq
FobzoP5PdXY9COrKzUSaabOefoTl76nCIsHd0itQks1aGvRzquMy7OBIq67klZmq
/EUWeYtFj/wJ5X2y3efxr4+xBBxH+Hg6hv3nZ5kPKqJJeNzRsviaqi0D9DVjZQzJ
S6MLR7ipbDuYFlgsd10G3VDDGF4eR6vUfiwkJY3ojW8zRa4/P0rMOw29Fhfy8CIk
0U7AJSJDYlPt2IFNV1he6VCC982zwAwgXnSj617mE1M0xl3vG4GAdVL4y4M/k07T
EL8du+5GtF3V5tawpNKYVAkAeSnZNa0wjA0xR7KkRAJ44I4F63g5Qhrlr9chEBCY
ENPNaVNpPypi7i7VN74ocvnaTRRgMj7hCGN9y9RhwSSyVs0HE4nBChZWhebEVIqL
zgfQ0gFQvRJx5VFhJKX0DKjty+7LKrkmdo7zQ1VqnISZnHT/MQqTHkvDnPRIBEd0
029makjZVOQHEUmj2Umaxvc2EJI2YwUvpf2i8VqoiD+VhF8DPqD5xIZ+i0mcn8Sc
Kaf0s599IuzMsQb1+RQkUDK5A7ODn2QJ28zwOIqa+/eU1KjOqh9f+fssoDUGo1Ct
AuAqJklb9s50cwL/diNQamF9pXdJLt53uhl63ppkXBULL/RlQPGB5ssKZHGCiOSF
WsfAhnVlqzFIvQG8hYLASBue8R+2cp9FaqPz1kOAO1jN0K5gXi89GXVbI067ucp6
gGgvC0RTdrLQOEMkNXHWgH96JPbNSY7W0fWpzlnKX3GW5JaGYNwf2Z3wNjRX1d1z
VOhQ4/pRa5XMrcs72O7SrwD54XLgZZg1lFNL7S7cKFc+y2ySbo03zCPzUSb6E5Ru
+/5Cd5KRU55qts3rfF0OICPKJvuYnJHw7cfkaVfR5ycezrsq68CRrVrPdRbzMyVC
zYsRX9gwUuowKwgzn/9jds3gJtvdQ19Dg5e7eaQ3u2nPM19MdOvn+mVWWvDjeJ/D
gJB7FePNh9ZTyPNPlsGmDgjDf+57mfvdAzDgWvKM4Weqb0ZhNOjd+fA75H3gQctt
EegigrIkNTZxGHL5APONqzGcePjrUn1Vs3JuWkngUqKnM6+m5gtZbql7wHgqC3Zz
WwzPUkDCyD1Y82k9M+qAAwVjZ19zq9IlTUCC+TFVHCPiclGKf7PeFKI8174nAqEL
p3BfdFPFAuNY3/opWzYHpHC1KS86EEWez8YqfmljzmkINacKzvFZZ1Kwg4aYf9yq
AI0VUb5XzyM/yxgtw+gyCWzNTCc5TO8GS2UiOatBFzw/SF7uKklIPP6HMgBGdLId
/t95qHTyPfmMHh6FlpgT+Uwfg7l8RDhpZ+reUPk6dJLIqjQ4vXRBcKpj0ogQZqcg
wcMDB1XAPHD/IF3/nbFhPjX+BYt6arMXWtJ5uSHXSXbBn5GP9OLo/jEQd5y88Vd2
pVc9oono6KcipV4/3oYTV5KCUTEnhAcrMv1J4a8eiIX1gXmm4h5sTbbIll885W/V
zX7zKZslBdbGKVT+9cG0Vpih8hHHykzLVAn8nhpR0e6R3aloZZEys5iHuxgkZrk2
zqWkducz/3o9sV2TsOSyyrW3AVNeSmPHKSpK3K0lYb4Mj8qu2gsLWCDMYDYGMli7
5cbVbzilsnOyWmUj/2eladVQsIxTnzeTTtPIq6o5uQs0y+ow1YDN4NRGVcKbuTPC
Bda6RzPqJm5345wlWKNxy1cs2qd7Uqu55y06BxxYO8JN9DdK+VUn2o+VEKtYL3Z5
qSEC6i8a/AGC5SRzCO6il+ZGZzOwLwl7o2HCEIWhVDhnYpSyM3NqeAXEFuvK+7le
8M6cjup/iKiDbaWyZCOFf9JjRL7R2rXuME2WUAWmDIAYg1edNyvVEw2s61xQL8Mk
FcVFeEclgcAyxVe11HFX9WVrlQlmKsDbPqoKNjkt2G8tYT/du9eDWvRFA1plM0JN
u23fxWPQr6bRPwb8YmEMevraAdnpIGyDdoA/emf4DRoHBfvUj2UHEUgUVfYIpZDt
p7Hl4WVdx+mNuL3USDV6csmDL8fFV9tJ8/1i2IKb2SoC0iJp2qwgK1rIjly/o//G
cKV3tIwGwLOaAoh2lzbOoeQpiLz5+BuSMO7x7nwIZ6uifMI2QWRttphF2SY8CFMV
eNUhh9mWV7l6QSQ6iTifqHo70/u2u3/jHNjXQMJu5aHpEGh3XO3P6JHEqzS3K9tA
W8vW7hPYtqmm+n4tI78TH67dGm/Cdq0LhykOfV/DwzrZu8hHJlKXdKvkCUIGQAR4
L0eLxApc4MmgElgkxOrb09mhsj7nTm4Mq2dwtRXOHqZ4Gf+ArsgNAB0HNJHfaqyf
9WDBsuHDMRe0Nv5qdVaE34dTVgUPrEdeqesLF9Il4zmr+tEvUpJDu5kK9IL4NL6v
Q/ThOO3WPZyXyBL4qUkewgJqbwUs1LWXGClGkwCYDaJgDXl9bIYoTzo+6tFh9agw
3WpiGPJ8rebaIcvzaSTbpMi/Af1wVryIPmwxnaVOdcV8+uQ5N9LW5Gt3xv6mETiv
G4IJJGJB3R/BzwI9rhYm0tjMGmCPkNA1X/KjukOSXhBdxtVfExwmjc1Ar04k26o2
gLzc575MTgSFKpiU228qLhFUGFK+vhhTh+sPGtsmzkW3UrT9HC89unhL/7Are0lw
ieVRpMkiQDQGwfC+3V7GcR4Il2dyV2zGMHXfG3EHKt6KoUNQW35FHxE3uIMIDlI2
GGtYKqaGttBdb58pqhHjrd5kw+gYieS4uCrdSOiXVoCrJGJzcis/JXjANg0/ZsaI
Hucdqv0wJwE0yYo8ZHy4TMou4TSUqWbbDlAGU/ZWXTkytCP5ChAYUXdvYlQAx32l
68tPjeKrG3pHcorefZ+IgQP5eHt3UYEzQo1F2xLTO95pwj+kvygjFPc39m4+VWUQ
6rEjWGOSrPCyPk49jBWJByjpDp9BdZJjX7q7CFLmq+/2X+bYYINmLU2Iq7c3Xnwz
lTJNUKS/PBG8V8LSOOn7s1cFj4VPHbl5eCuRjQv/viQrVAk0fgeaGMMoNZ7sxCk/
kOIHv4vaPZji1I2MTrTBGYzKAWWW0+1kokOE0eU4McUB6Gh2it7kMMyncaRVLc+k
QFT1Mvt8rINmM4/MBR/qEPardJEO0aZi3qY1CIEHZpizUxIw4F3stqf64+BglAfc
wdqqxgj2h6dV28xk/yL9rBIZEmhJlyoiNUdqQJqu2TjuyWlMu8lLz8qPV4Cr5C3L
82pm2q9RhRiKR94UZjNo5Pn39wnI2k/Fy6Kepi9MaM7gI+C/3cqPxNxZ4CC6laFp
utUXn7jaxVF34ifAARj4U4SHWacUtc2J+LgwI+ZeWQnhvYaZcV0kjla8DwvCnMKY
xE7GujwlRwK7robR1tz/8T0G8CPb5yHQkAomVD2iLAdfz2feQfPPtx0Pm4K16ddq
PuQO9z8H8ZDtUve7bftHHkmWhbCUJfraQaDJ/4VANK7VJtgFNk8kKhTbtPTENVMJ
rB336AXG2Dh7Hqpf5grkWI+ru1dVgdfrqkUvbL0PMKc+SsEE+bf57p/E8WWPC49M
TvdeOyDeOfujXpuO3pj83BPG8hfC4e2SgDj+IAqdxEM9DFQqJIbqb4LqSZGCekVD
WKCsGdMRfQ5tNwLmbwSzuJK+1cM4uaH7BbrN6rqrQEMPvu+KnuDLHkiO5wOxsk29
hkay/4ixfP7xwurPStIYz+niN7pnheqJYVARbFjJAO7nOPUW0jvVFarSaXJAqrcJ
dtrRehWUk4c6YofnvFEa6kMhkhQPx3gIDZMIV14rXPDeDEWYNhgO0TyIASIGjCGE
Xbo6gbJxE1hRpbgR5HkQQlBGBJ5n0AAr2/WBdLPsoRRDCgarXvgcAniYrO3x4imC
yimNMjD3LFkcULyFVyAnU2HMBCTx+zMCCp+M1LM7mS3heseKgPmepaeTk5PqQK4s
9JftPd4qcTSIW3IVcqc/J639UCDYyEFZ6kad+T9348p/5TDD7WBAKXngmCCzCTTU
c9BhPEnLKe4w/JVx5TGvGfepXnbTwGTd6SN0su/r4E3IB31Wd9mmgEy6q9mvGl8o
1kHlYRpsOU19f/kJGO/QJTTYHCvTb3HjoDceBk9YHy43FYwDIwNVQiwAZ+vkISzr
GubM/aHBQWiL+3qw0/M6Er0pPqGwPikIC7ocC0XF//7zRFUhjShESK461/3Lx4ys
GDDLI1TGMU3FNb8Cb7IOKreUVcXlZJXo7u+L06IVK8QjEuo6qypAVx/ub8loD6XV
hw4QpXvJsJj/BZak4EPFBT1Ty7TkGlcyxfs2XDNav7NrNSg4lawiZzgajlXYJA8L
Xc64f9xsQ2rNfJA0FI+cy+e7hXu0GQQ511BHIwAcGwVvoXaHvmWSL0H4lWqmMhaQ
C1FyyQ9Px4kgp6Rs7LVk4fBjyC+8pjeAadditMxmUoiR+uoj4ReFSunL6G870AhS
8bYy7OwrWMfvgUGYTqLmlx56V4n+KZ3UVHY560LCDUWnTg27xlrXzSExNoc0URaq
ptWwM+JyCeyqQ5NJ66e9qiwka2UYGKLsAXWZxUev8NV2EQ2WBdS5LDzwatalpRqb
nIth6Q8xdcV7fuheOgaWcFJIlUoC54yEr4CS3YaPQ6iMgQZ7jb/N/J8rdkqAUPoZ
dLAotwivf/E6mR+5Ao0BbosOvtlSFfdWtyar+N2pyaBGn5r/fhcINN7Fez7zbnPX
+3ImcM2pglcFDICaxQjZYTY6IOGbdc1T8eSZGOwy9M+dR3H1pWYHD5i5BgYpV3nq
87dFth47GTNbh+z86DJJbwAPL17JKmkbB+FSG27UXAksWtju/waS20E+6uv5C1/e
sPrpGg3MalCBmnUc7EhoxlruMOZjSrBaYOKxgpXgNGJ2OT48zoB1spLTT13x4UY/
7+MZVQ4hymb/SIXynNZ+eGRj2T8b8M2qrNrvk5AIY/8JBFtQbfzEJVhcYql2PWVq
gwf2v/Qq7dfZGmtv239X8sCRSFDxlKLU5H6d/EHtjsNDkIky9n9Cbo3x2lwb+vb1
BcAlI2SsAR/QpBXTs+OcGw+Q8hjRxzuKFnXdfUZ3qIaUFvnD5wfXuXlY9fpb9nFP
CVALE6H4SoNzLh9fnpRJb9gXxwmpYDK3Zwj9D3wPK827baggZRm/sfXs7OfopZjj
RrVhs13wy9PDGNDxos6BX8mfNOa/WFtw2VfMlosGhxYb5gO5L8IgJCTKhf2DxCf1
awPvetCv4qZaQxQ1hGpUoBIg/3fRm1H0Zka1NdHTmQ4Fgj6pmslX35xWFrYvFpzp
jwhtel4C5NTuuWUbvxgwhOOajFcqGNeYRc6hNgxLycIJtyVLW+WIWWVmspBSMG1W
M/kImkVnfPtWL497HLQjSEj7wkLHqlk633R+J1LFGBdH0rCiQ64L3RBf/jw5XouU
VJhrtkdE3HgUONwyBoKdqkYlWY9sAXq5l80tffbk8fnmYBLWTmggVKMcDcdfmgJV
Z+Fksc392fojG0Ixktwtqqvj7+pB9VjOV+D2E1J7TLBzX2roqc1lb8EMwLQu8T9e
relJEUF3qtKZ9PrT/B+8eri4QuHOuRdolavt1d00LcCDGuzwEao1Gp/OsUWSxaks
hm9vcMXUDn1ZOirGKwTPathBACpp5synYa4884rMdWvUhjHkXAjAZWOjlwtmOIso
bZ0epIm9TchHzVG2nMpxbBqa8qnheqsb5P+Krh/xmzJdAkG+GCkWUnPBkXgfynYA
JhhK1b2RpLMrHBYL3B2Q5hOBqRcxwarsGGxk9rThlI6VwuVhj+9GjLmET5SexfLr
vYFqqQg64z88/tqP8GCeMNRQF0SBbxa2j2b8Y87z7AEeGTxkvdLkzepL0pXgXMz7
UE1YBDI0ubh8X/wub5f8ushu1LlHmFtj7dCCABhbsgKOY0O1nMbQ2w1UWzkmbYfg
7ZIz/d8IY8F0k8EoCJUEYBqQ4DJ419/Dxu1YlwcGHd2epfM+GI7ytgXQvrAS+TPo
23tTqaSHhvuqwshKQOUUnX0eZC/PbqtMfRkea+IZVMMGkhsgebDCKzu6pFe/C3zP
OxvvOI45UHuVKytt6qFpXV07AG2qlXy0Ii9V8gSn/JT1043c70R1yicSlupN+2ZM
dhqTQDER6wxZ2cDEg7BLZA8ZHSSe6BgBYb3VKNPFD5xaIrcmUzIDesq4TfJ/f3TN
XMtcWsV3PRMm4UTARcRnXBevVt297kJHFoqF0Z9snhBwGH74+SWGilcd+pkex/Zm
6O7TFg4hSg9kc/hQ66aftXBPiBH1eDHKR4zp7ZYxBD3WGBEyRRMvvHV1UeATgbx4
dJWyI0igify02N79Hh62brQ976Xbk5AEKZ4PiOYm8oD98fNqlKqj6yEVitz3c8+d
1dhLAz3ZCWGVfydOqqNr7ren05ZKDbYNpoFTT02qPwPCMxOWSdR/ElVUKiWldcxj
BEdtY0dSiHUbKi8sPB7bNsICxOexGf8yjktS73MeBR48bM0Bb2SQnqSSGUyHol8i
eOl4FbfP1nqiNs2LP+ZuCiJvaYQYyxeKRH37okKfO1VmNEcsYEq7fzZcRmI87bPh
3wxI+6e2wl8eJ9yQl1MQYmAuS4jdV+5mcIHo0hlcUDIGGSWAxmhDZRENX7+2wXIK
2z9E5dsAxLtGTLROeo8HBkTIfXYVm2l7ggRFYv/5HRUM8/1MSqxpg4LX/b2bGolE
AReKajIuJo4I0Kp0tgxmQP8vpIHit35uFyew0NHcMtf38PK19e7kkTpLOGTzDBcn
mID7i/899iHFW6LCjS8cZor31R7rew866BzKsW5mi8BPh8WgP83T6/scmtKY/2nA
Z34qhxnFH3z6IxFswwF6RrMUB9HoMzecdqPiD9uPH5kK0Y4yUCre71BTjDHaBuma
THZtH863ohu38oDth048h6dvN29xhv8EPTYnFMiXVifF0gi6wFFxnKVPU6w3HfD6
Sbmi9IWx6OPg6aoobw44FbjRw0SkkvaAFmnf/EOTyFl150gxWdsNGT5jRoB2BwiU
/DemqsThj8HRsp6kgH+bhhxuT+Iyb+FheuNmHd9ICGKSOEkpK0kd6pApCKXY5n4k
G7yMYJKWXdEFw4ivmbRrMkfxPAPDEZeyKR2ebROQCu3gCy0iN5kZVlUJQ94EOAmY
4DWysvqXxTI/7z77/6SuZU1pPzxJwMGaD6qZ+Zac0FM60ZO8hMfOuFplHgr1S/wS
SokyJWC8LXmZkQRL++F+AIpjj/6/RYUGqB/5dTHhsmxQYjDRzajm51T0su7j9n9f
zJ39pNQ0vjw5lya9kJsQZaX2pz+RrZaEJkydx6Rm4IUuwXCpPAX9Lohb4DiY3iuT
2Qvrpf/ZNjTR8jUEcNlD8ggjF1EoM0PJS5JsoLSuRl4vrfkIuqDpp1qIZo8H/9ql
fgNBs2rGv9n/yDj01Tf2xBP+oLnhryT9uvCYHtH22B5qgEE7ogspVUR7AA9Khwi9
QXqOyFJHabcbkv2hO9yGKNjtudy5JK8hZDGK95sgQrrl2pzBaGhZYhziZ3sw9wdN
/zBk/DCvAoPzg+aAisNLiNoH9rC3B1WbV52Y7rPcvHWw8gNjDi4A4zuU70AP9jFD
EvsdzJ4+5uVoGvvy98RI9zjgyXGW2z43TzrLplUXOM6t1gj2cFRwsFp0CZGmC2GX
VZhIWUwv7AG8bZecibdPrXH52qRKYhi5o2rdM7GshnvRdA8Yi6kEzU9ZUVLodMMb
QEu2H0WUySCN6HzG1NihyUzGyqsemAsjtLlRIld1TYZqSHP1SDOqhZ3/TLmQBOFr
wPB/nQQQ0Nf7jeRGB6rIbRYj0BDQE8s+1U0+fDTtWtWr3ykCQcUcl8fF/ofoFUg1
gWNSFNFUF8wvFCwdxqP3AznCh0Jgx47Aq3/5gjpKway4C45kOtDXWZxdQGZ5SXQS
K7nZ0Q4ySpFuo7jIF0HO0YmTdBVVIn8lzqbKRs6ypjL4WHA2LFZqQOFzxaEFTBlw
YEBIxw82+YDrXYI0IWRxHh3kQJ5Ri5vouhUZHi8dAcssuQtur0lP0EvUNjLmNGuS
MsWzg2wD1wYj2hBef5DRkMLvgRdXsKCsXjPIK2OGHd3pAJvED1uYE6N9gVYzCSxH
xnHJHlcvWWhRL9Grmv5xJGYWatJ+tSSAohu8hSev4pP/HVmO4Id11Aq/rDz7pzbK
Tq9JcXTMW8SGD3iPU12H7SPvUfS/DU6TFzfEHrOEWUrDmhD/2I+Op1qyQfQTA7Hd
boAeCDengI2Qd2Bvi93UWM/nQ57FMIV1k4Bk92Nhvm8c52xiNVz8JsWapXLg+J7U
Hc/BC2OS/Ke6M08OD+ZO7myNTwoaWNp+SeYe4D1aPZNanpVivDKNPfYIGut2ZD+x
DwbintfWR5fSzY2Se9gJw7d9GGS1JtO1yFJ1k8PDm6GBJWPmT3au2wRiCluG6A4I
71knV3D1e1mCtIusJwQItyejMM9jY6pNhYMQUKSNeWZTRP2XyNnvPNHMNEosaGv7
wcDNjDjHLrRF/L+iigDAlRBbuMhaIWIY6Y37Df/qPuHkYpBorfLf4QJWd/rMEEUp
npW6FHDcrj3UKzpdh+SzFKP+dYXyXsTtY04F3uEyawCORYAoCOgjtLgjwtyVMWq8
k/pYFWvj/ggIUwovgIPgG0QU+CkvPTaZdqqfgE+IGSAsCeUmxqHEseXU3f1fM16r
lGTCUl5Ng0uec941815bic5tW6SbpxnbCte26MD+LGvzcY5WPgkm5x5fKosdMXjH
T6WZum5lcfzIkqrSIqdLKfAnypIlKb0ZHkjNT4ciaHjw/Wwg6VL7Bpe1x5nsgjpT
yVCHlTXbj/CWedn+htvdde5WrztVuN2IyTlRprmUeBaVfPEDoUXhDnAsR9zFlDPp
0aaA97jjwgibJPZyfldjjnJQm8KAnHMiE0FoTSmnZU82uhMo//qZKDa0679lvx2K
l73jGPM8sN8XAsgdIhJs5wNUAMMBOg/QP+UAOTXLDbJpiPz9BaOQLwu6feFoZ/UA
xoounOip2nYDpIlSV/xQb8YB0JUJWkork9dojhdGAnnwd5Q4RQYuZs/TweTzSlcL
/ctmOsOfHN/Lm0aLqwUcAoUWIf3OLpwfps9gGwd/sN9t1EUvA/qDJGp6io2P/5RO
/wCXu12KOlgI6L5t0rpJOWgIuUeOQyVTlZDOfAxN3+McIyacOHPPnx+se8Q0PkhF
TOxV+zJ+cvC3x//4Kjl5mm1okQ8WEIaf1exV3RUaxzzSIaHm5wv8NSj5eyzRa4NM
kkD8fimOpuuDNSHxxPdN2ty6k1AdaD8GIl0y4L0KMP9NqvkfShSGpg4d70eQThhx
Vo56Sk3PtV980evmpU0WMOFVC2RemI+GIhSI5lk+idIrszfRjWKHRi3zkzR1seOU
KWJT9MJ+jrjUcl4Um+Suu+w4rwGPWCjX7b8Z5Yne0T1nLSfYPWdSaI3ZZLnX969r
xGKkysFLz/ebI1kPDKFFjxrVSPCJiA5P+qZ5v4nlE6vTIC2LpCphdpizvEpqzZiC
S0Mn8A5cg7YOfMswHyXkdH3GLnODUww2aRxl4TcIyBdzahWM5xLSmhcxPwCA/V9a
MjrcUtjpUFXoEv6oj1X7zb1+7DWgyf0x4EMy7jB+rPl5t9NWm3hu/xNCNYPChPNR
fVKnaaARjhtRxJCMyQEjA7D3M7xOgBgufwGk89YTIteq8f2rbprJYSUOZfencWDv
7UFC7YvOGv4Li/BSkCDb+entlWsYjTC63UcuzS1Naw85rX/M7jhYodXx8jlKiQCa
koKKddHm/2PXYG6PYJmSNNtB3lWrvtdNYf7tZxhjl5G92gDPoCpnDYBEn9+TZxys
6AWmaR82aN6OT25OkbXLA/eM5fYSRlPFuZlGgjcd6/+dfxF1FGE65RQYQ4AiNeXf
JNhfdzfmevgm29bjYpqF83xkQabHBckm8eJUHypOgtGDM7Vq9YBdL6W5NrFxXOjN
iXkpS5FxZ931GFM4FIO7dsxCDPPSHF4rfAMnD97fJnjmJuuNY3qtlSqtjLYSrroX
KNykC/OKJO8sNJAKnxl7tGXjVQpA6rdykRPBcXOvkHxh3mfat6v+r3V2V/w+PaG4
eDyY/Cz5271weIh7K5ZOnUabliTjuyn+RkFhZVRpvqHB+YlYt/B7Rfue6+Aeh0+A
vMei+rlu485r66yl3v7eCzM4Vioub6T+zYgGyatZ5/3lMvFsXREdxJyX3vEAlwK2
nszmVqop/WUO3YzUrNei3/VW9mE0P0oOm0xyXXVRNFDSwODg6NrCWcneFdbkwQGw
olcjBjBEr4AOo09xJZL5l73hfAxoYP5/sCSzXnAz5ii67nu83RBgjfi1Mzm7pciZ
RdeFksOABYvB9uaITfM91PHOEByXRIPSUw3fuP3wCyHPE191B+BSUcJFvSHQgSou
8diCK1Xp5KsZSL4ZJZTvfOT07Bjl9ddnX/oBejBa8efNH8lH5dDw3pjmXBFchfXQ
KSsUE9vF9nJuBZ1RhiiuWW6oq8G3+yrNxDVtP1c29LjY2gMwWwnY8kT7jJBaAQt8
60i38KXjMzy4DoBLj82oOZU6P6DopLA1fV3RTUXBLrP5BP5OG/TReVuVz4W4dqVy
hHHsQCZEh6RUnwq51z5i3n0ew4EfE2BH0CNxfXOd7VnPP3goKRE9Jbqzo8XSlyph
le5ug/G3FG4xfy453k31e8vMRY+xWomyTaTcNQcR6d6R5rXLa9WpnOjdyKUdObGL
bfkN2WvsnlIqPcCUJz/KZT/HsvwZhVdDdV0dqHTbQM2IiN39owm4uTvo38WVXAjg
GPlOlqKHa26FMlKk/gaVNH07ebzoY6ADue5fG8Riu1rpkxs5qQpv3/dKKtZdGmXa
MaeN71GB/d8iHGGb1KJSRbYaNm/n/VYmdBefacVyL+oKvJ+2dT2P28tGzRbdGud/
TJTR1yezo5sEuAynhOYrHh+11213oyL2Vmqk0C+3j71CUjrUGJ4+BhuOCcLZy5En
OgpoidFXYxvKA9DYphSrEKGofMUljTrQcxl+5tNokXLGkuQEEge5QTUY5W1tVJrO
1RkUCLFPKmPAQbv/+c9lReeW6IKXnU+Cn5AGgxAnH/6lzqb9BdVrM8O23KybnQIg
/UoM/huqwn1UK6mLKoHizLiji4qyHeiQoZ+5q0gjTrFJtbcxH1jynl8lW2RC/DeY
oJn/BdDmn/LOdmVDuhb6AAenDU9RAS+m3JqPMxJ4SN6tp2LTxfDDLHxysYsyJl8N
4tsSMuTh1M+8ay9fMJRZ2gu4gGg3BmxD4OlY1PiTOP1VjNbtL1MVYar8+nIlSKyD
UrtAdTcu2IjlKxFi5ZZv29COOdmML/1OsIDkEvmhOyQy8BlQFIhK3obVd/egaedN
U/6ij/7YV4yda66phVgRKZ29hbcsZ98Em8AO+Mwkl3x1VOfLeGvEsbGdTPicI8B0
1CKO/5V8mXEklf7tRN41Z2Ah3XnSAK/Ce0Tw7X+sOJbk7zp+0h+ibnnn9jvbXHMr
ygHc+/HtXYC+wkJqvlUPm+kn/PnPClCyncMzytDZeUHe+XBHmF8emUaRQhXFlDRk
q+we0NKMH3gkcoTs99OsIhPpwe3g4LcnxH8HGvxtIA0bwbs4Y9vyNbjZLtIn+N0g
3WPs+PeVmEHvmxdG3VXvM3Mqzsg4M/TKefI+sRi5Ul2VjvY3iJ9xGralG5m+A9Fb
6XjxchmqNsotMG4mmqkpZy7z6AfJPYleOid9AZTAggFGVgPrYYy9ch+T8kv6kNel
AgTxpKwl7vMklP6Y3/O0Gyl88YVICd+2N6+uiQL96ZatpQ0WwZ8vr24V4fi4fNlQ
jSL41BtBU6bjcCOtf2AI1N952sEIMokbf99D5Iok+W8aWpe8PkjUKKlf9Gpqqt5g
vzL/VSTQM6X5k/sEX0xGTlBvVAzKyLniBawWEb1hssteAhatLDq3QTAObsJZouFO
/pIPj6cGANrLYk2GP3M7i9N9p/AVQmqW4p0yzTzkfLPXcn9e4Lrg5Bma6+hK3Yyq
fTAI1wYwTIeUUEtnp4EhL3G2Uu7rWpCz/q3EK1ReDeFGmQK2vSwzj3ZTzMYe4CJf
69c0qfG17YtCBdVtXrLDzvScD6tUn1EBeWTSfPoPYVg19Z2gdPt5ykwR1sFNfGum
Fz73A1ActtlaI/55VsKUG0hzrxQY5ySIZG/YOuqoq4WgiL8CKY/XHoR8N+xSdK1+
TsUC+W/R5bBkSrLyWLnLwY469fbDbeOXfygY2syVqOEgb7IO2m1PpUpk8yE9b9sO
Xncf+vjl6PP5k+yGCDjbZWeEz1eLYE2vh5spkfF6Sa7MV4DQFA0+s50F4Nhz03Tz
gG5j1AdMjBhve9H/BSp3/QaoJSQk0DvmJ5aUcul6tjr8iFjolgCkS9Oy4TTNkliE
lQd1rXtotzzP51ip8fpdHiAdikKD8ZsLW+VZNg9H1+GDAMYpG2qN9m+9znWl7t+S
2pzxOIPe1TgUYDdr/4D1jMhEblBClSPVgcqkb/3wRA2DgkLWKvzlUfH464pKcMxU
Y9SK8icLDS1H2uFFVHcgWTxv79XIfHl9yF5Cve6zKKR+Hlb1QgB6ZIyHup4zNVrs
mbkKlfL4JiiiVSog7yqOA1gxMgSgsEYETZvPNeBbj+29+iitKEEWFSHkARY1AnG6
AViU4vdbLwv8awKJYvknfOrxAY6sgOsndQDqAT8FyM5ubFMZN9PDEJh+hX2fQFQC
58bEpEJvYsxwCWTSQDNTUWtTOuFK+FugPvGPADeRHXeros1OEjwyNTNIh3JlU1Gy
mCx0irUn8T+zx4rm7I3ByAVDhTt8JcdjRsHI1tIeL0b6xo6w60UwMLIKS/ewKtUA
LNEImmRwnfpzC13d8y5+5/qzzk/eRNA2WcSldwlGHjt5YTifej2EzrGi/A7UlwAe
2KxLv9kJFEl1YGAbQDcDOW08AmIsd6qRIN10WRsxpyYUg/YCX+sLiIyqs6QfGt+T
vMofkfkxn9JpLwdjD5iThCfK9eUeybMRLPL/+PJKwSSgwz7L+PfpX855nUS0LtwZ
OSHt4UxyaFzVhw7E0RnU3zkf3O/1nWHu2ngnJ+UHvOFHljmbZriultFdUtWDPRWI
2YGjg2kaPs52MH86qNPuPXpumVLLpwuSyJtrXj7im7WZ0zxpoVoATiV6ehUE6xxn
lFhoAPsRofKGjonlfyR4htga8LEbsk0eBKvyUswMIWhLte6NQBhMqpTJth1JtAD2
I0Wx3UnwcBV0cSKyf0Cnz/SghmEExh3EEE0L4eTR2vslFF/575iQLzHnTr5ZzCjq
i224VVKrcfyB/WggA8rnIZkGR5FMbDJBZnNt94wtnuyvWpKo6bOhPEZFBJfNSdWt
zI2tL3bsb2V6+PFXmj+R17XgUHG6S0Ng3o9cMPMtYC5dKJ4Z1IAkmLY87v452Qig
IS4NtROnSYlzLPSH7jdoh+MHSLOXgrjHBDICiTSuqqkD1L0mamPiBEKKsDTmJD0f
wX0bRfmvApFpvLYiM7cLON1fYAeROr+Kxll1crrCks9cy9ETm4ZGP0MAErhldMQY
tLe4DJzaPfnLsUE6ZlF3SXfB9ZVViVkz5E13Lgx3SJOREkd6V5vFTHEZ8b5JF1Cb
btoU0yo8jjS5AD8Ovhd3AU01cGomML3SRZ8pXFENQhMAsV14u+moZ8T836/7My7j
ClBjbvFceYzTY16w0Ar6bMktnctOastflOQNKFBq7FaHhzq3D8x2Jj6cve7Fyxzw
u/Lv7Lh2JdBilsVllmVkKczhOzE9Rjpy1T7ggHQkB8IUwO9ZNTJS8giBh9xU0hO3
IOMvducW2GsQLTbvXzY0Q10gOGwpzcreVUf6qczVA++R4vTGk4S79Nd0T9eD+dUA
rkLtKSStgLn46wiTIwGOpg5OpE5IutVCPBAP5gmE76xYBzK9BfxSwUMZTHwS9i05
h3qVZCB2MDz3dr6g9VQfBqwoZp8uuTP9Q/MVEhCsYs9wN201lAm8odetbpee1AOA
c7LOBWnAiJO+frP46LJIZ6EaBuDGH9E3vJdi8ig+xSo9UhzhjvWIeeGV1N8DKBOA
kwnZX5PoeDHU2Mdrm9Mr0aIjzvKqhQrzrM8V+zdJ0L3V82d1kJrcw5l3NXN/WiV7
4eLcDwj/o2q8E8iQaQOQ8PKF5tivWLSB27xnPbU/eyJaFUFdjj55jTqtpkRCQ/PF
3r0Kq35HSozUWlnVV1RAv90T4Oc8UZKtGl8C+pvoG0wI6Tk5lBkRPgmZgC4wS91U
P41pnCupbILTRX5OIuebWWZM3s+HT6kZivDHchaAcviyoLMvHfnO6IGhCQUeuOVP
hUDXWRLQszxv7zmb3kUKKDJlQesIZnmKnD1q27yMFLmzsP+JAEPAEx4H64w9uUPK
16icw0Jgze5AKbLjQGcg1OiiVQsMys19Cn6o+jzQlGGdlOGN0yuNl/kT+4WvOOJd
l4MYX1Xh00uxQCMZ9ILPGlYMsN+WsofhVd1BjYcQnyaegPSrC2Nd4X69AK6rEtQa
mhvdzy93yyiEYMs3xWa8I+rNeF9NknvqdLShwM8ActlQ8eLXWgFy3kkaQx8mdMVH
C5sBGk1rwCowWL3YvznXYhw0TpA+QkHTom+pB8OHnKNSKvAmkJU7nM9ns9SgOcL8
OHNABVj4aLMw1/jCBI5zEy1P4X9gEJNdi+eD0h1VbU3U/kHPmTLi6J6WsanoYQtd
cIiyvt0hmJlxFuE8znufEAf/Q3gnsHJWbaa+Z6gHwn04Ckt80hgwkQAuyBlpp0i6
r92OMVhBCBrunUNNnV4Y1mE7xzP6u1v4LYAigZGInhARUnXdXfbW9LlgFFV19cin
tIej4/5QAD3C2Q1+LOPDID9M4/TU2cAsqS3W4hHA5aWOXBCXqjsyrSm3A3DtyhbM
mWyOxgQNMRUF8J4ZJt2pUKW9i7xdAnHX2vVxtdo+Jo20s84t7ss/Jh3KTWIvIpSF
nF8u0d7/opQblgDv9AdDH1wXY/VxXbNX1iJa703EVkKSy5bUGU0AdloO9zEALMBy
c4g6gFgFhCRe4j4bcKjR9fDNZOSfMo9cXG7fqWjqis7H10m0ZeWC386eGbLqHQNi
7X4iL0YlXh/CUhLPT9B0o/eEFBcER5zo4LoKA6Riik/If1P3nkER6yxj1ma91xsw
E9y+ZsumJdPocUBQY04gbJDK7V3KNDYtCvI5GWA4RLEnUYjucB5jCbR39qzpVa0J
xJbibIDm+3XOfbSD2DZpdzmixhNPkC4Ny4CwyXNiS5Wc9+UxL3Jbb0nzIavzSgfE
Io3CT47LxTALFlPIenyKM38RLKnqHJrLuHAiLUV9SsczMeVcSZPL70ZfY+2qYg1r
UfPg3qBu5PXHaeiT5avUrlEglsz5y3EO5rULfN69n4xYrdI2zEDsA4ltw7J42GZ8
iUchuzpJD4K0FJF6/Mm4ld6Yc0xu9G2SivBBJ2M7LSHCQqjF3zqlI0TjCE1ygbcR
MvTzHkplMHD3lXAuh5GxARNCmJKAkh0laJOCY8LwXZlssKCV4V6SjxWskeKM9LzY
MXEpvJRNhzNmkrqD5+BiA/29saOOonpr5IrlDKb8fqYsfd3aUI5jCGwJejrjUkjI
sEtQBKLdkl1KSuI1SLJ92Qj4lpW6+dOSPMQFWRPmbOHjfiPA7HiwUnGedulJFHL3
PhUDVSEHfPTpHL+VPLlgCDhmeGoGevHRveDEJ0u5JvBsNAACqlrNqcehNmGblW0p
3Bda+BsKe7cA9T479GrQ3028sfDTdyHl1C+OGWmLzZXDBS9+44B/SfDJtPJwMLwo
Q4bg9nkDnDpbKTOmDyZBU7deFrNrzik5SojeatkbtpEccoUakDjKplQ5DaJGIHpP
XOkmLhnapTOFuO5YiFstWlWu1P/BDt47RG0a2Os83+oH+zURiTOTWPKHuOWwaCUj
a0KFwMPJcbkzAKnV1XgVzbFkp2fakojE+2PIzK1VnNKsh4/Xpx+IJnagp5JREB8I
KUVYkxVUGolsgpwVRr8SwMVUIQi8t92xz6rhV32/ileT4+jkXpES1RphilUlItNG
wubMm2Gor3Gbs54mhCh7zKPppsf+j2kqFZiPZweOPThLfhpjxSeIGTz7Bdx/heSh
WRt1nkr30i5T2l6ooknL+xaM9x+ZWJzNB5Buuf2+yIRePT0c6aQueQwJRQhVk/+O
9wqKrCmUiLltZ5RxzcUXHFN9REyK3aAHl/Q9upCXz6ntnLedUeZLHURcvAZu9wqq
EBRKqWBoBBuynuznCRb9K/fSUxQjcnPyuxz9f7tKvKBfg4KWUYqfzQCQq4ZlQcwQ
T3RCpr+fZXuJBn69kWcBNc6hrnTtN2m1zhQJ+QxhoaIIXSH5bKFVT0kjMuezA0Ts
wfCvIonC6wJmgvYb5QK5ZcDjhKKDo4dGG5YGtxj6Wt7B8wN4/XZ0SJ85M9yzhBcK
hRkKV+xrHI3QW77pKBHpdHOHoS4yNMfaOBT0qlc9LebrQOXUk74v4IECFNunD+kb
9BRYXC1YGndJiHVR9fOZ//1/rA/23WcqtUTVeIDCogqbBNA1Y4p88CZBJX7oz7AT
P2MD24hnegY8QV0BElu1RfGDYLa+6KYMGXSGo5F4BZ+ai9rErgRWT43ERD8AbH5V
DzOGbFEmJxK3r83VyoXbFbm0NeJTARS/crv7u2KbS376lMaY2OoRA3czbeyDrvNY
pZnP55iIfJEJy9B1/lP9ZIAZePNNRGZP39OU5/Ha6LR3w/q2rD4KMYFwyr84lgCm
v1Ow/Z39R0GdDrip/29kqzgbp1rfYSU6HJlT+Z/52JbwYSLY90N7NLztX6jH/UXy
GUm5sWN1uwyyTB9a1JNJlyBiFMsAZkyzsAAsXiT6Giri6yYlKg4ZVdgnN7bhYlOL
dR7i+gqQsHThcBNyyyIf0r7M4Vm5ypAYCTPGneAbESi29DVRjjerkyVuwYTv1+eG
VM/+HqfdC9yzi1NJS8zYH23cktSws5JgzWn5eluzLsUuPbQXZVKFnh8s3B0XsHo7
wzzcO+hgh5B2zUwVaQQsZtICF9NM4aeoWYxBT8NkEnm0g8Avn+nb+gEElcuzENdQ
xNN7fX1IrA1g56Kg5dfqwjVWrvvY8ctnNKBoXDUswfKLcZH2WZoOHrGijQ6pRzir
WVrq+JbcS/cnmjSk7pSKms6B5P0on8HsvdFOD77BWX8Sjd4B15Z1BLQdA3NfzFqZ
nHfPvanYHTO6VaCFKMbhvoYjSjNK1m0ae7H8hYFjhaQOCl3Zb3O2IwaohJZvYjKU
wLTD/bUfAXxCuam24fqbD/+fT4mMvEh0wHPw4Qs1dVeQmNcelAPjuW/5err1OiSu
QWppzQhvnJWZkXn4TQuDEEjQZoXJeUTOdJCBNZtAwKbrNnasKu2PZCFHzV3l7e7B
MFDiqJOc8EsEyyTqeleqZ3Daj4p3AAvn0xsdvygTvEqiYeKfcl2UrhX/zFG6oSqe
lg4ICC2tUe76yMBXj6o2at4SLxvMsTB1yOuY/mRXy/cqob1xA01spAuAWe83dbgV
4M7+xq3UzlOGAuV60o3zdCJj2OYyWjd6xNhJmMwHKr64fR6qdHcyxr2VvSqrrovA
SP9aS/0sSxY9ppoAorQBB7Jo0+aXYhKcP/TIh2DFaSZc9qRmDHIL4baG9Yj8xKFF
NRWjSQd787ZatftkHWc07nhFeFp638PzOMnn5vTMXkf8la3Rkh6fpoQwqBuN5dxV
7TNmXVTd0vzEdxC4xE5oA4fxIRPJfVE9XoCys+I2K5swLtuJbmu1jQ9V4Di+TlUz
PP1XmwMKwP51H39A6pHeWw+ILRtlE3yG7R74mFnQ/XbzYFTJu4PT+0mM3VHQPkgC
qOcN6gMf1XpVDee1Pl7WQ5ABY49woszXlI+XEelgTH3Q+v+zLgt+DfGibm+eLSWM
bM13RrOMvGanUMC9F+b/4zddwz6hLo0Mm8ChKd6l6PdsR5oFBtKUKvXDIHF6xHr4
HQEsumBnkfU4DBIap7CQ7txFsWRUbFEdIC97UXwnNCfK9fwICBzEOKCzbbQUNNdR
X8nLtJyVabMXMHdIPNjwX9gZmhUTRseqcNKO9A2kdWPQ7Ovv2MMGVuHzfj1ekvrL
YGYkrkydb2mbZQJLbsZ5u5x9fA6gt74QySvMjf6epAKMrEZctYXIqz5ePZk2yEqy
b48JPjsVe15KMjx4N5GIyX+FCF3EPKYSE57CqyI7tbjzQxtHmGEXcTR4ni+jBrvv
HXcLdjxz2TXNoFv2cNWTx31h2eaSA4CbbWgpwAe55pmz8xdmY2Dxh+u1kqoB6muz
37w3hNqdqHMA9nx2X6qIMAyUPmUmz+AVFHddZ6nIHv8gqmpPqcolpnO16qCr5KiO
+09Jw00r80LTfpSXlV0EtRHF6UoHGrqCu6LII21QraVVDkrF2Wdvk3N1y1QDdYoz
4Sq3Z2lBCZibHWKpC+Uav+aC+KLAGy1o3Ftmltv5mdzTN2wQmKpdPb8H0BH6jEVi
JJP5lNst01+N7wTdvDMC03/dlaqpKvuXen6jg+W2AVka5XYLHIIWHRxqGU53zWHT
ZRar8ueagEINpMZcBu3ZgGPCbb4ARbcCCyP4s897ndyuaFpsNa5IGRrF/sfzEjPs
TkVmugcEC/Yz2ycnjhPwhKHHOxHf7vDJ0EEjyHUKmLsJ75YdZEvRuCi0bstzJaHi
pv1Vd9KyAh1AqPG3oYbJBKn+me88Ovtu2s+rOuh8fvyZ2mFHdv3xjlBjj0hjNgM1
QnI8xdXufUz7ejSJQwAfCj2jJszNAHkZLQrZOusYFoUFKAMcbpysDXYBrNM2TGIl
UDW5cEn5Sg7slPbNwCjhKfIxkWyAtft0Hvso6JzW9l+rA/YN7H2JQmrRVLpzZq+e
Skf1d2Rp4Udy90oxH7XyV4vYSEKbs4AI5YFVaSCmy/q1cUbmJ1H4SV2HZ8Tqq8DZ
JzbEdKb2kRgLRn3GiKYiUIee65XkWmVMsvdm5HMFVBaPL/U3m5VcXgcYQrVPDl0W
l4mpqCuLGabipfXevgJXBXocmdt+cG5+7TjPRY9plyeITGdgE0yJkx/zmW3h9xaX
zuLQ3KH/2dV2kH4aLTyQJwPY8QrGYCCh+6g2mgMSOQ9VKs9DLAcQvHNYUKjazsLm
Wo4J7xc75ITX+PIrsx+ycJ6ujAGl3fFa0ZxV77JsbeM0ddF1ISCI+wi3s7CY861f
HSeBUzpoRniqp/ThrYB+cAl/FabtvCNxpgMBrIpJZfW/KGY2VRBdk9AII6d1t3Az
9ZJp/BN/+bV6DXt8tjH017WdpEsiIf/QbKUAGSmc2d0StTKGHkB6BPd3h68ttUX4
KgfUFezVhIqWEtEg1hv6d5Hfe+MWF9J0rM0aHI09b5Pux1VCv9vby11PMFcEESeh
fpZwoPoqQDtNQg2DgJetzlPXy+bqCgBLBPQuFhxN8WfpPZnfBDw/KyxEzkd8MBzn
gGPa0qfc002j0E5EnE7vAedTC4G4r0TzGm+9JqnTpX0PMc5kLkJ3IGTo5tKM5lou
ySO1Gj/URaIJmOn5r0ve+LCpmlf1rRCK9MOoh/1q6zkt8vwgF+NYNT3Hvahvngoh
FVeGx9AWFbP/4BC3JxgrRDQAIRyko1tDiGGkyF6IVQmUY+BlcXrrEUnUiZ5rTSjc
e/lzwe6wY+pgndag9gNliQ0pGiQA67dAk+E717hcDSSQM8Ox9Q4UqS16tWYgPMAa
txDjtIi/Y17ay7unuO+AfNIrbEltLtylMT2Q49fNMsuvD9SnK3k2Q8bDkIBf3TBb
StfO31nWHjfarB/tT4N2Ml6HOgCMzFf1r+mrduBQtgV1r/3T15IatFGQ7WHngVRa
tUpoJuuVdVvyD+zAsCCGAqtJMHHkpy/D07ZKffukAOMn2r4X/7TvJjLrVREy7Z45
gqAN31AW03hVbzphCXKAPpgNSzJbgtF27e+fgrufIRyIP/DixCsI/97zee+K+QKm
ceLL6oI5phI4WD84TR7wNJoe95Ou76ZS6c2JvXq3CpUVdjsf81I8suSQVBN4WamB
8FPLujjokka+2RvZRMIjQ8OU49I7HpXrPHU08P3WxEIigkBbpZoQq8Cs6jbSLbGP
s+18wj+1YIGJBbVE+5T83PBMiAxrdr0i/MRzUL+eFH3Rt9YzrC9ypCnC96gfIEs8
FXnlZRTHpgftzNItaF5ijCbvpMqUtxXoe9kpIVf908hGS/cYKU/vu5pCYTIlYvQ5
D48OTEMrfqYW1s5J3aOFOZpqU5/ohLB32g+X/esXNWjVacHQs+lrDBSeplfOBUNK
mDLUiZjT6N29knn7BHjkNRRSdoYF4p6OONIk1J2rbmEWyK/2ybRDV4REQ+hOtXFV
sIHXzMvKOiz5mTrPvHqPj8X5Ljy9M6gU2sZARN9gww6zeMLnATQVJyp2LFJdjwFZ
GR/EkwE9DIAs96yfUBGwg5VbvO4cIdWuc+rAeW2ogHaVFPNELDjiIlbUUTQohuhg
GOhCLviiTrtkXVfzNP3TSIVbdF6hYyGqeqcTSnGhwLLlnm+MGqdnD/j6Ok3lFQAB
fVe6HruzHWur35eN5fm5Fr1uBVixG92r08R3486FFF9yZm0p2Se4G0I7QaMLlPRf
l61ioEAQOZHjtAsj8b3IAdZ9LO/Ttq+5NEBw9J5aFYFeDR3+BJwVLL68g8Fb3l7m
C5gPw0RIje5Vbj2exfru91UPmAaNCsYgY2IPc2cAfQJSDpXm5LE/Nxp/RPTkKQhz
JG1Bb9xZygMBRE8Razf37dPcAWdK7e7HG2AMJpcHgeWSCWQoNTTYPOGkH4xPnD2u
ev8j8rMuNas3iFvJv5Z5ZEWwsUnNDsD7IWxXNZVXVGQVAMhww9oy7/c440uX82/4
iKJcJFrv4Hr6h5eK096U7zpqaLyBFYWpy2/jYoAGHT40Agiea5gpTgrzILQoC80j
ZluYk/UFLJ8GPstT+B+/yrqNo87UJ7z8F0YAeGiMuJEmAfKz3Ba0JUw69ehpQ2PK
Lii0MDEfWYjOXnuMmw4zoCLwdXa8IWnOK+D4FhTRl/oVoM/E4/WZHkw+BRbUZYar
8YNzo5Kj6SvoKUxa1qa2/ym4AHpPvxOnU3ne2CHaCN8jIiN827WUVGPrsg1ZKZSe
y2iBkPy+9uv4cnLP2Wfbdg5c+tSMKkWW0SdZrR+LefZ60jJq0JhXp/IPvAn2CIil
89RuM7tidtnAQORyK3WxW2fcHCg3gJAYadtrVll9lkFCTF05HOIK8EKOBlfplzPc
RwWv2UvUsvdkMTZ7slpu8Thdb3LuXSuA/3fmvmWeu4wW0oGagqHukY5vAhdk40Cs
MCyTyrJv9ASFcJShzMmyAxRIV/PQcAV8Dj82yq6gR96sIzw8mZl4SbhHdhcxLAYm
j6bTd7lMdKnAY69eGdJjenO+Po4SdRbYhJaZImNVTa3krkSZEGz0Olu+lB/K4n7F
OXGPJvUt8xKeP2ZUeTgzDgIGunP1+yvMUfK18duynmRqab+ojnlFIfot+5cZ59Dv
pwRtLd2zVH0sRf206GJiqK5ZExNGyXyWDH/8W/lLfCQUw9m1iLsopmM7UoTcslMk
SJ7mpHikyi0SmCGpH1Z1GbzkxuJjv7rYvAPiI6vTsI5rdOKWn8y0qv+HvNh6kaff
m/OnY5qowG7nstG4ioPphhZjhj2i1A/RpBORli/SJ+m7pUGSJxnf/lh7g/02/e4z
La9OUfR4/PzEohQg0OdaAJ6+qmbRJvrB9U4zgP+FrYTyQMVmajurkR1oV4sRYxfd
nbx78sL+/oQTJ3GEK7VoURRSY2aaCyV4y/0VfxIemO16ry+EdSj9KELZ0YI1aJS1
dasMFkVcfzD+vU+SQPPMpGuqYJVU7KpbfZUQtHk85g3KOlh0BlnD6vmSNboDFvot
mteajpSjYys/2jcJliVh/+HdhfAsUn7p3K8mrV17AmqhuysRXhXII7pBllFPy2YE
9oRFFoF00THVRhIUyPOhP78+0k6OjFZzhQ87+atprQw3a6pXHCUOqbYARTP81XDl
mQm/cQkyBgvHlsgZkDTVi1GxwbeetRQSxVtc/xPo8/droJ2/n3vKrANmhz6vOnKo
XTKAsgcPVYmnLqBXpKTNlqFq514ggah5h2K5JQZI1T+/lXQJOR73f1bJVDZvw/2K
/eDPEIdlBmtN29nmj+ftR1v5yozRusxyFtBjaiYO8HEomTTfGWg7fkWE92Y90Puu
edDRMjJVfQqrArB5qr70THhSWkWFpY9pRLcUYKnDw4vxrBhXZye650ngbEAveGSQ
On1GjCtB0GbCoKjlFTcbpUYOojGwrZYxLBcbPU/2HoHlLSELxftXCbTaTsdR1C3/
Ve2B4L4brv2ON+ZkFMBNdgmZf+WfPhznEf/MgddBOVksB1MSQNgYm1NYISGojEbz
X1TXH6xEnw8V+NTwQZ1j8Da9hTwneBUgmV4QyYzttmLKTYwDJTep8ZMt/omS8q0/
NLGlxoEDzAHHnYu54WgQLZts31CRE3M8FV2Qz+qTrc5VFoGoBKqsola4kKrQY55/
uV89eKpF2ipNroGPZ0Y4Uzsn70eAVoJG+PH5sApHEdqSRPMFFER+rKQg1xJ+Ide6
JCCxF5frVfGp0s6xik5GwIa37CFoj+l2yPSxp4S+SXlWMn03zLo0UBSP2GG/GOKS
mFrvIqHLeWWgVSM0YCGscBS4s+j2mjXaurYmkggcckDuIkpy+s+UHqOWo8LuiaiZ
bA7eBroXUUuf97M9X9gTn7kORp4cMLLOZ0ztyDsi2wwj4bibltq2Brr+X3wUWZBY
T7UyiW1etEyi4ZMLW6EBqtcgiL4TxKMOzQVGC/WbXZnjbHXBZ+VlI7fklsp+FRM+
DZhDg3kqy+5tcBgpxHmyVwGAXHB5kSfAVEOgRSdQbEpWGGLjFIJiVccHFOmypxSL
SH/JtUf8Seng9ByftMfOsgiHGcp9Gk49WltUO0ocEtVWoj5eFIjZyJk5WQTfCx0e
AZV6ZJ1IF1elTJj45tjob1ByamgctPBpvekTMulncw7Ui7jcYYeTE7p186ywokJ/
7f19v7gwPkCttdYpbZJti0GWpjJcoaii1Rt2OSfzsd0/FZatCHbitZjEofqEkjag
vhRPL4a22I8oBYonBydjhiZrdwWgFNbjCy7d026hd9envOXiLtoQfUbLKE1+bMAC
/RvyiX6w2EMmsDoDyodMfX8LTEvDxfvlUOLXaoGauNJfUbyxnxdiI2YJi0of2DvW
ylfSlw3c+E8sdfPBjc9H/DUQHlrz065P18h0evY0eykQ0nxSprDlbRKyo3XHHrIr
f5UXK03nBclP7B7zInPBE4Bn+Ek50g89bYo+BWeZLPvvf19JepSkhmJz04N4N+d5
n0HctgYBtlE7lv1tROPV9AOEQXcI0BwGAXM/+0SpuaxkEdHpIPKJnpUWwJJfxnpv
FDCjA1fZWGVPFJcv0m0KC/fjUuRnbRx/mLBpguqs5dYnnUrS2Nt5f5Fj+lfz+cng
xmzdmGVOiXuIJp75crUTlfJQFP3rQkw5Sw95Ohzn9eCc8TyFHUarH9lBTfMumkQZ
xIiZsag2JFxCPyuXVjnohcfWA3JVHDKV2q55mrn3yH2rq2XvTMlhYNJBIYJLIYU3
vcMT6qTluriA+CwS53Q6LsBuLTNLUOTeMPLBBDIthSNckj+XHB9652W6Q9wFDeka
icRfhhAUAti2Ow5QtSRMK6hPh8KbV0kNpZHqHmbNStvArrrwKVqQKRyVuPl9pbun
YsYnXm13j06IH7taglZl70iex1PVbT/Iz0NOPn9Z4FzOHd+Fbf955Y6XXsisLEAn
f0Bq38e4vl+FcegwaZU9iH36d/N4oquJiiRIYewbL5B9ieQgWEHrj2gaHdI0JZt6
aLO0DFavGWAxFaHCrvJpozOA8+G1aZLloopND24DiUNWd/d8TdMNYBqbYqXTnXrW
XB88nZBGNGLnPlC28WBI7vostaUusMzzsWO/NsMSuk+3eZ1NoznN1X4rdOca5Q3G
z+5PR5MYammY+jz3oaqjZtAcAtbvt1LEf95cV161hiRrRw1ZVlfWdEAhOR6FpCHI
IXo+RFVyUfE5RWlk2ZeCvdkhCPBol8FrJzROpbW/z0g/2O4H3VpRWPHCv5trrLRv
/tabKP29uHSQwt7/sHaL9usRNgjgtKeU72oVJjxI+5Ee4vAs9zsSOjE41VAOcEqs
AZcvh1knC83NzlCRibwH3DvmTmTAtwSyOP6w8T26tp5/C+ieAWJShgDZoCazhLzu
+NbM0tl5UMlDZbXRpfBM5lVE5/TCh35ykTsN0jIYgRzppZxUHFEccJzUWK1oYRlY
7XXVR8R6EXy7pMi/7WI2QSoI73GiY3H17qT6EYf7qdEQDV+RmJmebjXpo6GvZlUA
QMtZ5WDMZkZC3hVEYWEZK8G+h9HIMzL0o1v4yhpRs+ZQbSWWBiyCgGQROc322Kcl
PbVNfIrtmvNQR3MdPvUrRtXYDAJ3M1PUx0IKLw0xwjncNSgC+yVtO3RmgWNEJSfL
IZq6TE9lw6WZCbjpKdr6jB6OmSHz8InKHCb5BNpetJRM7bCMlvzQH5doznHA3v6g
KUYroJou2ZRWGB4TDIbHztCt9hqsuhvG1+0ZEWlapx/ECsDWVkatXbzoZNSu8jD5
EvfvRhjuXHHKhLSG+VFryMTgKpwamBtPOHH6k8r+iWKv+vVT1l6RqX0ruMzE8W9t
495neaLVDNypIYLZqKy9Jf7owVJGgzD10oauKac4PoLCV8BmL2hjR+CQd2EM46Qi
mHBc06K7vSd4xhG62x5gycORQg3Th4bDXbP7fTm4/ZTBXwtPmbIYoGDJH0UsHz4V
uX0lQdYsWZTwcVN+fYssJUwdHUj5fcE4clUu1WTTP3l7x4/bK/0P4XlRqMav2bj0
rq7OcP6j8fAelsMvfFKjnTKW4KCuTej7zLPfKu6G1mYqAzk5pQn4mlkLJSV7Ktwh
t7+E+FsE5DMu6iVsNO9PjtsP74sXqBW7sniNN6lPle3bCCz8+CQh0jawZlT+p+46
Ly9dLc03w552cB1d+8c1fhe3wxNfICvyRE4mHJdKHaiop8d1mIOrb5rDs3b3EFGX
eOC5uHSmlLC45nLZQpxQ4oWQcNBckCVEWpMv2nO1CfpGo2kvQazkzPm/1kf7ATO/
CO/pCvM2X1MuyRYPPmLFwKqLD5xbFlIDNnVaIb5sJZfGw0LDwU2vs3RThuedG6Wf
21f9w+gA/cB80LhrpIQohOGGHpfi+amu9mXIHECqX6PwJ/u/grDIGXl5U064/tdA
VCx/7cb3SxLooC+3RdWQPIFtaP4PM0GFAgVOXxo2vKjHg9VQ7bV5kToyS0gu9lru
iRJIJIy7CGkuGqP5VNxbzAZ9tn8RKrqfgpFgOOf6hUqoCkheD1q07Pclh3wLBvwa
wywGLcmoN5HWn/4wKOxo74dWGdfjU/nCqDALz+ZC692mvX3LMPELq1VLyWq4NPZb
8XLDS1jCJsoCqSfkpFiABU8WDuzuNVnoqxCnm0MiLbC3P47bHSHsSrrs5RJek0RF
lmp6Nb1RmOVi8DL/F3fgBoY+HqgDaHB+oDaLXe/8l8kCjCDgN28271vwnj6VJLee
Q2wA6H8d/oNXfUW0JzBmZ0lpLj7Q37BbgQZIPzhblEU4oQkdCCkJ9ac6ECsnVnx1
v0yl2GuKk0jEkaeT7ygAysyH8ufGsSMo+bAfvcSrEh6D7ETkQmXBb/IjFbWbcETz
746MhwOPC0Fif3IurJkjVpfIiMCMAhYrv9c8/xEw0LxH3LkLmJY19ommqu4O//SI
eU/7mwF7a1yqEAW6v3OTCr40xOIhRIzsA2/cngeN+uYzDx943VVjV/7X0xUbr5Ta
1iu0Reu/WYyjrs21K9zW2CnhpyFzOGj3+Iibg7RRes1fpj8d94L5JFrrHrSn/Q4K
/b/mLab4y5RovDCT7DP3qvh+uBrj9g9MVcSeDpzD8UZJRaQNURloeSy6JtU/hiWW
k+HrxT4WaKKMIj3IMbL5Hpz9BDJh2gsexxBVKa6nD9PHfSp4VcylcC0j0e54ANHF
38QUg3WnuvrxZUP1AddCJjthI5cOSl+HdIbA4Qka7sqvlDRKKZhU04RgprGsidzT
v2RVBgXdEU81PEHVur5Q0MD+5e2ryDSVV4ooK/xcAfUzggunTgvY4v/rPEB3AY6K
CZPP9/vkxJFiL04E0B+5gtZoVTFTMcS9nZ4BHj9oRkpx7YM+1rvZ+1JST8dYT9Ve
xWX+NToRzoux20n6ch6dxizxSwX4KiwLofHMv+1y9A508l+2e7vwe/Zkpal023cl
r1E1YGC41bfGYDjbx25HP+hmGW9td7zpAM2upyY6zAbuJ0s9GVZBWJvsyxBW2uwQ
FuYP3mQlPIqbb4GSi4reKc8UG2qTGIwKqHOgP2B9UTorVpjgIuMN+95y5MXKkxyk
1hu60+iqTgkWKXe9N3/P0yBqwfxeJT186eNuG8HqOjobB8zJPQqTapNqr87H+MLJ
5xHz0zTCJW6gwR3+jUxj+u5HUEzvnNHpYumK8WvvJprvews+jjLQo0+bHy+irkag
sc1YkKsREHoUyUDdgsg0RQLIDLYTmMpUp1Ok4nn+5WXQjzJg0nebt8ioaGuieYdQ
rzflj27h/RZcWNO5XhJyCLCTI7GZ4vIIbuxsG5fSsAJrC8AlLq1vz1wKop6Ct4rb
4zwyx123jglgrkqekF6gW9noM58bwDWAKG7pmkKjCKyyTTjnRexeG/RzsIpkmugY
vzb6Uu7JThyJKBXYl+UK/4oGW5Hzo4AGEFQS1bA2tvEtP3NRwK0Gz9yWl8a058Oq
NBY3i13ERZi8k38TH2jmw462dDCo0fXcGeYZPjqDYGSdpy+yoM24VVozCWJvGVaJ
eVtRWIwgvZ6EnhOTUHCCmMF39mNBLAcKz7hjw2khZTGwweWwpzTfJiRkg0j0vkxr
u1ZE4ygvEBiyGjKm3e5XJDZC13mSIjUfhfyvgFjo/cQRXC4wSiBARq+uiWlMKneL
E0RlrJk5xD8V12z3DX2gKo+zUzV70K8hZF4n3Lvo6D5qwAt/aKIX046mffKy19tY
IWONpf/RrmTfyz3nH/wkAEkFRG5/4Gn+PkwES1m4HsYJ72WEIcmlF4TuGc3snj9M
EiQYeO4ZIqXT1ZoJUxWPxy086cmfSKED/y0f9KOdQ5E57XI6Brs9LUQfod3saywC
i3Jzo5ZaQ6X38NzjVWh4W3AKa0DOyVNxN+dMdWI1YGiUwZgl3ykMHCyNCGG89iPB
YLK0bX5XFw0DsXNZmRALCpW9O4Ck/K8sdQDQ6+QbQBQs+DOMHmVuaOTEkzBvOEN5
wgBUVDADIKQ53/tuQNwzm96w5U8iA6JOfb8PjjZwoVxvMXEwPFV/sOOotgsxBP9u
WgEQmnRjG7DkRd0LvGsZz6etbiK9fxDYza0F84NLahAhmoQqGJYMMHvZ4VbWmHiG
IfPvldm0BiRIAxqjaZ0Tu1TLJA0XUqNgZLE2zAdwOkTmrfDcFaXOOYLsoOmaR+i7
+B5o7PbnqkKnbKdMCom/RgC1PG5756DWH+Ac5UOSJAvFFdhVRtO6UOUbEjmvf120
MXAN5dNetEcUUjPa+LGoCywFq6AKLAyHGC3rJDiGHcG80q0l7z6U0MsLHQqGFgYj
rRTXWsNAvA4zC+/AZGQFtuF2fWx3FsiJVU//+GHS0tzluXylTxJ4x3px8ErstCnt
oD3kZlYVKe1gH5ZiYQV43QZbRCaNZxGMikjXXq7X4EWXPxaea54RRbMC9yjDZ/1Z
v0/39swLlhwgenTiJS4LDWliYNleWR6VqN4ZvChVQ6e0a+bznZTR45zQ9eP2tC2m
U0RjIU5KV9LwXRkBoO0FZUC8dA2IOkQ0nO6O0nHlHj9BmO1pBEAFubCTeBlYvrVA
q2AIHE5yKA+CEReJHgjX60xZwH6aOms62lNia/824PomSGAxM0ycpKlUJ9J69Wuj
2EH1Nad53DWPtguB/fFfjgv+pH3kto9KsTFMtjiT5KgaCKIYfVMHam9IuhVzVk1U
MbDS93CATucrezDH57hc+Nj53Ufnqi64KvtxKldw1r7s9FLDhVkAQrnZTNI5KLpy
noepVNkZP6oqUOkAWyCMY2bdXbRoGdhRRoCjLDSme6yEqFr+T1GEw9ui5RdSp2Qh
kgK+nBRcfDRd714flt8kNTNQIH1YQ0StWI1y4zbXa7sjie9CwZlcd3RR4IMmIezJ
UddZSgnm1EOrCdZi4glHOj1W/TmuR7u1tPkZUGyoO0WTz0QIV1rgX6we2c5s6MZa
8fJcQSP0NHcus+Nha4uBHTrmd+VLQcoSUs9vubmisMhseQhEK8nt6g7drimzUt0L
F/rEYQCmwIKFV0j84xfutJfyzllS9WaHoRjAdafNqVod8FVZ3Xc+ztWjiaFME4eF
mWXtSNLC4wsf2qH4tdcMPqGi6YKveOBWqSLq5Wodv8TXINxQam3Bk4O0hGpLhlGs
LbNKsFdvqbZzvJ6wwT0EpQMRMsGCsYdkTm17z1iX3poUaVqFntDL0KWvcynOND5r
fsr2PehOC8FN9cYEj0zG6yNXfzVBNOnUgRocc0YfJn+F1+sKpOXHM3SCel0UrVaD
V+WCLoKxdWUU1WdDtRFS1k88u2S1t78WGNJksUsByrLRn4xyxAlonvyhe4kxcHDR
L7Bu6w2Fj6YWJ7SutjrDdXhSgUmS/cxhHWwqII2SbWxnwgJv/tj+gV5g0az/FRCQ
ktLuXD/2PysylPHSim5MDoKL4mWfgA5EY4XaMbjb07yUW+U2RG0iU0lmzlNmzX8u
dqMNqFrQC+PAJs4t5RLXYNOviQJHLVaRODSQLj6ltIUsJ5tAj8Y/8yi7pNugHXeV
gg+zA555JYsD1MlnylWTBQaz718ldCdAcAiwOTyfh5Fb8Nw/A6MWM5U80YGCKfVn
WvdHVQSfApkLV9JzPBbvRXlPBQ/VssF57kJ/GypyIR5bbHyZsRttOIjE3tU6fbve
BA2FDq3bkXAx9S5d6NMark9INqAMfuI7IeLDF5/E1HEbN8Q4AZ7EFSrHDvOeXYV6
dhMFfHso8OvWc5fxTFNwAZNyizkS0xr8RFRmWoajOM+gujFVWstW0/73er1F9IQ2
lqkNB/c77poMIenJ+ufiKrkuikdD+GM4RZJsRfZTrEAetil3nbB3+WW//57YEu86
8QYyDT+WqP816Jw8thV+dDpQQEhDG/cJPs92Swd3LcjorN9kDbqrOmwSsvMaZe9H
0SYtAxxT8kk+lN0H7q9bpOi8hY8WxPTIBGa2A8Nn85fRM6bggP755XMT+pJEVhBH
eapRP5G3jRPQZgwPCkLiQtpFPs6oUwbB+IcagFB9WgeOQhq9R7CeeszhdE1vLprw
AfQD+tydMr57lAIK/OLbNL0sS3x1Lr1Fm4ef1iCpS34qoxBeXRA3vLn0auL5cNe0
yAm4GRJ6BcwiD8nABJsGhQS2roWxbFy2saCAWB3cu7iciIFLxx47vDWW4S9kqa+x
pnfUwGCO/mz/YOpnq5xklHkHs3jycCe/x7E+WPFzuGMz2gzlg9ZBQB6MHfjtlA/9
SzHAMJWiGfsDtt6kWAiOSB5Rwqa/yjds1oq0IcAVRZ3v4IPOejk2Vj3qLBn8aXQc
kUgbblSGgw6tRc/q4njqDpOAYXJI1UNNt7uXtxHYy1JNYI7PBK9aNXUBdCa8Fzh6
hus7uN308PLM7Ap+B3iIDG9iy7iw13jIBQBd5rKJi75rlBD4j1rBZx74tHozulN1
+tDJX6LRKDuLcsgMLDHie8o9O5ix3SzAaFs4+MBLD508RQEgg+b2UAozIRjFkTaQ
NpZ+8tZ6tNaYvZ/nr/A2g6gaomq3sEqTEdTJ2VFRQZbckv2+SaNEgfgzPTQ97fFr
jJ7nDz+LdbK2GlLLTQAcZpd1RJBneisi4GdH0LYld4vz/W3pTUiwnz133DOHZcJ1
Q3VKBPhGLP6jUyL3vuL8L/dJlEi9F/T01gYLhXD6RCFjG9jGvGmtBMeUcV3FTi9S
xqCBKqtgev617qGBCV4R8am2bI6eWQToxucK+3sDpfVld3nh/PbKbO3bLhOf6fH7
lgsLKKgOHTL433fjNzdebbCWxdXR4JDtEa3ikoJD6SuX63Rv3IWTkMlfZMAbSRMi
QnliOBvOzuaWOBx5+tbl8G/aFF5W08lvcey4AqS/q/lKNnDf2UFPol16UfV1bbRt
2Qd60ratH8/n0Y8ygzS35WjXViNMS6iCyOvpeS8vUKo9dWVHTeR/CkTCSvWcKSyV
XW6O7+ndEp5wNsw67sroeABgapuUkj7Qvg5AIl8hvN2aw2ydT09IiMXURlpOwWPE
EoUUlrc9f++iQV72tDZi/HNbnCRjb0sc+d0bO2HKb3vCowq7X8YylhZEe6tBINVe
z4hT1RkUc77GA0s/ogqMEvMWNCacESb+kE3HXfgI9nIVrS+w5p69fSuiFcTo6/y4
c0o4pQgYoYgxAP9oDbfr34fWm2h9x9Uljzuy/9nWSJ1/XWBhm8U6zL0d0z4Ku3oB
i5fxxVoVcc6APZYZ9Q97dV0KWh+0Nah9kFNeGhKqUu/91RpvXZxBoH6AqQEANsUM
6vGFs1adnXvM/4X4xK2m2+Ge0ypGi1WXOMIknlli3yKxNURdbHZlDlodPyrmAJnl
hE8vXXKK3IY/p4BrAS/+m00CQcj15BdC1yjx8V1aHepga2GHSdbTO3xkWzYF8Rd0
4jcqlY+hatvnNEbNufVcTu8oCz37Gma+sKR8SJSzrOGJc9ktrspOR4h8u/1XsxoQ
Bn6kNyKW/iVlBzKwMg/E1a0PWDbjipTpGBgj9R5zqSEh7iJJXILAP7ohp+EY69uv
mAZTacA4xjlQNV4TkQ98+Q==
`pragma protect end_protected
