// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rt7kZxP23zx1hHGgLd4WU+bP/NL0z7XAGDZ/fmiDACG/lJaCL38K4dcQGBFQ3CEJ
V7TpX7PU6yjFq5D5+KN2kspQZ2nZBZNAyodm/Uqx8+QKFeRajeWjmH/1AwnkhVZZ
3/Zg8+1pit6/cA+rB3fMUyvn9Hw01at5Z5RBs5dBCmk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29728)
m3qBrd2Ww4U8TzbC26GJSruID9bOrjwjws3iEsejgudWmlwqvijN+Yj77IkKfC2e
/y2c7jhGRzR3U4wvlrzoRLBK9CIFpHeVX20K3SgvQfic3z/Jf/VnYlX+i6xb9Oi/
2k08P90z5SKcscXQo9Frl4C0cBLE1QQpdQgwX+5lnjjta+CIdeVIx5ejGT8EhDUe
AWoGLs4zf1aN0bWAfqsszTW11M/cioj/ZEfzGaLviaStN1rkZwuTz2MkChkzV3Jg
rSOASg/qP/RHQZp/ULCXdn2EtyuUTNj6zcc8rqOv85TYJ64WBTQl7TGm5Iy7wM4K
8EVrhC1C3+HS2eyDjf0YQ4tQEJbyTlcx0Tms1Jv6O5Q79nLxb47f1ssSaJvX/iYs
FGRj+Y0HiNJ0KNZafnrEK2kMm98+wVLvULK2ZmYX8FFSfzZPPT9XuK57sPDghxHH
WL8JbMZd9Z8RECFbA+5hi03coh5gtieXAoOng/9a9NfWmruhINJcqdin2mya4mg7
D3GnNfWz0ZnGKHl1MTGDRPs55KrEhsgUFapdVPPL0YEHpTkXWSH7QQj0aIF+9AfL
TgWRI6bZa0uMcIzHeSGbGfwVrpGhyHsEXCj07Pq19ATPG4KDKi4/B7HmvQvQzU3I
Q8S+hPks+s6QlqiHBKCtQu5Q2Z4/2DFnOq6tQ9s5FXtMqazL2NaK3pqDwBSxqxAE
2gxACHaDoTFlrjCzlBwgB/VdtBC9Lp0pBpIhyPsEewURBvNuTKccaZ33TrUMfrQk
QQD6h7qz5Yiaws/H896MVTPdbvrUPHxjSx3odpqDPVef3KwruizSnPWPbl3hslCd
OkSv964OhKHan0rkRI0A5lBwj4RWRNbwJyTdHzvY/C/2xscbQzZUA8fgfQdtdKeG
75VlvK5giwMZ4730VYfkkDa20LpCdqeZhY4N9RsWk+Rux5W9jzSUvlY413cCHHxu
oDTK+W/BZSq1KH1nD7klX27p7ybAlWPULvYRwmqV4HXeCuENfZEJKxXJkVJGidgd
Zex4adTIE7SgC4E7y6iiQ5Idf8nJDo7MRjkkoN8FenXCer3HZdtDcFc9z7FO82VX
8a/IMldKlCCCc/P6DXORBvrN9gZrkkqBe1z+qaEj/HFJFvuY5hzVSjRvfcokqx6x
mZVw4uqb1KeI/z+v27bQkaun58NgnnZw4xSm4yVz0+TYaiLBYpDUJ/AHtl5DOVl/
Lnb1JytOhTujBs24z5MYD29KC+o3sbaSfHkveqLsMCEfCYZBM18+Ke6kSsZOpDjx
UvHenEBpMJMlwfz34oeSNnBWYOnUpdlB4DYRkEEbRJrEVeO2pC8WevKhXJq9U2+B
hfYjxNIaVWJO5hQKZp8wyZ+V1Yz/ZDa0TK/szj7uN/uVMOnEbpoTKFCi7V69wLQ5
EkTIo8jx3Ld/HPJ1O8vcJuKKC9i13nwsfSIrFMmPoUwquNnBytAHBaaJXNQBBuGU
6gEunr8T/i4C9OlqTeEHRECloKUquQBxlqRKEgE+fzg4cTPNKNWfQPz31RJAqqh5
aIdCMXHEjJ59gJhU3YJnVIRIwd2ZvVbXjPiEmvCpRPK6xib5DXoHw+4PpHupeTmf
xCPe9LydefT/z4OYCNfSfmiqhmSB0SS0EVSmiufkw0GH9hxuQZDdcy2F2/ceK7L6
ronJGlmzd7W2Z0WNgX1fldyL3gqQNWDsC8uIiDBeACGsjtiUtwWFKQZsnKVCaKZq
55iGTF6cpoFGhC8lXxuF1kXv9VdzSZU/xO6EYwd7jPyPK32G40Y0inIl4aANVSDi
rYUa7uwjNbLE6g87ZIcvM69mv2d2Torz4bvxADKZFiYzj1ckSZJkGHQ0CJJQS7dN
64J2pNRXwoeicrK5WofUx++rlUS9C+gd9AQH2P9gWY53Thc7aRiWpeylxJAcXfbg
A/3CohhkMeTZc7NkM3CQr+Zj4fon/KserOKGldXxaod7nT6xRsGRhWS03pi2YygV
X5aDFCK1H5t2QqEI52F3TpkUvpH084nHoIrsgCpVxWGf1ZJ8VmSqyCmbIb25iL1E
fIUm5/jtUbdkQLumVcnF8vYbw1SplAMlAXgUls50LBgBo7klthOKDnhQNQ5pgYjk
w8sCQwWWVVrGo9k+4CeeUQB158Jpr7wzzx4zuiGhg7Mo1PS7NMrdYpwAha83flO4
pBS82VbiRTEITumhWENL+ewp6gIDvJTIteoj66Ho+coFw0dFwsN5uQH7vce4csvW
g2G6mwm8GH2FAe92aMZOMf6SXQhJbl+T6jQKhzawF6huRkRLkS8BNeERXvDv5Kh1
M63uDKh+ztm1bQiDoSCknSxxo4R+DVNzboF/zZ244r5FRe0wkxZSetq2DU1QpEcM
MCThyngsP9T1Eixa2CeajSF0bWy7x6SlEl+/tpAyUcVlmLpUhXKMKRCBRokuF5yX
TzK6+preBiEZY31SBKN04ypbW29GndyS5CN+kkMXglI4buOIz3ohpCr+dpVDOu4b
KC+z00pMbypaiudSKDFnfkQR4YPEg3XO5IrGFT+3d8xWBKgrElUrgoNu4HosmqkM
omkiGTas9+W1If4Uo58wX9YKVGpNaZWxw8G/JX/n3ltwnEzwAcvArm9Sl9lkdBtg
SZUV0sTDSK3ns/brgQpus+tXuQ3rZOv0xLX8XFN4MRcWUj9+toH07AMhRyEB3vqa
RYxfxvNJxDHnP5JXuxQoOyKBLbvburzSghhfO/c4rjW6EXe9d8x+43xy7yFMqiKN
BeMkAWNr77yAMPskZYDfr11Z98YxDm9R/X0NG/PiZPl4z9ZZaiCXHGABygTDeuXY
zmN1bHcY822kgJMGcyj2hWfgHBsmwEyvD0XSl1wJtnA1sqMGh6KkweqHAZVHEAnm
491nQWnVzLL8Z+YbvUqquRHCTGgPLcUXBUhRErOr+NkJqdfGMPGRDawE3cA/cctY
Fci7U3J8jVMbOoMHlqd2csvK7vHUTJJfhPDf3OYiL32NmV4D9y+0p10ouQQ0Vmwe
NvEp90S/fqMJ8G/MdJR3mFIKl6swCvLhVeM+syvzrSkUKTlBRIdvO0+hCQIW3GFG
G0YwtFS4BWoYHIzspMG43QeGEAxIhlyCDIiNuWEw7j+ZaBSRNkMZMZX9t0N/PKkj
zIslxRtwj7KgUEU0b+w4FoDXWzbZF0LsyJvsY2xRlP4eIxtnmNnJL0YrS2byOkv1
wCgD/+nwtHF4yPy+bfPqi6g8XnxbV8rghbOgzoCVdLlCNN3pl1be74k4Kw9NEo+f
R37rE8PHdgD0NmpaV6guSDwMMEqreU9Ag6tUPzm1kyKrVlmPMmNfLWRkiAZslpJt
lHsjPXzQ+QPltznocr/ySH5n3xOZCMa7RTDo7LDV/r51ega25lEj39A1RBQt2qeO
R04Pk5bXBM6Z9hymQoSflPm6tVT83wJq+gVvmjDNLOKftMVHDy2ZgU22G7HteUD+
W4N/N0YOgTnvsGoiu8+fxiJ2PKLK1217NuXSVnsI43NrWeNjRaFR3t/v7avR6wI7
c+eo3eGW0x+RmfQ1BSp5lR17Y01SCW6SJNMKj8fkI7j4bLErFRJme4gFeMETmjxW
MsyUgp/UreoxkNMCqq+0uoSwDuwmBPmwoli0GNlG0BcvLkjCwbJDZ/CrDHX13wbH
bd24e0dF5fEBSnpx/PEWBkkPgKSIci2jJc0sw37h//lfxRV9H9Ds3p8elPFqJhLb
3rVexHcHF0/zYN5yw1fcp3fRdeKhn+YVmXrH/CBdhwElewA1L4oC5tAHtXoQkgjC
KauATLDYPFBpo8XGMRxBQ+gnOyTvpeaQkJkVbqrCfn4rMOdYID246JQQ0n+wOGpH
D1cykHH9gSAFWWzctRfnWG3yS/CC8w+pipAeKQqQjEN55cgpdKIQdth6mfTFrvtj
HNi2P9t8R44U3cLKht9VaNIKxUq1cDBZNp6J4pNv5EVq3vRJK02+eD6JAXpfxoQq
8/RNAqvV2pr+8i9hqfOxmOZSQF7HiuJmCU9+AuhqSQbMM0JcRydr8ZqADRPzuCOm
Ds1h+w0x/IqMcfsx/64u3nyrN7ToVJK9Trrnvb7CIJpEudMTc6v7KvcRiAypEnzd
M8ikSjE1ThAHULm+wmP0WZCAzJWD9sb4odmTmCQM1VaBP6ADJbOLSU0IXMWIfJlN
PLivxI869YoXRLmOHn/cpaGcuWH9cuThpIprWkbeYRggWNht4XPtDIOvM18+2yzz
Kg4wBPSImjzn1R1whEn85nLzsaXWsCYRAeBbBlqiru+e0kWXtoHbA4S++o9+eUIQ
Ijym1ajklZNLBVcXK2OnIWE2vt3xmsIcyKC/XLjDEnYrmbO/O1Ac26suWi98ZORf
rd5zxGz2IMW2dLX0pXNKa40X0y3Bq1z7qN0s8cyDbOgLT0JWUKvhjkGZv//+Y+s2
Iy+t5Tj4vbKiVWmj7yyJi3BIgSDcr+zpAtrRAH3QvXWV9VaPwSpmD0la0vFFwTY1
eK5Mr/7sgWLPT3i4Ac5YLBM5pj/C2O4to8U+LFL5NvB9MCfDrgx9q02a5UrrFXtL
7wnM7+RLgBbI7gObDcvi4Gz3CQk2sTRHhsObaLvQi0zk8vymNtmopbg4o5nFCtLR
7ugnAcA0hSeaMF1J6C/IxX/M4aGHWP94vqEwMUoFVY7Sy4h1HELUGIiFs6IgCQ4q
KDFB8YqLMN/HuYM/c0+IbtPCQkDbGlVu+mv3WSMeVU/66/IECWKZenLHgTK+UNXA
Wu6hhSrlXfWK4dWXLIBvSmzMiDC6MrWRkLQx3Ay3iuH/0abnF86g70CUaSyvd7IF
jPRhvipyyJxPAVzp0oAXjenG3xj3L6n5P4Q+kWv5cC+gwdvxIWWyZIS/cHbJw7Lw
5yPdqv0mnt02+4o9+pEGVdjGGmBNx3ivdPXYyA02V892fWqbv000WbkpGfjapy+S
+XmoS9o+l8fGlRR5tYFcB9PlOU4gpX6h91M+s93YyfP7/zbHJmIOR8hYuZmqrxo5
oYinY/7n5ezGtwFDND7Uv2lPZOd7i7dujjvZOMIv5ifXTIgfFAbhe+567ku+BTNO
7yGd6UBMMWrdBErndkg4xA+lOcIh08JOkh0Hx6ryiWyhAIzhk1AGLN945sqodxBO
iClhucAhb9BZeS8Ni3Zz92Hn7Ta3rElexbisIGdLGUwpgqfqO3lc9qpmtVH7497W
bQVJD2ZMTL5HTxRoTp5IkvNYGNKafKbMbHgE7N1qE9p7NCx+f/u6hwB8Q+gbbB1b
INAkZ8fW8cHbTXK4G+NThd+jCwodyzO5FR5DmE6GLzsPOl2mt3CxgTj0RtUguGOq
HKFsDeeP3dTu3nyf+2GS+EXWoGX2i8DdUWZzjys7pYzrMdpYaYftQWjJ1gqE/9XD
GytM3qyJtNegnfnS1t9utQb6s/7pi4BpoK4mg5pL/H9Zd9ISakzpTEnrz5f6inWl
ajZaIcayCM/7bHd7/qDGxMGFYxbZ+q6FUq5TbJ8iL6Tn/z7PJh1Npzcy1X6fEIOt
v8xn+ScNn5WnVQhJpURZXmahP7S/hEqsPOj490Tn+P0IsL8za5xRIkt8BYRyCxti
3NXLLf4lKiNYod7FcvevnsFjgJju8HfCp4tuP83zU8M7TZLkPZjSDqKOKDnyFrST
Jhk37dwTzfCHv3Zy+ySR/NT/2ClZqUGwdjA40nAt2ma1hJv4A3aXJI5RHcnANIp4
V+S8fLpE801j2lqKxEAG7lqEHBK6pYP9+B1Bk1Z7OkWGx5hHwhX1SaTBxxFEVZAG
JrCAKFQ7a4z8AxjiXavsydoqDWRxGf2uFwMpJ+NIZchZJwMNKogjmaLokP48VO+E
/BFQPDD7GCetNyOXtkDEIxY3wWHxFhyiLKziw0gOJr1/ToMDVBZvf9vDEvm0W8mt
nU2rgEjo4Y7joR73/14bz8ftgs354DDMt4HVywOqeuXJZiLHeVbgjuCykZduM7Iz
PAaMsJm86pR16kzvyV60rSDGvN8aCmMlqZEVQkqsYQKbPATxoeBLwmUtg5minhdQ
t44PyQigxOGbwxQtVx5VxJehfP1aLWK3SnyuOLypmZ4AgVfy4GFoCYm9bUQYipX8
KP6S3pjp3MKIzMGJNHQBZM9y8s+22G/S2yfKgtm9yfNXZfLREjphLW+j1AbrAVWV
tFQVtI/5WTFWVnLm47JXw+WGeKS4qMyeWJQwST/sxVdUgUOXeu9RI/UnPiz1pPTh
gp1+Vm+vqqi1Wu2++WpMB9EyPh9HC9Gq/6by4wmgfLfjxx8mwgQen3nDm3UNixGs
xdZ47RkwcD0CKkVrXe6mwMMQfqndTU4V0NijABjogd8UrQJQ/nHEzIxFwb1E3tYN
cAsufI/p8ceoeYEEHkfif33dkUW02Z+H9ho94HDXh+cEQ40eXcJMcXYmpXNFUx90
3e5Pqr3oVKjg9bFMxsSG3RYWfMnoDDJxAnuPIN3o3rKz3Yf2e2OWGITMbkhdN6mU
9+HhuQ9fyBeW2DVWjVuDK0C6pTh6bm6zuMd4rdQhX/vhh28QS1+b449ZfCcRTuoX
3tgr2fSTrhUUvm8duRH3J0TbN44zjQVuVyRDUYk1wnfFpkNuKxxSlr7KXP4h8DL0
GvGVWmXtKFdcx06wv70DA3kwT/E8lhaPr8fSPEqmgyTVhqlxTBTxoRvq/mgG013W
TWxrH9gwHKQx4FfZ0wP8jRhmnoOLY1X3fAX2DX1RdGFvu8bfMWsbax1y+BqyR4ZP
AbFS2NPfntBUw7NfvErDOZ8WOXFov1IDuODRai+YlgmRCfWuK8fJmDQ7lxe7ge30
J5Pe9v5oV4tS8WbUUq8QvQr9aAbmGP8KVskspplnY1a/srw1g38GwuEo6No6hyuC
5qf2WBbAPuE6740ua55vr4YjJD9RteHxo//IAkCMoGB5t2EELoO1PahSWCkD9QL/
4mfM4N7znCOEm7eqY80MznMlEzgu2Rn2lwE1dxKMJ787IAmq2OYLNtUTBc6hzks7
kunKghr9PRKpqw8dMArRP+ee4bPjYGHEfmEmzgDaufVMwph9cbSDt9EqmyWIoCMw
xClGDr/jKta+aZBvEzbDNA32/M4fdz/WGm29BIWKhD6Kky8CkpuqbjIGPZs2zshe
3ZY/29hU2/9+e0+xxWh90hDYEaXTwMYqZZPDOPSO8FtUnnirc5Ifq60bCJiUp7P1
gZp3kf5r6yItdEZapaCD7WY/zx5b085m0wc+j6aBrgXAXFTevT4HOZJifQYDMwbT
pLvyXbz7xLe2vK0DLq3wJYG064pq/T3GbXE/tLawh1CEHOh8NH/t/mXk9exdwBwB
f1b0CvSt4KtWJ768r7dDR/Jtoro9WF/adNvPHwCA0z9tCpy3VvFRG0Zl0dN7kvVH
3sleEsjwdLAetMIhhZ46XzOnQpX7cE0YRpDCpCfAuqkIQu58R7k9jTE0I5vZsO9a
N/y1OqzGYrAXKMR170fp6Ng3sq4HIIKNzo1rP8fTC6NIGAICm0FyQaMjQlyPIiit
ycGyLqZ5OsNIvDLVco7Wg2Sk0fL0kHUMln63dojohlRWTNRqQEmVVaVpcpNO6Tju
+6RDO1C+RPD48ECTK0DHEVMgVCeUF9DF5kPIdyDNu2B370RhwAoYwKCFlcK+ySTi
S8D553UDFWXT0ofx82BkKcXGoyWe1bxI061iT2Omdfa+SmEk8VmaEg9I14MSVQEM
zziBDBtEg6wRmXPnRofUj82MT2X61LAM6zyNloJoiRGW9ZScyrxNEa8YCYHepReC
aeRaY9Vm0JmZLhlnkbjUd9j3SvQ4xXetanRUnIJh3A1lG5DGhuaiLfupmzKA9jMh
7dftx0F7pJXzIv0kUjiMcEGED2kEXXjl9UEP/f22ul+rZmuHrR8zYt2NSEpNG6ke
HWcC0f7Jt3Jvl1H0EwbpUbIaz1+5B39vpOIS9k3U+1ntvF/mOvbRuM1BnZWYcR9I
0qEoHWIC1wVdgq2HckNWrRcpvfdZc7wTYQwY9U3eK+mSF/cDdFbDMzNGQ7nyyu4X
lx8WI4juvHQ77hHpeqkPDcVH89Ju3XOx+UrG+Us8mUoHZ8kqXgLWfRJp52eHM0av
/Ani1rQHe0Yomm7jJ5HGZDlzlKf2952OyaAegBi410Nn3l2N0ED3SSvoIhQStSLi
2IkjTJc7RMI5NZhf2eetu8SFPr+EaK0N0zPwWJJ7zgWLtg3Nxxv+77YZ6LVr/V0I
1fLHDgjSFWdvqYfr6Bwd5sVQi65OQXXaNNqeIfzq5yNXfTG5AI4wH/GQM+QlpB9/
dYy1bClwWrTGFe3XfkfQHhp4Iq25QD9hnkkl2mqttPoWd76Q3rndcZtPefiw4GlU
7KrHoSHeSHtS4rpVnFqP2BsYMPGD0DfMWl1JQd6TSLG9X1msJ7hWpwcM6x+vR7pf
2LqP16N6XN0y6s8jRxtJU27aMyINWAxECkpaX3li/yXImKHavYrEmQRnd6dehpPA
NW4KQNGbzBxUPoA9NeT4m5Q/eXUht+Pns93JI1UP9aB2d80Ge4haWX6ZtCqE5oeZ
m8PD+plJsSE9ZcHjvqU/8Eh8SJoRIG45mnNsP/mmRNJ1bLvHOHnEhJV4YNiupydT
njqTlUWpshPMAa2ei3/AHBFdPAZVyueBfBhTfNDmjSzH7Pa4pQsHTTCkdk808xIK
EL0A6AGn7HmcM36S6TDW2a0zW2MaMJB6l4wvJWj8ZB+Afq0h4KOCfMLaWU9F96zX
uY3DM0ciUU7oiLT4TGhijM5/5aI2bN/0r9b1s9pSaZk0IV6gx9xfIykRuF1zcs+W
lzMeid7q1aTZoPsNXY/pg28jK8EWGvwpovkuweJmqmi3m/m30T4XC9tBjjvCtSHB
NLjTEZW4SF63LzK73wMmxS38ecve/tuVnvRIp8mG5JjQVicdBjana7z5taydAwFz
MDnfyHLTiqtvosnbIdJwMJoDJhMd/BGAtgpJSaAvf4uc1mQ6Hu9B8GiMRRnkEP68
c5GFvuI3PUfDtBpBTZHfaLHxcAjBwPXVoqG8fC0BKQljpb3t3jlOwK0CT4aozTpp
nxShvE7x1qttUX0fLlL8j7YoZm1iA1ckv8H+gY06KzlhqdH+kfk45PAM2Vp6BD5g
KQPmKnd0EasOBs2uF52+ai1/JzTIk0H8ygCozdyn4JNqccwjWwtdcialupq+UUCW
4Q+k9GU2wHHoJ8jmm+VMw8wOMLszAermvswtIouCGfqJ4FhH7fciEAyQzw4Y+oyO
1P1HX5Tq4MAIA1I4d3RG5DGecppe3tgiXndi8UTjaaB8J00lQKLLOL2VRyG/GHDT
/v/EiNssk722tfwWwYTso0Rfk1PFowWu4LRfutm6mAQRicgDgZ4+yNW2qwRfMA+E
d9uTPmdDZJ2pirARgkBDzpHmsFlooOfB1xreqzmL54kIkZHnQ7IfQmVnRwlZAQE0
ESchevI41AAum+KR9csSzWu4FAMQcJSldnZee5wW0/7TZj5gkWPLXe9VPwxrM7vp
kotDRJN0jRIIowOxJHaX4lmfFsqBUkxSRtd5MpC56yUROwehsDV2wc4jBT7CSTuk
0J5vcA7KhVsvzAOCTzeTYNVKLq4jn9ybbVKkdUnBVxwEaZgUUFP8tdGaguUrq2Rf
ZwtoCSpECkvSnJbd7ViSU3H1Fkoq5jof95Md7KsmXMHJg9FHXGcCLjquSF1flAPu
7ZWemsuUOL9XQLORb4g7vgDAKBOoJp32aSrXJtY3lSC3a41lBR0qSIF1Xm0vmUA9
ky/2L2dthGaLBXfekESKM1Wo5/SLkARzge5blpxYPPEY4We3BJM0BcyQ5eeu3sDo
vdgDXHelTDGW9nAn2tlMm4fMcE8iyuFWBkve2DE0umyWGj4QjJHjmDcak15FoBfv
+gsR2bvqWUu+kci5Avg2sD7JiROZKg0AX63t5/u4KXEtPH7LPYHNnVepFvrj0Rs5
9nnsgFPSj86GOFeF/8sUQUIhohsNgMs9fXmCqFpDzIxiGg4SIakwK/6J2P4vp7NU
pDUiEzkDe057a8yQaV+7zaQWofEuZ5dTD3qq8H/x0ZS5Kd2gPAFLaySFPcznqetD
ZdtBiVJj6eW7EOoD+4y2bCCmfI/FHOw3O77wv49ez2omp3jIzt4Gk570LxkOyaQg
SfR21fiK11lyIAOKhT7aCwckfiJ45KLn0bKaM2a8uYW66gCDC9JlP/14M0K14PTZ
Nk7Dao5rwrcTfoVXyRMNCedHQcE46Ju6670euaKsC+4f6KAP3cK93ia4rA5gIVjF
N5kmfxMJV/2BqjlDunCiaSFn/mhloJ+zQs+6aYwUNa0iE4wr5/Cs7ZjgcpKyt5R8
sIV17tmfhnNHuvlAzJiTMAtlFDueWcUl02gPdEbzB4rN7Fx1Z5ONIq5vbqnxyJfG
Sa4cC6tSoSsb97tqSc0COWAJY0qwBR86IgGNRtMx4PjuCIbDWrN1HbRo3xMtyaXn
f13WN079YRNGyuc9SJglvwdxgOpHkz2QWVSfvBk5YC3VuwvAi6vAUlpeL6XU/Z6r
RALP3n0KvSivoMeEwTube1PHT9r5RU3OrJsr+vhR2fx4CpNKuViMcN7d1CvviEs5
DtyMI4C9rgR0UZVhrjjZi6vlZDIQgxTCO6LrZTBppNzLHSLXVM/9rhw7mMjaLcYD
SULKlLhF+H/DJ14FRNdQGf1giuK7SMBdLDXA8PM/m+cK2LwOY+3hZP5vFv/Ndx7T
bRBzDlpOs0D/QnoX2KMhGe8laFNvJv+0J4Ngvtanq8SOAwWQ1vOwJMtgAiFWXGLL
lQg6rF0E1Gqaoa7gQqo3r+wI9Ex4K/uKl5NmtlMGOcGnL3qsy1hVcIa3/Rw5L0Tt
b7+irQME8YqGKiXoWTZ0CW8NmuiYj1aX9hfHyyOjdvDyU6aavqdueF7GBHOdK0Vf
zIICIbPc2+zK3SUPVsKxyaaPTK9P2NR97elckQcEmTxErd6QrqVcztiDGmeNj4lZ
DBp3aeP0xu2T0dFv2KAP/jYWG5a0Gt38KUjdJnriRHAS3fWZjC90Slej4C5KILGl
RGW/2Q8z+Six/gsnZ5VKeYftLqOXLuYNw3nFM06ZpJWio3hye62NggCzJH4k984o
0C46bYq6FUqbX3Y4/8yS2eukHk/ZSB/fOF4q37C6KHW/08mawXqxvp8R/rkVtl1k
6XD/uggDnz8+BkOpvb/20jEutxpU3u/ZvPzujUq3jNBzDXZnoiIwibXNvT3yBHuB
dR1VYAbT+268sQ05fgHt/gtSTn5m+Bx2Jsc8XZdtvM48wOXAA9iAFq+dH4bqp1h6
9Nsl1VlgvgC1n0mg9x+U70a5NKyiD5fiHTjGKCRcPPWfW9WkR9+UU17g+tmWLMh8
roqaicgq5VjML0C4vOT2LxLYFcnm2hhQmrzie6PaYBnIpwnOQgICAU8QK+RKlSxt
tEWRuzdYrj5Rf6HLRLnoz6uNqsFpe4N9bWmS4RtqkTqaQbV0EGPBHI2a5qzsMx8M
hzWIM8TGeCWTjsGTAP2LUU5tNkLCsnAYH/hyclEiZhVx3z90LGFTdNFKE2ehuUn5
WUDgcZuuOvHFXYhn4lm7FO3Ehv7sMDoCsja/pec5qMSa5P1UlriPlkqNSRFg+CzD
ZW0FwR1OHikNVgV3No6BEMh30cOFD7+XOoCqyeTuqYz9Lvhic8Tr95uEACkTFrhj
RrWhRJA/QfeSpXJuwtQ6jw2f9N3sj7egkTuP/EjjcAOhhu1V3JQCP/eYsfae4ynb
m8Sr4F43DVNk5pWNJ+r9cfqt4Dy55Zps5pYHmSLWTnpLfU9giYf9O9G7Gu21pgbg
fo+RMMwOMc19XcYFLWksYyihfz7dHNGUQR0lMBzLspq3L6HyRDV/UVaHuE8CkVVP
AYupiEXlQ5XNBHdGAG+6BqJxv+mDLSK5IcBIJ3zUaOgZGZd0UN+5NZ4LbyktoGC6
5WW8LHKMfXOX1MRyktR1+aFqKppujxD6bVYC0Iqkd+5utvL51QW6hYEV8klKNuGT
47lwC+78afpQaaHc29SPo+2iZ8Wa+VcjMatXCZlW/1kUIE3x0AxM3EfvyMWonAi8
Wy5bIjYzGTNVdmBR9EDeFDfEoqebD2ufQW8at8H+o+qAoQe+7faXQ9g4FWNasrOx
KuhkhbUmFWG/uALqVOsXQZBu5oRzAs9KDo459A+LGA9garhXKYWRnnWmLeYFQyp3
4oFy974Va3Ia5Mhyj3EEwS8qrFlS5sAcOlLiEJXtcWcfLEd89aJdX40Q3tMiOnRj
RIg/aRJY0V5D5KZpYiW2TW6QAaGWrGd9F6pVrEgyuSrsGcF0h+hgIK1GvT/rAB53
kYMqvk1EAIECcZb3b/EKU+q/2FZgJ3kR+k0cuK1EBCwWyIrJDvGb/1Px/ItMsCCl
QeFpODwss/9PMXlNuEutt+uRMVGdxQ+rR/oD7g3OZfE9hbbjqv5Q1puWdfFIsFaf
WapMcv9Pe5mht1xi+0lz5pux/2/yp9J8mhtPlXoLExcGMRlCKgJOKz+EdPR4ObtI
L6odicy6TPLTgpDk7isK8qc91uG9Wh0oQr3oTh7KCh8oowNQNm6o/9wft/vQ1YJm
pme/xHHbGp52rnxq4mdRI45FwRF72/51799FyPLkSZkZl0yYyIWBxG6DEkQBw157
4bkcJWowv/6rxlGGnQj7nQGlPky8BEqyulwK5Xn/ReBkmRl3TscPgRy7Fs1OPxkT
nebXmxT4B07TVIdICz1/RTadj1P0F4VYAYsy1HISqRTvryvmWeqjcknAPG1l3EnK
6tHWBC2iNXCmm0JcFXOPbWyzg6F2/XuU9dJSW2+IDE7tmHWNAzrFp9L8u7JoI5+B
5WwODXUphf2vR55QUG8kWkAWwegl8QqsAH1qE8QrSN4Y/OC/QG2em344z+noAzSd
Q0taHn3rLCmnfQQ3EherYRrGMMjknuQ37rHQn9ICVGB8d4/auxa80xwx3cYiHG9t
Nh25ALMcLdocAZTAlqxWT/34/3k3mVJINzq3WqTVGr9KU4tLNCYzeSuEwKi8JQVq
c6qHX9RvxUCfMTPlSrVHULPIOh/54M+eGytL41Stn/ggnqYyi7MKz8QjswHqHTrS
cykzG74yxV+oI1zRFxtzSBdc31/u4GjWWyMfhoz5gcUuREWjqi/rgrjJJXZjNKZ6
0YxkClGIEocDUrIiyfP+VrQYRGbWjRZIq8XE3Vn9Lg5UUG6uqqJv5yl1l2q3BZ+m
KF3St1eGveUzegyaPtqG1sxNovhabG/e5Fnh01w131o6bph6IardInSsLJetFleG
W7xA4jay1JUaXik7j0UXKSkR6EogWk/hpsoFVCh73kjVk00Tbtpr/kt61IOt0ZZD
pblALYNc0UO3NQU9Cl+QVaYIfdYMK1mPU87ZU0lKDJGaol8rfbrP2nDLgOBe5wSB
OFgBh3LKeuRLknGYvoM1y6rUNDQZM1gWdE3xIJ2Ldu/YC9OWZa3x1wETuHxoSoaW
YsFZ9hrbtK2BDmYTAk0GBHmoZBsgvlpILGu+kx+yqJjDtmSD8oH/urgaNY/3RRIJ
FdRJr7kbH9PjUrYj4EhFYy+YLjd6bMhnWzIEclcBtoyp2rBj19SBYZu2IK5xZ9eU
bKD/BRzrOKovoqWMkxfIW+yibBG/q+/lrXaJIOG3NYVTpbmTA2WMn7GdwQiPCzh2
JFG7RBgQar0hLe+Ryncl5I4/FrK4DUKWfPPsZthnGnV3XnuFQUz2sg8JUi8Ypvle
lgEbHZT1dhAKnqncImPNG2sZ94GOif7/e0+ZKQNqXf4BIue7h3GSsO/IfSIaXpX7
pmhjBBfKY2RySInPh1fjAXpLWNx+I97dwW/RMbRKfAW8G9Ux3jDq7DK0t1QKhlFP
DJU1vqmt22bmO0oq8ZiHahTZqsJeR+SyQfH9gAGfBXn3IxQ3gnwljH1RkZXilCR0
R6fganl51FMWJV7JC9kTwxIoYf0BbebFxErg/EkWvTVX0dXhEQlzYQmnQHvut2l4
rPDOYNwpWI3wg7o1zToybYXZePSLhuSLD0G0Gb/U1T1Ss75G9MVhncwWeF69pkZY
J+7XP1DKZDKxnabnXohaSddLrcsgJUJ5su6Hf2eb+KKnURqK20NG2KL1q0SbJM2a
BPID+hb5QjYXEfBT1yddqOEBp4d2u2nYRvle20V/BRZt8YHJoTdpUNqk9zudRKXG
BfnAG5du16hhPduIMTEGKzCjoZDJ2YzTB/N8cu4gq6oFsNlbWWSgueksHbfRJ26H
DYy7WRtXolSSOXkKIDMlxPkCd9AloDjJWsVrb2lXROcFqmErkE20z5xbshRJU6Sr
rOmTbI1e2uUbzb3EH0LjlMzfnkuHSyRgwjVpUSX9l+tnrAADEG+haadLv4vUtxTi
wEn6tKpjuwyy+fAZ97LdjaMobBklZeoNxUVEZJlmaHmLeR3Nno0K4ZGCq/fcDDIb
rHWPxojYYtHyxlaMfE6eiURMFw6tPnwsiKooGckAYAwmpDEkd0fX/vvoTsAWY35o
vqWdqxy7GtmxS5uqox5XmKgDBD6zap9NZdE9XQLX2WEVz9ibCaO9wVtuHaPQ1rUH
Jy4/Zuq8av0EBnhp90lToXGFjaTlYQ7OvfMVvgTz55nF66xiF1OmIS9GGxC0JHPe
4OeW9t77kfxCDwRnMhmvQWk3oCo9YLvpYCzoiqi1enhUSHj9rq7A8TFJwv/efw6g
hZga7l5DXDdIQABt/VnEnNlKBVCtbkPs73duqKrh1XLbFkjYNu8XBrBoSz20cB3s
9+qg/DclHuR8cLoxn0whXQtUXA2CbTE4Ou4/ZkOYdw3s5ZYMrEWaDmq5yGD4eT+S
Y8W0Djeb7E7ZiU/UEWSXIpV4jIijw9HaFhtm2JT4DDNG4oOOBGlYlGMUuzZFfKoD
G9YNOtaDpqmmBCQCAEaNUjNXeByC5jcrVkNPrenmFuK4AjRTzJ8I/lSu+Ms73Vi7
ZWasW61a2+Q/76SZ2EBSWWi954miKrsDyfckCr3FGhoWwUb96SdUEmUFsW5CHyC1
JO5tr8RK24hscwkBj3y+Kgut5WC1NisyL1aiSNnHHL/6U8pZKqJ3jR3hgpdkQ8Nm
6IswtX2puu0UkiOov+Vs79CmhoyskJGOVRcBmX6/nk2MJ8bNUpMGxWRpzoaOdnWR
4j+QZ/XaU5P/uG3RPRtotmtorOgMUHSgDaN1Pi56vcVtgdZSbDqagmdGeCY8NF5/
j6w9ksDf1MLfcAlAH7FyjIfdM60OB9tCSANEjYZZnur2HSlAJk43QFvWhsZKa7oF
kt2TkyZVC/s1EtLiAUotEXE+zt5d6+Xe7U2MWnpM+QfzZhtGZ06gblixEHbuS0Ob
DKSQLCw+sVv2Z24oRJhRjweSOrTcy8F5GDywC6vn98a4xD8O2fl5o4Tm4y5pcDEa
Awaq7t/s945XqHvCF8+MOOXE/Bh2L3fy1n9SsjnyRAGM5RLJf+FXDKcvOco5nrHI
/20sc0CAFSbAhQLHVBmau+fte98d/Zr0AAK1xuLDpyoOENBb6o1q5Wtn08h5RnX8
N5naqLMSLFZtrwjF5OZoQXAvFYNH8ypEaCRj6i6A2BowqArEUyzOQPwi9XF0lTCc
qwm5slPOGMb6aDvx4SODzt2I7uwcphq+1c6U4ilfNPb4V0Rd+sUVdgxsCurLvZmJ
2RT6YXCymBrnv0lM1T8t1+CbYwhBnyIZ7QMtqQnve/uxYn0Z11pObz8JTtEdVzAt
VgO+L9djLRbwhxPz4nBOqet8BXpfNYOmGcK7RFitie1SITOPNVkrV+6xu1Hszucb
JRVCQv61SCpAmcw6HSBVsMWCpn8QaqfvFmJkDMSBoQyAyRHNJzJUYyOtxE8CKgD9
LbtToVBZVKojGNf8AJlXu3/c+lcqMVjKkE2qlQzILKwkGE6At0Fa+qOm1FTGEY3Z
MuxyuIJxfoDVP/9cRl8qk33YXhJL0DgkBR5OX9f+oju410A/vK4emxlPeMKK4I2g
/SuegcOCMjoI69mtPGhP7yLi4AB/JiJXuLqHo1k8LwwnCA/1RveWetF0dmNoqq9G
6I02kOD59pEiAVeESMJjkF4H8ii6jSPUymIu/NmNnV4JvfzXkpIW5mtRKs4K5wvW
T6C6PRJ3XA3fWVODbValkJoQLndh3pd+ZSiR0oEM/uvRBmvxV5oAiNpc73OWV6nq
IaWtNJmb7gcwrtI5ui/xkKzhuFwpMPpq5zhSTxG0N8pzPW9sF8c+H9qjF56ltdqw
mByfINcgaI4ojJokKs3ENCpFecEtRkbnj0yBtjbSlIj+Sb6LwhlqqmCPC94FdOH9
AppJfrSYZLOOgy0tDBxYSFszA4f0ecLCpPl6hfobL8CqM5tclxotmZlajRQCXC33
mZHa68JgLdt+Ja2sRkmyFKi7drqYqZb01Q8uYfZnaf7AJsS5mPwfv0/2DgpH/DYy
rpYg9Oiehd/KSS7EGjwbLHKXSuFx6GD04IYe2r1ApDUgFt7um/Yzdamp0BYutGY1
b+h+ZN+RZ5RUKdCGOU58+/gh5JAHlo8sf4N2ptDqmynolQtiQ89yx89IWXgbswUV
t9gG+dqoGRSZk4bH71sDecQPW8h+RYadwElBwbCkGcwnB0mlMK7yG/8O4X+6CwOS
TRCSKoiganP3epgwyBgd0Irqs+VTp9qyxIhiM9XbsvncozgQF4wojqFYcUtTO7ST
CYjPoGNqGQewIHXox9Br5YLHxwLH4VNTExlKj3039evj4tdiM1EAstZmc2zv9QmF
LY8znCtZS5Ysrt49Yns+8VgttALPuEL/gaK9maqj6BF/QPSKqfnwTFH8w15AfqRk
5TLTGSN8d8b+DqhgDVVqsHgZpV5w1CtChdG6jXOFzERwAdAH496wF0VGXADVq0lB
auxpEVbx4oxw03tJpryFih2nX0eFhYAWRqtI40yXD8Imzl5gojI1x83rBHCZjnHm
6ikqNMmuorb4y28QHdZ+HTecVoHwSwIrafyfCI+elyIFe0MIX89uv/gMYJEsRKFf
0LybHM2QXC/WBDiYZXC3n8P5mx+M/8EaCQbR/P2SVoOZD8MQi0/2IudQQp3vk7VC
p6ljuQgr7iNBrIYYmsBuZ/6L7uH5GaVRPnP2skx6olrKugsVj5V/vHc2jbj5aDxH
Xcx7ymqghAWaP5OcXVGm1bbKy5YKDihCoK3/Fg47JxoZmUh1I6GD5KZ6LQwZphA2
QTvtz7NeRqnrYotmvk4zrXlSCF4QAQqfWh6+tSaGuFWIBvsOwV1YNVJPkzRJOTAx
nKFiJuU32eIgsRSyNK2iHzveFb4y8mkVDKBrqHUmpfZwXrFRfmz0ZeH8MQmiDqNl
v2LpSbO3p4FAIZ8WzVPJdQ8f1u/dWukNMRC63nDk0PccuKOT31JHYY5jXXZB2MQP
vS42bC098kHlOCyOikveR5Pqc1mYZFUYzqMY0Aix7v8jl8zNpmX3WC2+XEck1sNO
JOAtc1OZFo2RxiVwIW4nqH7lIXw3q5FUggAs1YTSlh6sNWJ2DRiMGwoTNM4YXmBS
S9idnK58poXVRsdtLoe/EAiGQdMaMSSY2f/do/k+VHjFBqZZovtHhTkAfwB1slz0
DLU4px6wrQy3szLFg72aBL1KdmzT9zzQ2bCnjj3TIOChIZN9j6f7qzQ6YGak9EBr
NZzNNVdLTW3TxJ0Bmxux5uGX8xHZW/PG1voH4sToiQxz8xuhCe6gKvErwoaUf4tb
aeB4j53cZwxrxoZ26D0Hj1n2+SrI5v9LFPe7d7wFm6hD3iMzoIQ+pnyuDAauPjfq
5MFbAb22IooJ+K8etd3lxd1uQDg4Et9FsGLcWkW9Exv0jRj7Bt4ph+ObcKFHUeUy
EvkNhXqAGalEmmOmbuMmPulou1lkF7xhIxIyzLyk9E5ZWvXvk9skx4YGimMk+eKi
ljk2Lp+rmOkaq33Zv3z39DgcxIX+Yx31zvspIqftNsEBE508X/3BMJfZBi1MPS/Y
j/XJXxFwbBjSwjJbrVU64NVGYQhUMzViMvGoPDszrd1vRG+L5W2tGJDPedhErmgK
7YZNVHlvVnLjcBuLkK2AY8nLq3Zl1N1QdZIy+15x58Kk85qgqkA7sIsZVmgNuTwa
70HM7xjY6KPC/QO/CNhr091dVuFgZa4R6vb1oX6Pabr1zpTxtpTDsHxkYoXP4SHU
ejZof+3B8cchFKLkLn8OEHQA7XLSyJpCM2atJE+oibDmeM/VE9GfuQS/ODbP8v5P
nbXwxPTdwuBHq4/y0rq7vsK/euKjsPNsTs0g25GpFDGkjQlz6nHUWWDkKci1+ypT
htftigiM2bR2QKUhugKeio3FMMJYvePfMJvuR/BMuMphQGOEoBD2CiTlS19Uh/Zr
x4xfjXagkDXxMmUSKPexeXgb9CW69aoWIK0WR/TLP8PNZ23meUdyzNOBqqSwPF8+
pO3YbXWzV2MD1KLx7vetODpwa1QaSILJbwW45qixBHAi8BQvRPn3EXYdPdQfyHMD
OE+tLv4cENIXAEyMN58y4UC+ACeKG2zcv4MvNksRmXHrSupkUa4cTBzDXpWX5IA5
uJ1gOEwu+We9n7D5jl72HSDwLiwfOcBL3GG4irIFNlVlb1DeDsFhbP0IuJomr5Rq
X4xM5zypDZbFvsUuG2XCkyngYflTe8swrzIVQ43Cgxa7/P8hMib9sr3Ubx1jimlV
r3EicH5Tl8pc0y3G1r9Qp4xZs8/K8FtMv47g8Nd10tj8y2fjtswxXqj6ppfQcC1V
qp6t+oVtxtuXochD7SjQHs7UM6oDnRB3gOh6eyuwPddcZZNkuvNXCIYr7DlJa5pr
W1WUeTReAgD02rB8SMu7948dVee43tG4DkazJy14sifpSk0Oe2S6PO1wwYSBByno
m2GlzD2BBBPa3w6JrvtAsji9kpYC080f+9gMldnkXjz11dDawEyl0l2DH+I6AbS8
KKTw2mRqg86Q0a0FOF9759vd8P3j/SVBEfGKm6FRC2TDoju20aMSHPKCq6lIsg8D
hazdQWSEsIYWKEzIN2QzkCOhOyv/7dwixaj0haZmMSpnCvCkWN1FWVS9JqdVOtUb
SPjyOiCETKY7TYEzejaXScrSmAM8Q9E16ZKXB6kYfUIgmk0EAPh2agINe8zSfKY2
1t0uz/kL4b86MTUqvXV/LHgQv7dN8uJVOHXFnqExlDcNqKl52vZD2GMK7pV9mCBs
7DEb5a5m40ZQYSyqqdd0u3nzDXsflX9zWFc865oJCXmciyuyoFdkant+IXOuCbhr
5z5l/kUWBJ6NmrgY0jjtac1YazonlyBf3tdcJjfp7UoaNXkLVEjyO//9IPDIVWed
jXb9sIS2Wj14j4xoMVmJ2CM/EhOc3L8sJggraChtqixwEDZgv3FvXilpYAtJ4ezX
bOJiPttNEWw9OFOSbeyCzyK6FlYZpUYFx74cgVi+xzqHWJIUmrI3tDN5vZuPQ2GV
Ctk07sqcN+NS0iBfi6Kmxp1vOPZxNVHc9JF2rTKQ8BCUFXI8CvgsJYvmou9sVDLo
qghliLMqAXqa5R3JpQwQ3kBN6VY5qiWOfBB1M2cWud9C3JIw+P74nGOhwBznpstA
rQUwiF4BDqkuwsnw9wHHWWJsz3pnJZJobSNal4AFvgVwILaPjxzyH88dxFWiU2Zw
S8Aqr3Qo+IQFGoq+v9uOA6SKdHG7BdSBUY110Z6tXehvaQVOB/G8eo6BJwfcjW+B
4hZO2Re+5DSNf6Lc9XaIHzQpJhRYQkyAt/IchcXAkzIFuFzWLYMaYrFZxRktUKm8
tQFbK0ueddnjKjtHb9jJkFXprna2SbwIFAWyw/6C1gZP9oac3joDsgZDs2xHcENK
r5V24u0eblt9U9R5w2btCd/pJHQQ6ZQTreqFgi781d21P6E5Kv+mizYATABVH7T7
3qFPH2guQ+smKpDaZGIY/K+iW3/ijmzm+dUy2lJmZS16C5yjsFnWBD9j+8DU6DgJ
wITSvVFirHvM5nr+6cgdiNwC67xOQdW6rIgCr7+TqsLT7oLOZXLseCwVEtXsXPnp
OthYxZYp5p3kXRuzeMZTCsqZgJlTN8E+R4phHWS0JDjLi2lk7XmLlq1J3qdSX9PL
FnLR13NJGFgqfzQeRNtG9X3kYLTAZYUFr10y5XsWOXPRVgzdO+qIl3F996EGjBmZ
353o38L9d2CQgY3budQeYTRtQEBMNzc30wX+/u5sNaHnBqUKNxWDsvr8qypxsbAa
ZHqurG9ivk+lYpp227kq7BEaSzenAuWfj6lT3oNYiR2ioroExVufLLO8g0i9zhGJ
ObJQuVnAEIsbqOOx14NLJYAv9IkqyZdTMvFokF+d165J4uSM8yqzZBqOdpA4DsSG
omfTdVUtIOoA/+BLoyShif8Psrmf/TphD1z9uz+6Zzo3AkaJXLunebfqlWlMg5Ew
fVZBMBzk9tgD271FcX/hhzEuO/LH5Ypb81sanKUiTHClmsClGsOjkXnI6WsrI/W7
8GFrCykWSbi3bpNpOVtaNiWnyYQtGOFhM1tywHG0YKgPXJaz52cyiKzFmEj5P8TI
FMSIb1ryyW1WIpejq6KZhEzv26sdCnMcgWMmHPOIBMnVpNc4Kxzuq4QCoEg2SOFR
aR7Qfrj2Qew2G6RyU82+Z2hgr/GBMQRYkxesOva2F+k6OHLxcmF0q0mvrnAj4JPa
cOfiyJFiwLGU4tlDH+JoI8vsyEFuCFjTWa5aipjLYbblYmgtBxqSzziIQ2jLa1xj
2kxs9bEk80AIAnuxUa8Vcyn6xU83CaNvT6CSIp1YXWPVALmcColfVvydSiJE2Bie
k+3vAlmUGh5Dve3VHgeze0QIzLeMjaByLaqaZr4BxAx4JQEY+0o2tC8VSrm2wKUr
NjGmVBE/0Xv9mwq64geeKqGa2qFk+MwmDYhJdXe2Ot83wa6Um2Hp7T3obLjmYeys
7Sgtk3N54YWtsSr7E+oNtE7Hw4xjY3PNGuWvJnr2mpgYmS571r27Xm3Jy3wYEZay
MLuSsXrg4txTGesm2i4eOVcz8qcgFxnrnCvzxokBoFKR1d8ts2GScAO9eaqb0hqa
6phmXV2Dbnv9MizSjtFvmTO1CpIyq8xasPCfIgEJTyurQYCM4fTlRcS2ilSUgKlR
UHhSOMD/Wdjv8/dgpNShpBNsaCvLEHGU2DQgP/OcuUM6/wiNmkUlG3MzJoz5QpFy
T+isoOAVhgSyQrXDoOF7C4sVsbNv+3+XZPIKXoqIspJoqfXcFHqHMFd/5T68ZIqU
JRSMrQjTOdhIgQE64CQ5yjX+ajIrXGGHvVvvGEdbnwr8fOhyfAP5DZ7ExWA6TatU
M47rYeUSsT4bxEHa6DAddu6uTpc/hMHqBySCg6qdQ1BvKvouvBfxFMPR36HsDxSf
QX6IcB5dE4ABJaqpBnPoRigV7F8+PFwVk63EjPAn9GMy/FiJLYQ0FdtN3Bit+1/R
MBVz6fn5xUgYW8NKfqQMsaMrfYmBI66RkM8HC1PSPlsRfHNL7b4b9WnqxFg3Zup5
ZachrPk/tqaF7AOJGbRCrN88SDrybETUGNDW3TzI5KvaL/SzJ2EWCiASfbJ1x1Gf
i8xWU7PY8i1eE1E4TSnsbfdlCnDNeiBw0gEIANm/EwlvpY33ZURIF9KmgUDQHuKq
OfZg8v18smkHtcdRTMEw2izhOQn2QUKFAFddEe1TS1qc0z3dAiy9NZRECKGcojo7
N/w1qjmZMGVnw4bBSnY4HeyRCP+g1GcnBvn+F47xyKx3bisGAoNNyGBIMXBbg9wg
eLmP4pf+1SeIB2Tv37hjihZ6bNXKPII9SAdKdC7YCvkTCBWRiWCdhIm5tAXGd3ke
sg1PQFatMbJHU6Nwhr595+Nhu/1r96SQVINHNIE32rAUzW87aD88zJh3NKOoPUY+
+VdeXxbozhnYJXWdl33QSymAOBVkFNUKMTUigo+9JhtDoh1syYGwdLX+BstH+JIN
g9Pr5IdrvWzInxWMx+UZdnPM0q/hJgTTdCBB5usmrCCjl5UZ85XKILT36qhrGK+y
65vTQWsVaIrjn8nBMiPVfGChVvXP07+zpe5r1ZQxrCdVdtWK49iWqPWX0XR9yKTO
Ph3aguTAq7iVcBbg18hw8K4bh81CY6WKBvhihpyKYAegYZG4EopQWzh7Pd0+U/WL
sG3qaa8vXLAfcyklKSwpPBxx4fXHACkEC2Z/YfmjPA4x0VAZ5Qz1aAcqFjR6KBRY
L0EUVTVkn3URQa7nEiSNSGsr5I3UYqZs6euba+mTnUFaaaZgW9AuUBa4Scuisxb7
31lgX48OEU5D8KlQtdwvyxghO8qfM3iUXx8+VjGo1OAKwWLyEJQAHzeLcAh/6xER
hjJhANQV3ut+rWHJ0PhI9iGWWbIUnAEeugp398RvqbVqmRn2rZj9QcypXs20KODZ
9wPSToa9KmoAK3H5N17SSqf7rWzegQ7zmhG5EO9ZS/XO+6D3hy58s9R7xbcONzo3
Y+6fPdoPOddKXZsWxUfTslBX4FtHJ0BzOb2egOpiLQ3xnrTCug8vW+7H+Ye0deRf
vBZGAX++HYw+4SyIyC0IdBsc0qJebQPZvYL3bNYaVpPIAhDp+BHCYF5l7VtnhSM/
lriAjp284+pAxSUyTlIW74I0oYBtkVIrBlUa9J8GcSRjL0xQ8rZUoYsAs8YQRzMd
x1yIm5wZswut2uBd654UDnOjgmmtZ8mQv/cbutKn2/C3jbmZvqjViXS+xJsQggw+
aP4qKrhjd2oVe+fg6bjUrrTbRwTN2qqmfeoXSJ3wzBYspLFVjVHXturnX/7l3MQU
ywufHackPJoZ6XqoaE4+z6QLSSX0xD4DBvMRPZvuTQL9Y1/T5in2oJPBCBqb0TBN
vzSLhuJS84J9y2otu3fkIdBcdM36z4Y9l70USkrEu++nQ/9Jl9yOg9UR+vfPfyIF
/Pnw+sQ0Q5BGusnFyz5g9Pyj2CO1Jzo7FMMsfV9qyLKoFRvttI4+Y+dlkjPCtThV
L4qxvj4pS78pgEdpX+lwhv1dFsZZkh/PPIyacK3E/P5ssAmzTi5gZ5KcP/tUg+az
n8l4EqnX3XlCm/eUSRO1IiIyz4TXxuRylOaRiOcjU6b3ZSW27IunLryVxf9etI1D
VvI0QH4XALuDiBPl4j0JsaP+s+BN6+p1cKiUmNm93Zztqci4EVR18wnGckxJLSGk
0IilhfmYFA+mCwV7vgV1iz3DhaTKdMbxO76ParMk1mBpuPF23F2O24iTbk0oq5Lx
2qzM0JFsj1lXYle4KHQUbmAFTOztERItWpsa/FSO8LTYbh+T6EWY+Y73hHTxROz9
fLzSZfpQzLtCAfKB/oEvueRtrHDlz4mA/CV+f+DQSYsFrrzUtL0ETKdrL2+k9wAL
UXROs+mRaRzomMuetxNcndxrtKJjJqWJOzFC4bMLuNUfiTK9RmvKISe6Ijlr9sbb
BXXm+yOXpm72XXOZj58ypgAJnrxS9jLiidpFPUswYElINoEXS4pQNQf+tzuK0n+x
k2uFVkXMjajxejj+2WrJk/Pm1TeQLxeZ5w1gVHykrqajQjncF7wdFW6giwZssNgk
gN5fm0VPLWSu/GQ/3wmh79nfNO1t3OgND0V793cg6tt3kGMZH+75u39zfmYgIOIf
+HQ3ySvOfdr9JhR9DQ4kXsLxHQnJgoMuqZ0QcMGzrq+P+jx9fPRbkVPxt8xYp5yI
XSWG4BSzdUO7KGeRvNKOjlfYlG9Xa+9awNtn/BIjEB+n7CYPG3XHlqqau6DwmGva
QQ07O4coJpzLpc/5iHaeWKuNpnz6VYXEWad46EJoOHv+iKuCleOF5w4bVouT7Ulo
/6o8bK40Spi7aJBza8DonC1mcoB4poodQfEb4Nkz/BUALmiykE9JDez5qb0LwgDQ
eBI1PC0Wo6MWGgOHNfIkcvOXrlDxsAIoJpqFcHamxZYfzm7OvCKL8HPTD1ZhTtVS
URv3nylim2ZcN5kAXUJlBwoRLvfPLTnKUNQRBvlngYWGrqs7JRjGWn1zK9FvOLGs
jrJAboTky22nAYusofwmx04O7byqLSr4y+Kp2IQ/to1+wop8dQtd1MClZjaXPiOt
uWzmDGDRULHWHJPTE/Q3wobQhiP8yZgBFBtDlfsf1QHggJD5iOmuiLEDuT2slG97
qaKWKoL7k2bOkUPHBFNoayooqzbgtDzLgoPVeg/nhXYGzS8+yTWLYt+tPC6f109Y
YEow5BMmbnGRMl4BICKTY1e8vBTeQG2aZaqKQQnXveAliYi4lOVz7TrQxDVVGgGG
6eAKdaPlVFVcCGY2X5O4wVgtMwV1aYZcp0EhdpWUdHLXXiG6rF/XkpE7wv75viCP
6r7mnH4UBusm0FksF+OnWYttReQ6aeeea8e440N5C1BaBHXXe24bOcRGV66HgV7w
dEtjFfehdwzvLIVCB5QgKpWhZkjvE75S8XcOWYXAqR+I/I5pvbj+YD7ViWfj5B7x
WLfPfWf2516j3oN8+Ofk43HqoFnUWjcjU9es998VPimgSQWv8c+zoBg2Mkzj7Dkr
yrC8GK5cwDDhAOUq8aQCT0oZbOprOoBZPcfMTpPY7+v6I1CaPbipLp4UsgcULCMd
opQoFZs2Fi3rCbFkaJkNam6n39+OtVFrd3qHanMQ5vwOARDSO7SkXHns6bsgjyXn
m022dHKECNjXHVYcqbWdtixzMnPuCGzYT9S29zk+/oC/0VWTKuPSsNTTNvHctHbh
GOIzfspQQcMygYyM4RB1wulwXnJoFMbnp93gHSq8gPzUSuwOlvL89DOeHSI9ut0l
5hzU+XIp3w+ylURXQYdEuTKXiSTqvbY8y74mwhQHuuwyo7zKO4bGlrRhLgrYU1fT
hsHEIbiCsibz/K8hs6N4+8zqlzmZKZ4cdvkL2wSUMctX+lttm/TdDKRyppDYHyZx
1lKlcbshxuD4IkHHW7pwApJChl6ILlRnUWe1I+YK1fR9KiRWUF5fwfp/Rb7PJyKe
CBNf2ZDtmzJHd5tCCoLW6Kh5ufrOWQ1211ulHeTGQEVRJG/0zab2SR24WdhvtZJ1
oM+d+bAbE3An8jbuuZEOAihp1aBRE7DzAhmyob4KJYREdAAERMs31CRBRFdzN3ox
qhWXlaz6QGdezTgCz9f5kOjnRVzo58ip0aH5caTdYymXj5EqeuMoaTwRGxMCttwO
cOSDo0qZf1XPG/KqHsPXIgvOP/XJK2KbW7ufnlrVTQF5xLetV9biXQ/88tihxn5B
LzG4atJVxA2c0fAkUyAIwq4FSXxoHgMiiEB4fWWJmuSQKvgkmpc/73IwrhaRrkJ3
rK9w5fBjuIf7mZRJJShcZcW0/FpOb+bsWXeH4Rxj35pnEBKsxJw5aiikOgqIX+67
OJaZOmWmnwdaxamRUx11w5TioHr2VMZu4foKpd7iPRSSqZxApVGgeIIb1F5Mubd2
EYfv4vfVci1n2l/KNbYvgMoISffD1To/nL3IP+hB9Jb95ydwumNE82IDD7fLnsLm
kVSCi8MDNL/JDg5/cEmubFgQxzX/s8qIKSMewpwPZ9WSicio1dhbudC+XFtJEkwq
ApuI+o32vquswE/u5ZNblaD7k1JgNmJqhmvclzurloSY6McwWcNjeN4WetQx7r76
hMjfEe1qZZYJbQjleffknFZKYl+ovWs0q87DyVsrmvbZUr51Q9H3FY+fKNqTypJl
XB7r0hoo30okoHz8xqaDCcT3EUItKzNSH0745urXE5i8PAYEsuTD34W1L0dSGq+o
hNLYOUpqCYvnHVI34ewKrG4Ny1akRPniuO0im8lr/3M3rDjeb/xUwePrk930BxPs
FmSxwsFRRzRbJgKb2XdlCT1Wx2uDImF9mOapci2X4v6Ihq0XQJPwz73Q7RXg79Bu
arOILjCWZ/UAJylgdgRh4zpWL0YnEUduDq6Ix6CUleeRfEl4ZmZWVj+2efkEuJsD
qzAK6XnX4VYZ0yC4bC1vA5CF7I5GrLBqUlDqPKAinXchJpnMiDgtcfLMEItwPeCg
pE6OiyASWZunEjyL8nHALGS1ew3Qg6HCSVe1iLuaLskUbK5rAErgCWN2eEFp9Fgm
k6u5yTqnQyqj8juTvhQ95saz2LREuuigLTxmWvTCfArxO3HaGRB+0zUUiaEBoHH3
O0Wvm387lIomyge8u9F7oAuukmKAIlgCED7tls8ONAKDRtkd6/GnlXC9NcAH75Kp
twUMPMQL6zB2SlWvT2zhyulMt60he/L8ehrnCdDFrYRM/OEF8uc9UGAm9ad00ZSZ
4lLBz8MECIFTzeFRTuMZFtplfZ/d2py3VoF3Wu93u09Fhw7JethYdw14j1ONN96Z
EcdbH/s7ktxQpN9fBsxuTYXNmiiVmx5A97oAhMW8eo7QBjcDso7inGFEF+ZkYk16
d9LRkXKsYdBJm9DS70Fmw4nE8QxOHiK8tH4auUHRvR1R+4iAabd+4g3bNuoNPesX
9A4tUCfyrxyCAGMPtcDvBpxt5w9CsptrIieUui2+6rSJ24qyGeuKkpIEhF80xPhg
JAnTsKMRE4rPw77qksOCujBNpXM/fH4vPaw5Kjn6S6kuv77oOpUdlpgC4rqdNnCO
Pguue93rUptqF0MPSGtK0bDKd6cc/JCjfnJk8/EeGLJVpkUbh9EDugv5Siz/40aW
R+G/sdgzFzcaUp3SR4ILgnxL9ynQrhjqL0GKMxtH6gDPDcn0StnNjvGNgWbButyy
K8l1/ke6jUBvVUHM8/FB8Y0Y01zY0+L8wKf4MDTuxpzGVGxmkY9137vXeqjjJUA3
T4/73gBUhTcKsrPsFXMXiizvBaLW1E39La/gg8hB+4Hk6l35QsVtgl/1IGGcU9Zg
C5ruBb9YW/dnsnznZ49/Og/FIu2Te8briYod+gBpI33XDN4WypDNs9y8PzIHFBDH
VvhdaKVYj6jHuJgKKKx4i1HDLmYY0hldWfsmKIljuAcFJ9YwebOhQdN6cfBLvcd5
iQmWxXszSWIX+VMPstuQI4DUssDxNZO5iJs06oCIZ0tkkfaRdV1z470OCGpu9UtC
08+CHz0PsAr95VuQm4t9pZ0OAZv1CESS0vkWQZZEM3e1Eoaum4C4/3CNNVzy+zsc
DB1+btdBHVgPR7/bsD5vZ/aXjv3Udj/QzW+ZXyS9dtHU8LIxzrgztiYxrVrrJu+1
wUEUy99O2uAZoX9l8bksk42VSb8/ImyB2tMKmAD8WD2Gul+x1+mM97ilJwY+iqtC
L7wQL15mMvRwZUoWvxW5dPfYwY7ADPheIPdO9YSNSXxGctEKiv4ocIw3t5ZGERAA
0NXf9LPu4PthNzoi3lDijkSWXsQNlfZ349V17OZasS3Dp8c4Sbkbq68nvygAxTKs
Y8/s5raGiRULJbBkZ3Sub/Su+YC6k/32q7BY6VZNXQBk0Qx4kwk6dpl3AafCf+Bk
1uEwCxCLjanT1l3BSq/5ejyAJSBk7q6y6/ndpKidoSXyxwVgkrdBRq52iHrUfPub
I72l7R4BmpY5YLB+5a/CcSL90ysazmZJcy+DqEQQhjyyLd9JQL9pavecr6F7SY2N
uoX5kpqnSSMD9R2FzxPVogsKA6MC9E44iGl5NTWRB8mIRnecHzVTFjntZvaeqJm2
2X613yeogBZGabouC4dmtKZScBzwSF4YOvAPifbxM8dVdpFzEwk3MqBE8ws4x+ts
6X7vJjEh6cIm1Kan4aaLoPvR9DjUMmh00LP4okOW43u5XMdcdC2nBLJr2/rMgBAD
gMnEnLGmXCTrVoCXlj+SmASNJTdjJV1bjTlXCKHhq6CxTXSnXhdc68K/L8gT/bLf
WeJuXPZeUfL5wf+EMUYH++wGeTjCfRNsBkelUwjPJU1XpLtTIDjnPtsJ5IWL08lI
ggdJrtbRbrvyXHoQBQP/0AtupN6P1OXO8u9RvCR7eEUwGMHMq4gqUCEa55NkFpsF
cGH2HqRuiPBaTJvEEOsHR5yYc8TwKPXR0ZQ379ksLiB8+GKBIOtAg8KQr1fKQehl
8UamYaib9w1dLvs3mjVE36t7yRz6U3cqKxCW29v/V2REaZrUE3kRMvcLsxyg8Lzt
Ugoia/qBY6boNVsmQsw2CjGDOn30t2jgLTiaa1eXmHwllJOsT21zbJKtRFLbOTdt
4uxsmSVQojo0q3Yb56XsNOs11zHDEU5kFlmNqLL6cbs3/7nTdoMQ4VwRFbHh1x85
qlQRwwBQ+ddds7+gNQnCQHnkBeGGUzycBuTOnJGbv4w1D3o6WQNkswqeRpPwAf2K
pjJThHU/5dTfEXDZz0k8P2Z3Wbqs9HIr8jMAoV8NzPROBLb/o107jt/JdsiFKf/I
qWgVlLx9/QP4XdvFTHTPDM8HIPSJjn6wmryTOnHiwxxgmJ/cUFeRJ7e5dmkVIcAE
jjK0U+j9+UooQI00HCtNc3FhAsT886pTTpIzrMZTqv7HU2/cOyzkhg1RoXP9FOCe
ZUChMlwJryU+JmlzvEBWuWBhLFpIvoF1zkuPjlgTL1lPBisByy8pDv0E2JMfLvkl
0NuA7PvmonYGkfcFXM/6728ZoGURS+jy+Gcwnb+l4aRaBrCrmdFeN113Q6ydW6NY
3Ero4voNRm+ARHAk8Aa+sR1Tw54cTl2oTta3zUfl+7eFfLXRyJdPTOHsTxJvdk92
25sFBft77Ync0UJOlzKD+vRbWAJND5nBJrBei+PoYP2tni8yWGNxSbIP0LP84mzX
EgATkiAIeUuUELmqOoP89Tcb/KuKKu1gPi0Sx2VChrfapIe9ymFVuXsf0BnVQPD8
0oT9SosSnHmANas9GORpDHqvSQJbfxYlhP00xf3Eo3B/vrHU8YgkTd8FSZD0VoEz
KFFSxn6f/RwvStE7bO6tynx3yGTuRQdd/jLz6H7cAZSgnaT/DVYD6EkdxUDeRQH+
yaEkXMzWXLahwvnJOQRRkpsrea02DAnFkgbhN9gSVu7HZJgTwvTdRNTo3LxJwD+p
po4Lw580D5rvb9Y5esJUb8syfD35EY+9dTxfsdLAegsPaVRBRsfBEiSgw8BtPE2V
u1xX1Z09W+dKwo4f4AupKWfwYOcvM2hPIXLR3pqXSlCXfegex3GyrXwJihqr3WlD
9bnIPFAwzaPpIDAfk12KCp3FJCG+dOC233yhh5DSgJBYk9ndyzfHoOGqkmR5Clhh
BwtS/TYEzX8NfG1vY46VYlol0ZFMdpvQbPQirX+Z89Fa13EBW78+VdmuzYCNaRwR
72Sb3QJxDx0nS82JN1tsHX/vMJyF+b/OIZrWS0v2A6HJRuXwveg7mb7V6O2jidOR
lkINEpMmXqONkemZ8Z3qh7giRPqeURvLUCX4jEaNkBm8XDedv+wpX4XxKYwd9GS6
0qUB5TLQ6MzMXOTLjFgac0AKhUb2wXwJ20ufU/t+bA6MY/CZVyu+DPpf4H80mW5W
NuMac7zHCO2qVksnVayqZb7GoTUuLJDaB13MAQSBhs/QAAr6xQa0MXcoC2d/af+a
jIdvYsF0lvn8PYizi5G+NbdDOXv7cZBjDK+pL+jeqWnyibBt1euTGExopzWm/PuL
6zt6lsrN+7Vlv4qeqb3tZ7/2cF7JR9/ostnybVuKmbpqQqLR9SsVQDgmV+8+RG5u
eN2zIWNcj4e4M3WlPCKGUFcJjDZM5XRdX1vvJBiPUFKvm+X4n2Xc+mFWJD0Gs7GU
wOZIlttyHHoI+Ayk7kw+PTagFt1i2zsMVPmrhO78Zqle/Vogz6BNhDJC/3jexVFh
LeDLslV6WOT03qd566DY4ufOkFW0rNovUWkyvV+tFZ+kLVNVw2XNZCtJ/2/n2MSz
VjdNbEr3t1QEzCWrxLKihj2C9smvd8uYz4lOLFE3C8hMf4WhEdwygQt+eLseYQOb
/SDsndWs1875w949/lkLjrQnGd7At+KddODVxkyqFJDZDyexWAvSmNIMfXwcq5fn
nU2GsNqN2OdFy9bDR2eUNWcr6Jn9iqwB8i82ihLIA4M2LBvpJJZeYHZBe0J7JgDB
IK1soaC4y3h0Ww2muoZC7rvezjIH7mcV69G4hTOFWNDt6pqoVNXFMlP8UxEDP8tW
/gJbtdNmo9cLhLRp0F9rydaZ2Kqo1PXZw4tTinq89g5R01Ujoh8WVVihWLkMDajT
irEcUtJbZY3Utuesp069uJA6CKzPeGfLo+iusuzPFd9qp4ccUF05SxPOT4ob5r/S
p4AkAUALZtkGrRfwQNkiLbEEiw0R9Bsx3/HU52DW+ikWViZjU53lLxdRZKGkDq/b
r3rNP7Im8XvU68fSZgHEE81Eu/Gh2qqFvS0dLRtBIo4YMRti4O2YBVwQDLhZ8Cfy
YBL3o8L8crmQtTcARKnBLHZimxb6ZEv6ejtp5wDEeIiMj2GbzZjuOxWLFwNwVnR0
sOlLCOeh/eJJuchcgFRB5FG+GzhP3HZSNgocDh+HC0PkwaFzZSnGKg+zohx9zPXP
P1NYwAR8ehTArf9HhTSEm13RLH3bLyXyky/PczfQWWglh8n1Fer4X48c0DJcAgjB
LTdYqtff5FBjhNMKHw24bto8YcoQsvhpnJJPPazYqJtnZdxW8K5Jb7sWgUwb3KiT
/7yOjc0OPLvTPlUD0o52b2BUOgPVwfF/956JMyKSiRMe0QRe25FdqMsj6x85dM6Y
QShW3z13GRCba9Gx8k6nc2ydBh3R2Wi8ZCHAH81zn1Z+EVsX9a6J4b9tkU9H8IKJ
wWnKO3ZgyZgU8X0ks67yug/++amY1ajN5IrgPcpyCJovRWwAkU35R5W9gUKMoXCW
3V9yY1xQMvhRf0HapHzwLlJsMyyOv2+jmIuGnjS4S2qajiuqyeBvQJq3obtSHJN1
ZiWRgK5dfS7Qlu02kVKsiB/JKqyCm8jrnIqESCyT7eO/TbUwEXkXQ1r3u/cYdZXJ
cUu7+j+XdS7rR9xX5r3nHbU4zo+iIgpSt7A8+4c2Kd+6leEwDiduDlqicoCCPCfs
EORb6sO8+J7XM3w2jTQWl8y/piu7YDSHxiJjtIOAP9yGnZ2Q3QCaf3qSIzHCnhOE
jKo2bwpRWetkGEj+YjN37C7qX8QfLGgQ3XbBJsmqHZMlbVeQXA0oqnKKZh9v1K5+
Jq72X9hvoScjaGkmlFksIcUl5DxpxZFi/croixDumoojGjl+6t2131EfyBpu1ryp
n1nJtLBlC+gWLWzYiT5QlqE2sB0XOeFMn8bzILrYOwOuDOygmYZrsBaJU79itz5C
qM+RINn2bJ/JooMSAMbjvrkMh1H/45J5+NK17gekesC5Yp1iz+++VI8y6tYiTKJL
lb61UOqCt8Zx9yknlEt/Ae7s4QVMH2rawGGMrKQDYoFlemwdjYicZO4pyOEe8znN
cE5acaQ7M/JUmeOP/e3MRPsLdIg8RNC3M78VmD5dfj50dD7xra1ghYCxmKL6o5wm
7r5RjlepHohnsHKaFezZRzLRhLZly8TW+vh8jja1W8XVOruZ0FHB7DtjGIDDRaK1
KzgTM+hdpn3q1+CRcZZYUTRObLPN8TVyua0uUk+u65oIvfZlLEZbe+au51TzYyQe
bseV9P9adgnQGdIALOZf4DtEhigbPCMhJbKeKj7g3t8Yz8hw1Vv6vGzduTnEN19F
+Oim3UEWA0nnJCdrbCINdTck3eWTs82vHU7jLHKI61P9kdHtp6609Sd+dEE/RXpS
U9kuOraZC5rdQgU1u/mNNW1uWREN+v7kIdGMTsYLLpdQK847Dj5rzNCm3s8N4Nrj
ZUr73hb3OdXyLhjWMRQ73XTRtahpCH8fHev72o2zvlJy2l5We4nbnoxWsdYIdWj1
X1/cACM4975Ljf+AcuoVg9zcmrOvQW0HOxWZrRVhx2/VavTpJMlVuFeJ3DRMtQYe
m0khomWoZEZjjZYVFYqTShRSLotaJZLkFFwAYlBFOhwZaFjbn8ap0mp1Nd3dQSBr
OZiQ/bxIYNXwMa7ce0EkWq0zl8t/jxA3oSBDHD0E556d/XjNIbuKKzTJDi0R4e3+
RPDxvDhWbzHzz+IX8ewVwBCOKulqBGBTbbN9ASBM14hFgBMABQHnJaNofzi99bNv
guyaZ+dTvZWQ3fTdYEJih8x3aTJKp3cfjgNVYfF2HIdZqKbH8UhIxYLVbMn/gliN
MuyTJCR5nEmG7UTQPE+XvYTzxoWSD4wBv8/B26dlPJ/Gt8Gl6Dc4XrZSioFEoY5E
LCI/pMJGGlN8WRL+1xP5qn7dc5AFJ5nCIYdYwhklJf5xz3WL54aiB8yZrEB0vadx
xALFtkWd2yxOLBaYGPuFORTpPP1SouxSXus/fER9SqmFDw7WrMDfZx2IDdvv742c
8Djqa5rjDCAnkfp//Y+UaVDI79Bt4p3WBCVLk1x7GFltOY4psKMeDYcETZ6GEvwJ
mu1o5zpfGZ9U6gPj1gv2pGWNfGgu8tM9vkaFAMWDwdPJoRM+LPkzZ4JdWu7Grb47
NzI1KWwqKD7I/0cB9bHyMWdQzStUY4VBjB1tObeP8m0fG83zPeIobCxkxuAv63Iy
LplRuztowgRr9mMXflzwzBqKD/joKYQk0AhUmbTncYUQQLFcl/II7DkgHLyFt3xX
uuki+WPleDWZYmgLT148uJsgHVYEATgxI6mt+96MjGwSSycyZnrBhp1MlxsYd2ed
gDFNevW8Ef45F1l36YWR28SAXQdVGR+umkbYQsd/Aq2VI13Quv5+2Pe1KWXQ9onc
n+jz0Ff7cpFpGudW0lbf4PrFc4GYOOQfaEdMC8TgSldXpEons+mpbQQ0bdsfb0Gs
D+toq9c+IXwmhX7ihEFRn23IEksMELN7txHMa9aglp6nj9g8LvjFNOnEEngbyzhT
7j+v1pO5xcBsJPz6fQptPiS4p3iVi4/OTSqDjc0V64P+GuCfdJ7Ujbtasu6S294E
cW8zNFJnLVHbp3u417PQzCteT7eskzfTpJLpDfcj2FjGl/YPfdLpSpxG1KGl4fQT
03XBUGL2qrUKEImY57Y+A6flZX9d2ZVqMUdXrNCsXdksSDtVKig0FEXUekIQ7lMU
wlh2yiC/njPrLpJz84Wo8yWpv32MQ4pjDfos7M5/xILiTOV7MRN94JyTeSTYJ1f0
iO5jPCgJhkoRAS8wSAJmT0VZ1G34t5wkm5qK2/IsSH4fOIVbdss4IaNLU/5pVDfS
eS6GqRLjhiQvHBD2PbQ4trcvAt1J6ixnboYHLq1V0M0lmX9m5N4DVy4Ktxjec0xE
UI1Seqp3+CO5rM2AKx1utXiXr5QuISsfJEVff5FlcRuTQmk/JhAcfiEzGi+8PEK3
+QI+tbYTs6Umn+/j6yc8+//rAugD1NJNsVSv88jFBg2qVh7bLMeW1tkd40+MfurF
VilB1NWjot45+CaF3zDpMquxG9OZARHHhG+X9TV6+KdFwaHYIc99lzumAvmxUeOo
wG3zgbgaGHBPI6JWnxL5b4HuMjLJfbgd5PaD7obeI1U6Bs1E233c1OdA9xHFrkSJ
/juJCkBnPX255bIzMYwNO661LTy4BURlj87acK8tlK9XbAbeo59y7gCDCcypqj71
Xq3ZjJqmr9yLPm0Q2lnOwH6fN4ZeNHQEJiEjEq+uigrY5DFOzqAh/0a9xQecma6P
COBljiXtsZK0FbTYGF/HxpMdLHB0eaO1MPics8dq7uT8SMJ+38HYt/CCSn4FeomP
dyyL0YSayY4XI+8bRMVDJWZzJb6UarJo/bD0xoskYfssvWAFeutSyaEOhVs8Nz4M
7+TxuEyTOTSiQO/XrsjBOWYuKaJI+t/8ZiV/dcJh9eBDF3g+66qMDMn4tQu86mHk
S3KNAti6QmxJEaUugBhOiB3/kSBrrD51K84GLVmEG3SRf8b717fwCPKsoIChOZyt
erUDhH/cwWjaMsDxbsScAmNeeQjOB0t0qCCX2/4prEq/uNA0SjJ/EPJvoGr+h3nB
NqiCyZ2WaRAKctiRxKHeCvnXh8T8JOWqX/l+d/Q+X7M7NyQFSVlZr2nSZ6apr67Q
17ofEovjomQ0xHfi1bDLhJ9fjqzHYg6pKFD0PsV84s+TXf51OlcVza9s0wX4Nm4P
/7Zo3WK/W7qxk+eU3o5MTTnx7GOVobLSUKI4QLGsWfohSpR9ZpT7WrxwRnSUiiAB
cNhCEZMuK1BaXDdAjc4K6yurwYh1poCPh4y7I7dzI/SD5EPvg27Vc9j8PDEEcRej
DtT6GnR8YLVAfuVKyeA03PqiZDeXO8A6BSqgcP0BvI0aPv9fw1k40Gl10PEIWaht
gOk8HBJSWkyd4m9PmIbBDXL3C1o1m6r0uHialrBdpAIf+Ey1hUq8/gYSdEzp4r2K
3h9+Hk/sNukjiRZnXoe66UXH8DGtaLyHzUb3oQgGL8jCj80iIZ022EPJ5IVvposE
R/teiw4dCG7o56f64d9s662P/IXdcOEWw1k1ALNrGtxdErwVGLIm8oMiYQYnNiJi
yVKYdELYokOInU+WVR6e3wT9xJEreRjaEPes9+cqhG+M07c7WfU0civX3SqEdNtE
8TgJbSUOPsvq9nhS3w5VvnnUW/9el6YIkqKmpwmy8KirKfrAfPvLYNgA1ek+3iTb
FcU39SC0wUfyxvs15/z+zbn36u4TtOZL+V65dBgplXJbCwx03u9KZ48MRCdL6OZC
jmRTbkY1AUQwfWmT55sMEZFbbzdOOdwyRbdT+3Bf/yf3k4PkP4Uh7g9lY/S8sjiA
o/QxaZGXrwMuPsmqzYaxDWUfbHCfaHQjE4ulSp6IHFar+D3fk6AmMnb8XqCu5JEu
ChPYYjDdcjwmC4u9MgKvAca91Pv+XL9TRXhpLXWsl38/JrDJh9C91pI/sC/5QfN6
pP89BRt3lPuSHDGWpGuNdqlwWZTayjFNBBZJ+cbxT+iKcwsz8DGKUOwiwtnCrgu9
JWVI0InhCjvTuzWhce9yhmk+7S0BhuxIVauPNtLm3KAwdTT6LmRJkgb/wwQNgCq5
C9cQWIkJt6Neix2yZ4jLcDxajPgTV5B5iwL+Ji56mwJ40UloQBDEYNjXY9iuCpxc
aG3ELc8X5i2rMxMyoy53RiwrWitJ878cTWKXTtDio2JWyU0mxxMw0XUXEFzbHkdG
DBDeFBOXJetzvYIeNuG8M7JgSSeBkpTzZDe2FakoPlut9wPzvzC71ci9n/Or7CzX
CDZsRZMiDciKshoecetMyO5WrHpUG3khdGEOJVMSDLRd64PrOjd4JDYGWuXQ3mim
cfEklRVrPusji6ZnX4t8zUH06uJjj5m5DdXL8eShCeH4hHnZZo71uPyIiUskKX+m
Ov5G5UXW8S6kVoSmJBRbEsRYHnlmB1xk/7mVgxGRb5ZBcSrWbCpXqMzZueXOsTR6
5MSozg2tljnMK2FeulluXl/khST1P7LYG1hv7OwiQryYcERThzoy/jzbPRmxR/h6
b2QPc/aY2pJgW+IVDzsQG083NYtKgUYJl1NZVCBVLqUPfuFZvZtftQ/Nb58GN+R8
NOf8Omj4DswlV2wMs3Yx2i/KffYwx07XgNu1ZV2H2Gc0UkgskZ4vE4fmYJAW9KU1
rydQLTbwBaoXqCWVWY8rJ+2D8Sa7j2dWvYB2wibtZj8E5jZl1MafbckD09qVTv53
qhSw38xjpTLZ23YapA16GspOYKU/teaJ7QPdatugJvzycFxjl4IsRpYLaH2f9Mb9
cbKYCQ+R20fGr8S6S4A0E3Z9KDKSeDAFjzS6oL0S08Gn0GgdsF8Ssx7MwhWmZibk
HaIUM1H9iWrbxe6dbH24tdUqb9YnPdLU2vA2Lg7jqPe5sgFt4YI06SsAhMboydON
FAhviCS4zNifREv5fruQHzNrIwMEQme3KwmhPoXTMGRuxedL1veQ7GuNMrPwY3fv
IktX+cjIThHOfSYweyLpdfaz4uHT+velNg+WwpJGk8V4Vo4Ki1yRvI6v53OZrHj4
9JDfY527eIcuwygF6NVyvDbR9PAw9H9rVJxmyd40YBYidM7womu0UMNC/LvDfqc7
03RKBUlFfLRDjevTzbnQcgV3/NmTwYKGwMUG5KvwxLFpP8Is0VqY6NXAgSWglARe
VktjxV6mdftvi8reYxvZ6rnLwjTA3sQYXh8GqY347ysn2XSe77umwFEGF8iA1BFA
3SsTz7LxZoo308PzJ462GgBUjrotdyuEqOj2pag3xk0B68JEqdCVMhrDEd3PjXWg
1jVG27+UpbzYghZmxA510QFLVm8qIMwCgJBdCUTbuQbcSTSkzCmCWQwJgimkIoRd
LASJgXNQeFugSZSczuEEX6GCa8K7kLpEax+JGKyDLsnf1rqklLFgUzfvS+iA4GcQ
WwAKVm4tAmoPO5y3O19eoE/fKOJKiP6zzeWBS0s4nnTG1zdjvoX2Wj+jJkCfAoER
A8Jr74DdIy80fNr2+ZRgkDcYwg7DWP5lV82tv1C3LowHpaeKonkcshrqCopE/QMu
upxAGuCQzywGq5/V5nnHb8yC3mbe4JqBzecsArXNj8c6m86OVBFh0vJz627gm+Nx
3IVIZg/zW3OzqbBM0sk2qzLdXgoik3TDVEBKokC35C4GiBkXC/nXflDtXF86bFDo
/D0XMKTPAGBl3v7uKvZwOzd3M3rdoTkbEwgmwOVjkXp2tiGTzHKE00e4MzEllEDA
m89wcUUY/W/2+aQeRREblrvh+Haf6DMZj8lsIjNjX6srdx59FyhOpZQuSRHDYDfx
Cp7w2tP7jM9p9kXwjFBOA2/OBWYTIZ8tu0fAbknEaUvmetL3Ri5+Pvi+StssetDL
OBK8ZslWB6IeFnVDki/SetLzdgjkt4MqnsRJeo/tCZrAHNpZ7Vc3+NoRVAQ7OFvj
cwwP0UqcL9ix6761+gJ/9aFEkYVF16w3Y+Zi2nuQ7ebCzrKbuPcSuJxumx7s9Q/v
JunT7DdY8I27c3P9G6qVvwedkRNC+b2Xc+pU77OIP6swziB6eawOXwCNcyWclAFY
P05XV3FPB8V7VxZgAfGyD0O6BczcZKgGBfXYwlpt91WsQtUMRwhrs0/lC6kaXAKv
vhhSX1MQYFRnuGj15nf1wYA76SuNETT7UlernPxQi/YAbIlsQheoV20P56PpYpfO
aSSZaiVn23whNkggbn+EvAmpgPHTpXg//PHTngh3HYC1yc/L0f382q5OWrXHdIro
6oMJZ9KZmtWwLJeelnAxpfthixthKN3Ddvz56toNO3ZrQYI6sznqIFQRQmmlNaYf
h2bsDscD4rnP1U/r6f+25ayV8RjILbCfyN2H/uwbgDUim0gTUVFUvr0vmzUKw2bJ
MpTEYUiQ7RULqbNde+eACNHRhxdnLek12mzULWrczjQKf/wDJwfS3FpL5unR1H7V
lQYoKU7oSBL+I7ELNauh2zv2i114Fj1O3ZodTSYL/yxs/fYRoh7TY2JW2CWNF04b
OFs1tIcUE+X9NZqPhklfNZJ+HALcca6KFbDayMz9R5UC1U1QfWT+kkEw3BvuY5b2
ypxuorSJuRNKpXbCfXU4l3BtYoTWpbYpossV4+LFPMwDsal0BMdLXweFmpSJ1jkC
/roCd0BNKSoRErKyx+Q3UP4pNzE3768LOBqrb9zQIxtjSEclcFsHByZD2t+ZXOyH
JDpXt7WgZ6Qm8uQ0GTZ+oHyahF/eSz6YiOOOZ0WArGSDt78duZX+97qMA0YU1TRO
oWsuin4f/wU/LztlaJrpH2qmVjFC0tJPJfzuDd9Mrb2ADkDT/U8gil6Wk7Dv5dGS
cM8J3ajA5uJwuFEnfurvhV5Fs+2lrzVCOSvjEwOTULrjfQ6Qkx2aJPYgJ54eA76W
WLh3of6iw8ALbB1U6xVV7I8tcClbqbhgJdwt4zBCdxiP9nZ8062SK1cPPkmq12Js
x5AxEFy284Aa2SW3IDKfDmSp0YYRhhMFCPmfFCEg0MufyingI8ZJ1wfYW+4yWLya
w08ONkSx0ffGFMRd3O2WHhd7YTuY3jyxK5mQr1vfcZQXNbYL2K+BdeOZ+fAaggwY
CW8ORf5SnfwvX8VzpVDNNu9rj0bfdBOXaLLFqI28jjEkmdhG53j0GQWwmTWHvlhO
AJ/dWCqVK1Ih2m+OuA1H55KWAPbCfGJKxuxW690dNFOOPzV93FNCS278wXLegtTB
UrfbxwBWvGvuTzfz2Y3MFXTIFNWwoPQm2sk6+8H2LBiOwBXeS28D0r5jHiG/5CqJ
2MGZr0J7zG60VieTXdnJTZKn9+IpCMttuIMeWTnymAyafuQcn/F5i4+ffT8EMumD
7wnQHMUZTGzFr7M24l/C39qRC9gZUH+zwta9DNfUbIr0SZ4Yt+XVRlp0TcIthb6s
80Rd2kZgOqH5IW6Opz+/fv9lkaKxyAaVIqH5F69tPSPzWUf24PxczInpNIgI8mBX
X1HcirnqVlQeivGge7xkl3NvJsd5siJMZHnmFqkUnoPjWh2ahhX1mldCcb3SlUnx
5ERwqQ+aDSLMMxw5I5CwBrcgznciQ8EJxN5iNKyXh3EtpptZRlzQZKR9KHiqDh5+
3nz4WTvnTnqsnsdYFsg7F8++24dTV7ZZg9Vh0xduK3LcZWuoVbyEDbq0hKuPsVyh
v5bd/FPsB119TXugxAGnq37b8RM8v2S5o3yaHnn5Zw/ExuEw4k9kJdaTK3wHBLSh
Dv4HSX3rrxvhe0IeF7W4Mlbfdj5yNNMtJlf7+BpTqt3aAxKveKxWTqFg0mjIAfIl
XfYraQkNnmtDi0Os8eGydxsUZJLkIfxFBcLbUWXH7MEyKaxf2pVbOecIvKOAndm5
/A7BPiZzs4uHz8BhO5D8J9uugk9LT+z22pHBA7ot1zq9hNmpHt0ZYxF69jZMiJ0U
9TGJ3TAqzjJSa3f9ERb3scYrGWGuYWh7PpmRyFYpiTvuI6awhS2fQ7HlCBb3r3KW
zfs0ujG49yza3uxTdPw96MazJ64+5ZsV4inUcNDvueZkTFnAK3hT6Gbf/U4AZ4tV
JvuF3sVgB2NF79nmMq7cvIxMtGaqXoKjH9vVvwZVuWA+QIIO6f768vrQsGqm63y5
9YZ46beBHvK9DYMmeXGrTTW0BMQJ0Ocz7FF6tWuxwg8M2LSkVRjqDBEesiwgEgdY
8GWhUjUJRE477syCZI0b/W+DSvDh32VkSrwB/tPmnkT4RhCOxU0XxeRZGR2+1vC8
sF8tzJSzTbt1Wa9tvE5wu7NpAu//mPKJaAXUsh2S/io5QS55irf6Z8nLOiXkTIsK
u3YIK231OtwsHMotjO0h7l6VdQHehO0mgQG6KvG9w171FfnZqSE8GNB8vAIAvaxG
E29/m0WcDUWa+/+4cEyhdY4oz4oR//c643k64BiFQQsulV60ueqhbG3ycKEsXySi
7XGsC5esbBn2dBiZrIyItXtkdgo2oJnZ1MoVAjlEZEyuNaYRNrB0/wuG5nwPbnvO
J++eumnYnncWGZ6Ele1EYZ4k74Iagt7H5y5wkfNqkjnP+RWr+ZWfhfhWla12qY3G
JVhRxrAGXqcer/uoiw62wpK+JEh5gCtRyC25KCgLnitMj7aryECxrHgmLQMl6Qao
8MYyuIJj7a5749TgkfgIXXjbYoIVB0QLmAFYbiZbqLtXjL3TNyDAYLy0M7xWDu7x
/e9nrOyHI0WpN2bJHfjG6/CAsPZXMk4ZNy1QWUfzrrbEuQH1UNN5XFTXgApjEMNv
tfuhmwJkusM2NgRi+VToXpJHXHgsjm4OKLLwiGLd/qhLt8uhPRSq0Ui4quvHgd24
r6RfXHdQ4tdXIXGpMori99ElB/gdjMXgNRLonHNGhASk50kmnKFxRKAYqJk8bzPn
i9n/GtYoLoyxj1mBFPqQbA==
`pragma protect end_protected
