// top.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module top (
		input  wire        clk_clk,                                                 //                                     clk.clk
		input  wire [2:0]  ddr3a_status_external_connection_export,                 //        ddr3a_status_external_connection.export
		input  wire [2:0]  ddr3b_status_external_connection_export,                 //        ddr3b_status_external_connection.export
		input  wire [31:0] hip_ctrl_test_in,                                        //                                hip_ctrl.test_in
		input  wire        hip_ctrl_simu_mode_pipe,                                 //                                        .simu_mode_pipe
		input  wire        hip_pipe_sim_pipe_pclk_in,                               //                                hip_pipe.sim_pipe_pclk_in
		output wire [1:0]  hip_pipe_sim_pipe_rate,                                  //                                        .sim_pipe_rate
		output wire [4:0]  hip_pipe_sim_ltssmstate,                                 //                                        .sim_ltssmstate
		output wire [2:0]  hip_pipe_eidleinfersel0,                                 //                                        .eidleinfersel0
		output wire [2:0]  hip_pipe_eidleinfersel1,                                 //                                        .eidleinfersel1
		output wire [2:0]  hip_pipe_eidleinfersel2,                                 //                                        .eidleinfersel2
		output wire [2:0]  hip_pipe_eidleinfersel3,                                 //                                        .eidleinfersel3
		output wire [2:0]  hip_pipe_eidleinfersel4,                                 //                                        .eidleinfersel4
		output wire [2:0]  hip_pipe_eidleinfersel5,                                 //                                        .eidleinfersel5
		output wire [2:0]  hip_pipe_eidleinfersel6,                                 //                                        .eidleinfersel6
		output wire [2:0]  hip_pipe_eidleinfersel7,                                 //                                        .eidleinfersel7
		output wire [1:0]  hip_pipe_powerdown0,                                     //                                        .powerdown0
		output wire [1:0]  hip_pipe_powerdown1,                                     //                                        .powerdown1
		output wire [1:0]  hip_pipe_powerdown2,                                     //                                        .powerdown2
		output wire [1:0]  hip_pipe_powerdown3,                                     //                                        .powerdown3
		output wire [1:0]  hip_pipe_powerdown4,                                     //                                        .powerdown4
		output wire [1:0]  hip_pipe_powerdown5,                                     //                                        .powerdown5
		output wire [1:0]  hip_pipe_powerdown6,                                     //                                        .powerdown6
		output wire [1:0]  hip_pipe_powerdown7,                                     //                                        .powerdown7
		output wire        hip_pipe_rxpolarity0,                                    //                                        .rxpolarity0
		output wire        hip_pipe_rxpolarity1,                                    //                                        .rxpolarity1
		output wire        hip_pipe_rxpolarity2,                                    //                                        .rxpolarity2
		output wire        hip_pipe_rxpolarity3,                                    //                                        .rxpolarity3
		output wire        hip_pipe_rxpolarity4,                                    //                                        .rxpolarity4
		output wire        hip_pipe_rxpolarity5,                                    //                                        .rxpolarity5
		output wire        hip_pipe_rxpolarity6,                                    //                                        .rxpolarity6
		output wire        hip_pipe_rxpolarity7,                                    //                                        .rxpolarity7
		output wire        hip_pipe_txcompl0,                                       //                                        .txcompl0
		output wire        hip_pipe_txcompl1,                                       //                                        .txcompl1
		output wire        hip_pipe_txcompl2,                                       //                                        .txcompl2
		output wire        hip_pipe_txcompl3,                                       //                                        .txcompl3
		output wire        hip_pipe_txcompl4,                                       //                                        .txcompl4
		output wire        hip_pipe_txcompl5,                                       //                                        .txcompl5
		output wire        hip_pipe_txcompl6,                                       //                                        .txcompl6
		output wire        hip_pipe_txcompl7,                                       //                                        .txcompl7
		output wire [7:0]  hip_pipe_txdata0,                                        //                                        .txdata0
		output wire [7:0]  hip_pipe_txdata1,                                        //                                        .txdata1
		output wire [7:0]  hip_pipe_txdata2,                                        //                                        .txdata2
		output wire [7:0]  hip_pipe_txdata3,                                        //                                        .txdata3
		output wire [7:0]  hip_pipe_txdata4,                                        //                                        .txdata4
		output wire [7:0]  hip_pipe_txdata5,                                        //                                        .txdata5
		output wire [7:0]  hip_pipe_txdata6,                                        //                                        .txdata6
		output wire [7:0]  hip_pipe_txdata7,                                        //                                        .txdata7
		output wire        hip_pipe_txdatak0,                                       //                                        .txdatak0
		output wire        hip_pipe_txdatak1,                                       //                                        .txdatak1
		output wire        hip_pipe_txdatak2,                                       //                                        .txdatak2
		output wire        hip_pipe_txdatak3,                                       //                                        .txdatak3
		output wire        hip_pipe_txdatak4,                                       //                                        .txdatak4
		output wire        hip_pipe_txdatak5,                                       //                                        .txdatak5
		output wire        hip_pipe_txdatak6,                                       //                                        .txdatak6
		output wire        hip_pipe_txdatak7,                                       //                                        .txdatak7
		output wire        hip_pipe_txdetectrx0,                                    //                                        .txdetectrx0
		output wire        hip_pipe_txdetectrx1,                                    //                                        .txdetectrx1
		output wire        hip_pipe_txdetectrx2,                                    //                                        .txdetectrx2
		output wire        hip_pipe_txdetectrx3,                                    //                                        .txdetectrx3
		output wire        hip_pipe_txdetectrx4,                                    //                                        .txdetectrx4
		output wire        hip_pipe_txdetectrx5,                                    //                                        .txdetectrx5
		output wire        hip_pipe_txdetectrx6,                                    //                                        .txdetectrx6
		output wire        hip_pipe_txdetectrx7,                                    //                                        .txdetectrx7
		output wire        hip_pipe_txelecidle0,                                    //                                        .txelecidle0
		output wire        hip_pipe_txelecidle1,                                    //                                        .txelecidle1
		output wire        hip_pipe_txelecidle2,                                    //                                        .txelecidle2
		output wire        hip_pipe_txelecidle3,                                    //                                        .txelecidle3
		output wire        hip_pipe_txelecidle4,                                    //                                        .txelecidle4
		output wire        hip_pipe_txelecidle5,                                    //                                        .txelecidle5
		output wire        hip_pipe_txelecidle6,                                    //                                        .txelecidle6
		output wire        hip_pipe_txelecidle7,                                    //                                        .txelecidle7
		output wire        hip_pipe_txdeemph0,                                      //                                        .txdeemph0
		output wire        hip_pipe_txdeemph1,                                      //                                        .txdeemph1
		output wire        hip_pipe_txdeemph2,                                      //                                        .txdeemph2
		output wire        hip_pipe_txdeemph3,                                      //                                        .txdeemph3
		output wire        hip_pipe_txdeemph4,                                      //                                        .txdeemph4
		output wire        hip_pipe_txdeemph5,                                      //                                        .txdeemph5
		output wire        hip_pipe_txdeemph6,                                      //                                        .txdeemph6
		output wire        hip_pipe_txdeemph7,                                      //                                        .txdeemph7
		output wire [2:0]  hip_pipe_txmargin0,                                      //                                        .txmargin0
		output wire [2:0]  hip_pipe_txmargin1,                                      //                                        .txmargin1
		output wire [2:0]  hip_pipe_txmargin2,                                      //                                        .txmargin2
		output wire [2:0]  hip_pipe_txmargin3,                                      //                                        .txmargin3
		output wire [2:0]  hip_pipe_txmargin4,                                      //                                        .txmargin4
		output wire [2:0]  hip_pipe_txmargin5,                                      //                                        .txmargin5
		output wire [2:0]  hip_pipe_txmargin6,                                      //                                        .txmargin6
		output wire [2:0]  hip_pipe_txmargin7,                                      //                                        .txmargin7
		output wire        hip_pipe_txswing0,                                       //                                        .txswing0
		output wire        hip_pipe_txswing1,                                       //                                        .txswing1
		output wire        hip_pipe_txswing2,                                       //                                        .txswing2
		output wire        hip_pipe_txswing3,                                       //                                        .txswing3
		output wire        hip_pipe_txswing4,                                       //                                        .txswing4
		output wire        hip_pipe_txswing5,                                       //                                        .txswing5
		output wire        hip_pipe_txswing6,                                       //                                        .txswing6
		output wire        hip_pipe_txswing7,                                       //                                        .txswing7
		input  wire        hip_pipe_phystatus0,                                     //                                        .phystatus0
		input  wire        hip_pipe_phystatus1,                                     //                                        .phystatus1
		input  wire        hip_pipe_phystatus2,                                     //                                        .phystatus2
		input  wire        hip_pipe_phystatus3,                                     //                                        .phystatus3
		input  wire        hip_pipe_phystatus4,                                     //                                        .phystatus4
		input  wire        hip_pipe_phystatus5,                                     //                                        .phystatus5
		input  wire        hip_pipe_phystatus6,                                     //                                        .phystatus6
		input  wire        hip_pipe_phystatus7,                                     //                                        .phystatus7
		input  wire [7:0]  hip_pipe_rxdata0,                                        //                                        .rxdata0
		input  wire [7:0]  hip_pipe_rxdata1,                                        //                                        .rxdata1
		input  wire [7:0]  hip_pipe_rxdata2,                                        //                                        .rxdata2
		input  wire [7:0]  hip_pipe_rxdata3,                                        //                                        .rxdata3
		input  wire [7:0]  hip_pipe_rxdata4,                                        //                                        .rxdata4
		input  wire [7:0]  hip_pipe_rxdata5,                                        //                                        .rxdata5
		input  wire [7:0]  hip_pipe_rxdata6,                                        //                                        .rxdata6
		input  wire [7:0]  hip_pipe_rxdata7,                                        //                                        .rxdata7
		input  wire        hip_pipe_rxdatak0,                                       //                                        .rxdatak0
		input  wire        hip_pipe_rxdatak1,                                       //                                        .rxdatak1
		input  wire        hip_pipe_rxdatak2,                                       //                                        .rxdatak2
		input  wire        hip_pipe_rxdatak3,                                       //                                        .rxdatak3
		input  wire        hip_pipe_rxdatak4,                                       //                                        .rxdatak4
		input  wire        hip_pipe_rxdatak5,                                       //                                        .rxdatak5
		input  wire        hip_pipe_rxdatak6,                                       //                                        .rxdatak6
		input  wire        hip_pipe_rxdatak7,                                       //                                        .rxdatak7
		input  wire        hip_pipe_rxelecidle0,                                    //                                        .rxelecidle0
		input  wire        hip_pipe_rxelecidle1,                                    //                                        .rxelecidle1
		input  wire        hip_pipe_rxelecidle2,                                    //                                        .rxelecidle2
		input  wire        hip_pipe_rxelecidle3,                                    //                                        .rxelecidle3
		input  wire        hip_pipe_rxelecidle4,                                    //                                        .rxelecidle4
		input  wire        hip_pipe_rxelecidle5,                                    //                                        .rxelecidle5
		input  wire        hip_pipe_rxelecidle6,                                    //                                        .rxelecidle6
		input  wire        hip_pipe_rxelecidle7,                                    //                                        .rxelecidle7
		input  wire [2:0]  hip_pipe_rxstatus0,                                      //                                        .rxstatus0
		input  wire [2:0]  hip_pipe_rxstatus1,                                      //                                        .rxstatus1
		input  wire [2:0]  hip_pipe_rxstatus2,                                      //                                        .rxstatus2
		input  wire [2:0]  hip_pipe_rxstatus3,                                      //                                        .rxstatus3
		input  wire [2:0]  hip_pipe_rxstatus4,                                      //                                        .rxstatus4
		input  wire [2:0]  hip_pipe_rxstatus5,                                      //                                        .rxstatus5
		input  wire [2:0]  hip_pipe_rxstatus6,                                      //                                        .rxstatus6
		input  wire [2:0]  hip_pipe_rxstatus7,                                      //                                        .rxstatus7
		input  wire        hip_pipe_rxvalid0,                                       //                                        .rxvalid0
		input  wire        hip_pipe_rxvalid1,                                       //                                        .rxvalid1
		input  wire        hip_pipe_rxvalid2,                                       //                                        .rxvalid2
		input  wire        hip_pipe_rxvalid3,                                       //                                        .rxvalid3
		input  wire        hip_pipe_rxvalid4,                                       //                                        .rxvalid4
		input  wire        hip_pipe_rxvalid5,                                       //                                        .rxvalid5
		input  wire        hip_pipe_rxvalid6,                                       //                                        .rxvalid6
		input  wire        hip_pipe_rxvalid7,                                       //                                        .rxvalid7
		input  wire        hip_serial_rx_in0,                                       //                              hip_serial.rx_in0
		input  wire        hip_serial_rx_in1,                                       //                                        .rx_in1
		input  wire        hip_serial_rx_in2,                                       //                                        .rx_in2
		input  wire        hip_serial_rx_in3,                                       //                                        .rx_in3
		input  wire        hip_serial_rx_in4,                                       //                                        .rx_in4
		input  wire        hip_serial_rx_in5,                                       //                                        .rx_in5
		input  wire        hip_serial_rx_in6,                                       //                                        .rx_in6
		input  wire        hip_serial_rx_in7,                                       //                                        .rx_in7
		output wire        hip_serial_tx_out0,                                      //                                        .tx_out0
		output wire        hip_serial_tx_out1,                                      //                                        .tx_out1
		output wire        hip_serial_tx_out2,                                      //                                        .tx_out2
		output wire        hip_serial_tx_out3,                                      //                                        .tx_out3
		output wire        hip_serial_tx_out4,                                      //                                        .tx_out4
		output wire        hip_serial_tx_out5,                                      //                                        .tx_out5
		output wire        hip_serial_tx_out6,                                      //                                        .tx_out6
		output wire        hip_serial_tx_out7,                                      //                                        .tx_out7
		output wire [14:0] mem_if_ddr3a_mem_mem_a,                                  //                        mem_if_ddr3a_mem.mem_a
		output wire [2:0]  mem_if_ddr3a_mem_mem_ba,                                 //                                        .mem_ba
		output wire [0:0]  mem_if_ddr3a_mem_mem_ck,                                 //                                        .mem_ck
		output wire [0:0]  mem_if_ddr3a_mem_mem_ck_n,                               //                                        .mem_ck_n
		output wire [0:0]  mem_if_ddr3a_mem_mem_cke,                                //                                        .mem_cke
		output wire [0:0]  mem_if_ddr3a_mem_mem_cs_n,                               //                                        .mem_cs_n
		output wire [7:0]  mem_if_ddr3a_mem_mem_dm,                                 //                                        .mem_dm
		output wire [0:0]  mem_if_ddr3a_mem_mem_ras_n,                              //                                        .mem_ras_n
		output wire [0:0]  mem_if_ddr3a_mem_mem_cas_n,                              //                                        .mem_cas_n
		output wire [0:0]  mem_if_ddr3a_mem_mem_we_n,                               //                                        .mem_we_n
		output wire        mem_if_ddr3a_mem_mem_reset_n,                            //                                        .mem_reset_n
		inout  wire [63:0] mem_if_ddr3a_mem_mem_dq,                                 //                                        .mem_dq
		inout  wire [7:0]  mem_if_ddr3a_mem_mem_dqs,                                //                                        .mem_dqs
		inout  wire [7:0]  mem_if_ddr3a_mem_mem_dqs_n,                              //                                        .mem_dqs_n
		output wire [0:0]  mem_if_ddr3a_mem_mem_odt,                                //                                        .mem_odt
		input  wire        mem_if_ddr3a_oct_rzqin,                                  //                        mem_if_ddr3a_oct.rzqin
		input  wire        mem_if_ddr3a_pll_ref_clk_clk,                            //                mem_if_ddr3a_pll_ref_clk.clk
		output wire        mem_if_ddr3a_status_local_init_done,                     //                     mem_if_ddr3a_status.local_init_done
		output wire        mem_if_ddr3a_status_local_cal_success,                   //                                        .local_cal_success
		output wire        mem_if_ddr3a_status_local_cal_fail,                      //                                        .local_cal_fail
		output wire [14:0] mem_if_ddr3b_mem_mem_a,                                  //                        mem_if_ddr3b_mem.mem_a
		output wire [2:0]  mem_if_ddr3b_mem_mem_ba,                                 //                                        .mem_ba
		output wire [0:0]  mem_if_ddr3b_mem_mem_ck,                                 //                                        .mem_ck
		output wire [0:0]  mem_if_ddr3b_mem_mem_ck_n,                               //                                        .mem_ck_n
		output wire [0:0]  mem_if_ddr3b_mem_mem_cke,                                //                                        .mem_cke
		output wire [0:0]  mem_if_ddr3b_mem_mem_cs_n,                               //                                        .mem_cs_n
		output wire [7:0]  mem_if_ddr3b_mem_mem_dm,                                 //                                        .mem_dm
		output wire [0:0]  mem_if_ddr3b_mem_mem_ras_n,                              //                                        .mem_ras_n
		output wire [0:0]  mem_if_ddr3b_mem_mem_cas_n,                              //                                        .mem_cas_n
		output wire [0:0]  mem_if_ddr3b_mem_mem_we_n,                               //                                        .mem_we_n
		output wire        mem_if_ddr3b_mem_mem_reset_n,                            //                                        .mem_reset_n
		inout  wire [63:0] mem_if_ddr3b_mem_mem_dq,                                 //                                        .mem_dq
		inout  wire [7:0]  mem_if_ddr3b_mem_mem_dqs,                                //                                        .mem_dqs
		inout  wire [7:0]  mem_if_ddr3b_mem_mem_dqs_n,                              //                                        .mem_dqs_n
		output wire [0:0]  mem_if_ddr3b_mem_mem_odt,                                //                                        .mem_odt
		input  wire        mem_if_ddr3b_oct_rzqin,                                  //                        mem_if_ddr3b_oct.rzqin
		input  wire        mem_if_ddr3b_pll_ref_clk_clk,                            //                mem_if_ddr3b_pll_ref_clk.clk
		output wire        mem_if_ddr3b_status_local_init_done,                     //                     mem_if_ddr3b_status.local_init_done
		output wire        mem_if_ddr3b_status_local_cal_success,                   //                                        .local_cal_success
		output wire        mem_if_ddr3b_status_local_cal_fail,                      //                                        .local_cal_fail
		output wire        pcie_256_hip_avmm_0_reconfig_clk_locked_fixedclk_locked, // pcie_256_hip_avmm_0_reconfig_clk_locked.fixedclk_locked
		input  wire        pcie_rstn_npor,                                          //                               pcie_rstn.npor
		input  wire        pcie_rstn_pin_perst,                                     //                                        .pin_perst
		input  wire [3:0]  pio_button_external_connection_export,                   //          pio_button_external_connection.export
		output wire [3:0]  pio_led_external_connection_export,                      //             pio_led_external_connection.export
		input  wire        refclk_clk,                                              //                                  refclk.clk
		input  wire        reset_reset_n                                            //                                   reset.reset_n
	);

	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_readdata;                     // alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> pcie_reconfig_driver_0:reconfig_mgmt_readdata
	wire          pcie_reconfig_driver_0_reconfig_mgmt_waitrequest;                  // alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> pcie_reconfig_driver_0:reconfig_mgmt_waitrequest
	wire    [6:0] pcie_reconfig_driver_0_reconfig_mgmt_address;                      // pcie_reconfig_driver_0:reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	wire          pcie_reconfig_driver_0_reconfig_mgmt_read;                         // pcie_reconfig_driver_0:reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	wire          pcie_reconfig_driver_0_reconfig_mgmt_write;                        // pcie_reconfig_driver_0:reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_writedata;                    // pcie_reconfig_driver_0:reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	wire          mem_if_ddr3a_afi_clk_clk;                                          // mem_if_ddr3a:afi_clk -> [mm_clock_crossing_bridge_ddr3a:m0_clk, mm_interconnect_1:mem_if_ddr3a_afi_clk_clk, rst_controller_002:clk]
	wire          mem_if_ddr3b_afi_clk_clk;                                          // mem_if_ddr3b:afi_clk -> [mm_clock_crossing_bridge_ddr3b:m0_clk, mm_interconnect_2:mem_if_ddr3b_afi_clk_clk, rst_controller_004:clk]
	wire          pcie_256_dma_coreclkout_clk;                                       // pcie_256_dma:coreclkout -> [mm_clock_crossing_bridge_ddr3a:s0_clk, mm_clock_crossing_bridge_ddr3b:s0_clk, mm_interconnect_0:pcie_256_dma_coreclkout_clk, mm_interconnect_3:pcie_256_dma_coreclkout_clk, onchip_memory2_0:clk, onchip_memory2_0:clk2, pcie_reconfig_driver_0:pld_clk, pio_button:clk, pio_led:clk, rst_controller_003:clk, rst_controller_005:clk]
	wire    [1:0] pcie_256_dma_hip_currentspeed_currentspeed;                        // pcie_256_dma:currentspeed -> pcie_reconfig_driver_0:currentspeed
	wire          alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy;                   // alt_xcvr_reconfig_0:reconfig_busy -> pcie_reconfig_driver_0:reconfig_busy
	wire  [505:0] pcie_256_dma_reconfig_from_xcvr_reconfig_from_xcvr;                // pcie_256_dma:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire  [769:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr;             // alt_xcvr_reconfig_0:reconfig_to_xcvr -> pcie_256_dma:reconfig_to_xcvr
	wire          pcie_256_dma_rxm_bar4_waitrequest;                                 // mm_interconnect_0:pcie_256_dma_Rxm_BAR4_waitrequest -> pcie_256_dma:RxmWaitRequest_4_i
	wire   [31:0] pcie_256_dma_rxm_bar4_readdata;                                    // mm_interconnect_0:pcie_256_dma_Rxm_BAR4_readdata -> pcie_256_dma:RxmReadData_4_i
	wire   [63:0] pcie_256_dma_rxm_bar4_address;                                     // pcie_256_dma:RxmAddress_4_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR4_address
	wire          pcie_256_dma_rxm_bar4_read;                                        // pcie_256_dma:RxmRead_4_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR4_read
	wire    [3:0] pcie_256_dma_rxm_bar4_byteenable;                                  // pcie_256_dma:RxmByteEnable_4_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR4_byteenable
	wire          pcie_256_dma_rxm_bar4_readdatavalid;                               // mm_interconnect_0:pcie_256_dma_Rxm_BAR4_readdatavalid -> pcie_256_dma:RxmReadDataValid_4_i
	wire          pcie_256_dma_rxm_bar4_write;                                       // pcie_256_dma:RxmWrite_4_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR4_write
	wire   [31:0] pcie_256_dma_rxm_bar4_writedata;                                   // pcie_256_dma:RxmWriteData_4_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR4_writedata
	wire          pcie_256_dma_dma_rd_master_waitrequest;                            // mm_interconnect_0:pcie_256_dma_dma_rd_master_waitrequest -> pcie_256_dma:RdDmaWaitRequest_i
	wire   [63:0] pcie_256_dma_dma_rd_master_address;                                // pcie_256_dma:RdDmaAddress_o -> mm_interconnect_0:pcie_256_dma_dma_rd_master_address
	wire   [31:0] pcie_256_dma_dma_rd_master_byteenable;                             // pcie_256_dma:RdDmaWriteEnable_o -> mm_interconnect_0:pcie_256_dma_dma_rd_master_byteenable
	wire          pcie_256_dma_dma_rd_master_write;                                  // pcie_256_dma:RdDmaWrite_o -> mm_interconnect_0:pcie_256_dma_dma_rd_master_write
	wire  [255:0] pcie_256_dma_dma_rd_master_writedata;                              // pcie_256_dma:RdDmaWriteData_o -> mm_interconnect_0:pcie_256_dma_dma_rd_master_writedata
	wire    [4:0] pcie_256_dma_dma_rd_master_burstcount;                             // pcie_256_dma:RdDmaBurstCount_o -> mm_interconnect_0:pcie_256_dma_dma_rd_master_burstcount
	wire          pcie_256_dma_dma_wr_master_waitrequest;                            // mm_interconnect_0:pcie_256_dma_dma_wr_master_waitrequest -> pcie_256_dma:WrDmaWaitRequest_i
	wire  [255:0] pcie_256_dma_dma_wr_master_readdata;                               // mm_interconnect_0:pcie_256_dma_dma_wr_master_readdata -> pcie_256_dma:WrDmaReadData_i
	wire   [63:0] pcie_256_dma_dma_wr_master_address;                                // pcie_256_dma:WrDmaAddress_o -> mm_interconnect_0:pcie_256_dma_dma_wr_master_address
	wire          pcie_256_dma_dma_wr_master_read;                                   // pcie_256_dma:WrDmaRead_o -> mm_interconnect_0:pcie_256_dma_dma_wr_master_read
	wire   [31:0] pcie_256_dma_dma_wr_master_byteenable;                             // pcie_256_dma:WrDmaByteEnable_o -> mm_interconnect_0:pcie_256_dma_dma_wr_master_byteenable
	wire          pcie_256_dma_dma_wr_master_readdatavalid;                          // mm_interconnect_0:pcie_256_dma_dma_wr_master_readdatavalid -> pcie_256_dma:WrDmaReadDataValid_i
	wire    [4:0] pcie_256_dma_dma_wr_master_burstcount;                             // pcie_256_dma:WrDmaBurstCount_o -> mm_interconnect_0:pcie_256_dma_dma_wr_master_burstcount
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect;                  // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                    // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;                     // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                  // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;                       // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                   // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;                       // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire          mm_interconnect_0_pio_led_s1_chipselect;                           // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire   [31:0] mm_interconnect_0_pio_led_s1_readdata;                             // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire    [1:0] mm_interconnect_0_pio_led_s1_address;                              // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire          mm_interconnect_0_pio_led_s1_write;                                // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire   [31:0] mm_interconnect_0_pio_led_s1_writedata;                            // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire   [31:0] mm_interconnect_0_pio_button_s1_readdata;                          // pio_button:readdata -> mm_interconnect_0:pio_button_s1_readdata
	wire    [1:0] mm_interconnect_0_pio_button_s1_address;                           // mm_interconnect_0:pio_button_s1_address -> pio_button:address
	wire   [31:0] mm_interconnect_0_ddr3a_status_s1_readdata;                        // ddr3a_status:readdata -> mm_interconnect_0:ddr3a_status_s1_readdata
	wire    [1:0] mm_interconnect_0_ddr3a_status_s1_address;                         // mm_interconnect_0:ddr3a_status_s1_address -> ddr3a_status:address
	wire   [31:0] mm_interconnect_0_ddr3b_status_s1_readdata;                        // ddr3b_status:readdata -> mm_interconnect_0:ddr3b_status_s1_readdata
	wire    [1:0] mm_interconnect_0_ddr3b_status_s1_address;                         // mm_interconnect_0:ddr3b_status_s1_address -> ddr3b_status:address
	wire          mm_interconnect_0_pcie_256_dma_rd_dts_slave_chipselect;            // mm_interconnect_0:pcie_256_dma_rd_dts_slave_chipselect -> pcie_256_dma:RdDTSChipSelect_i
	wire          mm_interconnect_0_pcie_256_dma_rd_dts_slave_waitrequest;           // pcie_256_dma:RdDTSWaitRequest_o -> mm_interconnect_0:pcie_256_dma_rd_dts_slave_waitrequest
	wire    [7:0] mm_interconnect_0_pcie_256_dma_rd_dts_slave_address;               // mm_interconnect_0:pcie_256_dma_rd_dts_slave_address -> pcie_256_dma:RdDTSAddress_i
	wire          mm_interconnect_0_pcie_256_dma_rd_dts_slave_write;                 // mm_interconnect_0:pcie_256_dma_rd_dts_slave_write -> pcie_256_dma:RdDTSWrite_i
	wire  [255:0] mm_interconnect_0_pcie_256_dma_rd_dts_slave_writedata;             // mm_interconnect_0:pcie_256_dma_rd_dts_slave_writedata -> pcie_256_dma:RdDTSWriteData_i
	wire    [4:0] mm_interconnect_0_pcie_256_dma_rd_dts_slave_burstcount;            // mm_interconnect_0:pcie_256_dma_rd_dts_slave_burstcount -> pcie_256_dma:RdDTSBurstCount_i
	wire  [511:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_readdata;      // mm_clock_crossing_bridge_ddr3a:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_readdata
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_waitrequest;   // mm_clock_crossing_bridge_ddr3a:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_waitrequest
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_debugaccess -> mm_clock_crossing_bridge_ddr3a:s0_debugaccess
	wire   [30:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_address -> mm_clock_crossing_bridge_ddr3a:s0_address
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_read -> mm_clock_crossing_bridge_ddr3a:s0_read
	wire   [63:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_byteenable -> mm_clock_crossing_bridge_ddr3a:s0_byteenable
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_readdatavalid; // mm_clock_crossing_bridge_ddr3a:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_readdatavalid
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_write -> mm_clock_crossing_bridge_ddr3a:s0_write
	wire  [511:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_writedata -> mm_clock_crossing_bridge_ddr3a:s0_writedata
	wire    [7:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_burstcount -> mm_clock_crossing_bridge_ddr3a:s0_burstcount
	wire  [511:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_readdata;      // mm_clock_crossing_bridge_ddr3b:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_readdata
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_waitrequest;   // mm_clock_crossing_bridge_ddr3b:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_waitrequest
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_debugaccess -> mm_clock_crossing_bridge_ddr3b:s0_debugaccess
	wire   [30:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_address -> mm_clock_crossing_bridge_ddr3b:s0_address
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_read -> mm_clock_crossing_bridge_ddr3b:s0_read
	wire   [63:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_byteenable -> mm_clock_crossing_bridge_ddr3b:s0_byteenable
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_readdatavalid; // mm_clock_crossing_bridge_ddr3b:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_readdatavalid
	wire          mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_write -> mm_clock_crossing_bridge_ddr3b:s0_write
	wire  [511:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_writedata -> mm_clock_crossing_bridge_ddr3b:s0_writedata
	wire    [7:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_ddr3b_s0_burstcount -> mm_clock_crossing_bridge_ddr3b:s0_burstcount
	wire          mm_interconnect_0_pcie_256_dma_wr_dts_slave_chipselect;            // mm_interconnect_0:pcie_256_dma_wr_dts_slave_chipselect -> pcie_256_dma:WrDTSChipSelect_i
	wire          mm_interconnect_0_pcie_256_dma_wr_dts_slave_waitrequest;           // pcie_256_dma:WrDTSWaitRequest_o -> mm_interconnect_0:pcie_256_dma_wr_dts_slave_waitrequest
	wire    [7:0] mm_interconnect_0_pcie_256_dma_wr_dts_slave_address;               // mm_interconnect_0:pcie_256_dma_wr_dts_slave_address -> pcie_256_dma:WrDTSAddress_i
	wire          mm_interconnect_0_pcie_256_dma_wr_dts_slave_write;                 // mm_interconnect_0:pcie_256_dma_wr_dts_slave_write -> pcie_256_dma:WrDTSWrite_i
	wire  [255:0] mm_interconnect_0_pcie_256_dma_wr_dts_slave_writedata;             // mm_interconnect_0:pcie_256_dma_wr_dts_slave_writedata -> pcie_256_dma:WrDTSWriteData_i
	wire    [4:0] mm_interconnect_0_pcie_256_dma_wr_dts_slave_burstcount;            // mm_interconnect_0:pcie_256_dma_wr_dts_slave_burstcount -> pcie_256_dma:WrDTSBurstCount_i
	wire          mm_interconnect_0_onchip_memory2_0_s2_chipselect;                  // mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s2_readdata;                    // onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	wire   [13:0] mm_interconnect_0_onchip_memory2_0_s2_address;                     // mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	wire   [31:0] mm_interconnect_0_onchip_memory2_0_s2_byteenable;                  // mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	wire          mm_interconnect_0_onchip_memory2_0_s2_write;                       // mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	wire  [255:0] mm_interconnect_0_onchip_memory2_0_s2_writedata;                   // mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	wire          mm_interconnect_0_onchip_memory2_0_s2_clken;                       // mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	wire          mm_clock_crossing_bridge_ddr3a_m0_waitrequest;                     // mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_waitrequest -> mm_clock_crossing_bridge_ddr3a:m0_waitrequest
	wire  [511:0] mm_clock_crossing_bridge_ddr3a_m0_readdata;                        // mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_readdata -> mm_clock_crossing_bridge_ddr3a:m0_readdata
	wire          mm_clock_crossing_bridge_ddr3a_m0_debugaccess;                     // mm_clock_crossing_bridge_ddr3a:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_debugaccess
	wire   [30:0] mm_clock_crossing_bridge_ddr3a_m0_address;                         // mm_clock_crossing_bridge_ddr3a:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_address
	wire          mm_clock_crossing_bridge_ddr3a_m0_read;                            // mm_clock_crossing_bridge_ddr3a:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_read
	wire   [63:0] mm_clock_crossing_bridge_ddr3a_m0_byteenable;                      // mm_clock_crossing_bridge_ddr3a:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_byteenable
	wire          mm_clock_crossing_bridge_ddr3a_m0_readdatavalid;                   // mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_readdatavalid -> mm_clock_crossing_bridge_ddr3a:m0_readdatavalid
	wire  [511:0] mm_clock_crossing_bridge_ddr3a_m0_writedata;                       // mm_clock_crossing_bridge_ddr3a:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_writedata
	wire          mm_clock_crossing_bridge_ddr3a_m0_write;                           // mm_clock_crossing_bridge_ddr3a:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_write
	wire    [7:0] mm_clock_crossing_bridge_ddr3a_m0_burstcount;                      // mm_clock_crossing_bridge_ddr3a:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_burstcount
	wire          mm_interconnect_1_mem_if_ddr3a_avl_beginbursttransfer;             // mm_interconnect_1:mem_if_ddr3a_avl_beginbursttransfer -> mem_if_ddr3a:avl_burstbegin
	wire  [511:0] mm_interconnect_1_mem_if_ddr3a_avl_readdata;                       // mem_if_ddr3a:avl_rdata -> mm_interconnect_1:mem_if_ddr3a_avl_readdata
	wire          mm_interconnect_1_mem_if_ddr3a_avl_waitrequest;                    // mem_if_ddr3a:avl_ready -> mm_interconnect_1:mem_if_ddr3a_avl_waitrequest
	wire   [24:0] mm_interconnect_1_mem_if_ddr3a_avl_address;                        // mm_interconnect_1:mem_if_ddr3a_avl_address -> mem_if_ddr3a:avl_addr
	wire          mm_interconnect_1_mem_if_ddr3a_avl_read;                           // mm_interconnect_1:mem_if_ddr3a_avl_read -> mem_if_ddr3a:avl_read_req
	wire   [63:0] mm_interconnect_1_mem_if_ddr3a_avl_byteenable;                     // mm_interconnect_1:mem_if_ddr3a_avl_byteenable -> mem_if_ddr3a:avl_be
	wire          mm_interconnect_1_mem_if_ddr3a_avl_readdatavalid;                  // mem_if_ddr3a:avl_rdata_valid -> mm_interconnect_1:mem_if_ddr3a_avl_readdatavalid
	wire          mm_interconnect_1_mem_if_ddr3a_avl_write;                          // mm_interconnect_1:mem_if_ddr3a_avl_write -> mem_if_ddr3a:avl_write_req
	wire  [511:0] mm_interconnect_1_mem_if_ddr3a_avl_writedata;                      // mm_interconnect_1:mem_if_ddr3a_avl_writedata -> mem_if_ddr3a:avl_wdata
	wire    [2:0] mm_interconnect_1_mem_if_ddr3a_avl_burstcount;                     // mm_interconnect_1:mem_if_ddr3a_avl_burstcount -> mem_if_ddr3a:avl_size
	wire          mm_clock_crossing_bridge_ddr3b_m0_waitrequest;                     // mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_waitrequest -> mm_clock_crossing_bridge_ddr3b:m0_waitrequest
	wire  [511:0] mm_clock_crossing_bridge_ddr3b_m0_readdata;                        // mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_readdata -> mm_clock_crossing_bridge_ddr3b:m0_readdata
	wire          mm_clock_crossing_bridge_ddr3b_m0_debugaccess;                     // mm_clock_crossing_bridge_ddr3b:m0_debugaccess -> mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_debugaccess
	wire   [30:0] mm_clock_crossing_bridge_ddr3b_m0_address;                         // mm_clock_crossing_bridge_ddr3b:m0_address -> mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_address
	wire          mm_clock_crossing_bridge_ddr3b_m0_read;                            // mm_clock_crossing_bridge_ddr3b:m0_read -> mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_read
	wire   [63:0] mm_clock_crossing_bridge_ddr3b_m0_byteenable;                      // mm_clock_crossing_bridge_ddr3b:m0_byteenable -> mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_byteenable
	wire          mm_clock_crossing_bridge_ddr3b_m0_readdatavalid;                   // mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_readdatavalid -> mm_clock_crossing_bridge_ddr3b:m0_readdatavalid
	wire  [511:0] mm_clock_crossing_bridge_ddr3b_m0_writedata;                       // mm_clock_crossing_bridge_ddr3b:m0_writedata -> mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_writedata
	wire          mm_clock_crossing_bridge_ddr3b_m0_write;                           // mm_clock_crossing_bridge_ddr3b:m0_write -> mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_write
	wire    [7:0] mm_clock_crossing_bridge_ddr3b_m0_burstcount;                      // mm_clock_crossing_bridge_ddr3b:m0_burstcount -> mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_burstcount
	wire          mm_interconnect_2_mem_if_ddr3b_avl_beginbursttransfer;             // mm_interconnect_2:mem_if_ddr3b_avl_beginbursttransfer -> mem_if_ddr3b:avl_burstbegin
	wire  [511:0] mm_interconnect_2_mem_if_ddr3b_avl_readdata;                       // mem_if_ddr3b:avl_rdata -> mm_interconnect_2:mem_if_ddr3b_avl_readdata
	wire          mm_interconnect_2_mem_if_ddr3b_avl_waitrequest;                    // mem_if_ddr3b:avl_ready -> mm_interconnect_2:mem_if_ddr3b_avl_waitrequest
	wire   [24:0] mm_interconnect_2_mem_if_ddr3b_avl_address;                        // mm_interconnect_2:mem_if_ddr3b_avl_address -> mem_if_ddr3b:avl_addr
	wire          mm_interconnect_2_mem_if_ddr3b_avl_read;                           // mm_interconnect_2:mem_if_ddr3b_avl_read -> mem_if_ddr3b:avl_read_req
	wire   [63:0] mm_interconnect_2_mem_if_ddr3b_avl_byteenable;                     // mm_interconnect_2:mem_if_ddr3b_avl_byteenable -> mem_if_ddr3b:avl_be
	wire          mm_interconnect_2_mem_if_ddr3b_avl_readdatavalid;                  // mem_if_ddr3b:avl_rdata_valid -> mm_interconnect_2:mem_if_ddr3b_avl_readdatavalid
	wire          mm_interconnect_2_mem_if_ddr3b_avl_write;                          // mm_interconnect_2:mem_if_ddr3b_avl_write -> mem_if_ddr3b:avl_write_req
	wire  [511:0] mm_interconnect_2_mem_if_ddr3b_avl_writedata;                      // mm_interconnect_2:mem_if_ddr3b_avl_writedata -> mem_if_ddr3b:avl_wdata
	wire    [2:0] mm_interconnect_2_mem_if_ddr3b_avl_burstcount;                     // mm_interconnect_2:mem_if_ddr3b_avl_burstcount -> mem_if_ddr3b:avl_size
	wire          pcie_256_dma_rd_dcm_master_waitrequest;                            // mm_interconnect_3:pcie_256_dma_rd_dcm_master_waitrequest -> pcie_256_dma:RdDCMWaitRequest_i
	wire   [31:0] pcie_256_dma_rd_dcm_master_readdata;                               // mm_interconnect_3:pcie_256_dma_rd_dcm_master_readdata -> pcie_256_dma:RdDCMReadData_i
	wire   [63:0] pcie_256_dma_rd_dcm_master_address;                                // pcie_256_dma:RdDCMAddress_o -> mm_interconnect_3:pcie_256_dma_rd_dcm_master_address
	wire          pcie_256_dma_rd_dcm_master_read;                                   // pcie_256_dma:RdDCMRead_o -> mm_interconnect_3:pcie_256_dma_rd_dcm_master_read
	wire    [3:0] pcie_256_dma_rd_dcm_master_byteenable;                             // pcie_256_dma:RdDCMByteEnable_o -> mm_interconnect_3:pcie_256_dma_rd_dcm_master_byteenable
	wire          pcie_256_dma_rd_dcm_master_readdatavalid;                          // mm_interconnect_3:pcie_256_dma_rd_dcm_master_readdatavalid -> pcie_256_dma:RdDCMReadDataValid_i
	wire          pcie_256_dma_rd_dcm_master_write;                                  // pcie_256_dma:RdDCMWrite_o -> mm_interconnect_3:pcie_256_dma_rd_dcm_master_write
	wire   [31:0] pcie_256_dma_rd_dcm_master_writedata;                              // pcie_256_dma:RdDCMWriteData_o -> mm_interconnect_3:pcie_256_dma_rd_dcm_master_writedata
	wire          pcie_256_dma_wr_dcm_master_waitrequest;                            // mm_interconnect_3:pcie_256_dma_wr_dcm_master_waitrequest -> pcie_256_dma:WrDCMWaitRequest_i
	wire   [31:0] pcie_256_dma_wr_dcm_master_readdata;                               // mm_interconnect_3:pcie_256_dma_wr_dcm_master_readdata -> pcie_256_dma:WrDCMReadData_i
	wire   [63:0] pcie_256_dma_wr_dcm_master_address;                                // pcie_256_dma:WrDCMAddress_o -> mm_interconnect_3:pcie_256_dma_wr_dcm_master_address
	wire          pcie_256_dma_wr_dcm_master_read;                                   // pcie_256_dma:WrDCMRead_o -> mm_interconnect_3:pcie_256_dma_wr_dcm_master_read
	wire    [3:0] pcie_256_dma_wr_dcm_master_byteenable;                             // pcie_256_dma:WrDCMByteEnable_o -> mm_interconnect_3:pcie_256_dma_wr_dcm_master_byteenable
	wire          pcie_256_dma_wr_dcm_master_readdatavalid;                          // mm_interconnect_3:pcie_256_dma_wr_dcm_master_readdatavalid -> pcie_256_dma:WrDCMReadDataValid_i
	wire          pcie_256_dma_wr_dcm_master_write;                                  // pcie_256_dma:WrDCMWrite_o -> mm_interconnect_3:pcie_256_dma_wr_dcm_master_write
	wire   [31:0] pcie_256_dma_wr_dcm_master_writedata;                              // pcie_256_dma:WrDCMWriteData_o -> mm_interconnect_3:pcie_256_dma_wr_dcm_master_writedata
	wire          mm_interconnect_3_pcie_256_dma_txs_chipselect;                     // mm_interconnect_3:pcie_256_dma_Txs_chipselect -> pcie_256_dma:TxsChipSelect_i
	wire   [31:0] mm_interconnect_3_pcie_256_dma_txs_readdata;                       // pcie_256_dma:TxsReadData_o -> mm_interconnect_3:pcie_256_dma_Txs_readdata
	wire          mm_interconnect_3_pcie_256_dma_txs_waitrequest;                    // pcie_256_dma:TxsWaitRequest_o -> mm_interconnect_3:pcie_256_dma_Txs_waitrequest
	wire   [63:0] mm_interconnect_3_pcie_256_dma_txs_address;                        // mm_interconnect_3:pcie_256_dma_Txs_address -> pcie_256_dma:TxsAddress_i
	wire          mm_interconnect_3_pcie_256_dma_txs_read;                           // mm_interconnect_3:pcie_256_dma_Txs_read -> pcie_256_dma:TxsRead_i
	wire    [3:0] mm_interconnect_3_pcie_256_dma_txs_byteenable;                     // mm_interconnect_3:pcie_256_dma_Txs_byteenable -> pcie_256_dma:TxsByteEnable_i
	wire          mm_interconnect_3_pcie_256_dma_txs_readdatavalid;                  // pcie_256_dma:TxsReadDataValid_o -> mm_interconnect_3:pcie_256_dma_Txs_readdatavalid
	wire          mm_interconnect_3_pcie_256_dma_txs_write;                          // mm_interconnect_3:pcie_256_dma_Txs_write -> pcie_256_dma:TxsWrite_i
	wire   [31:0] mm_interconnect_3_pcie_256_dma_txs_writedata;                      // mm_interconnect_3:pcie_256_dma_Txs_writedata -> pcie_256_dma:TxsWriteData_i
	wire          rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, pcie_reconfig_driver_0:reconfig_xcvr_rst]
	wire          rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [ddr3a_status:reset_n, ddr3b_status:reset_n, mm_interconnect_0:ddr3a_status_reset_reset_bridge_in_reset_reset]
	wire          pcie_256_dma_nreset_status_reset;                                  // pcie_256_dma:reset_status -> [rst_controller_001:reset_in0, rst_controller_005:reset_in0]
	wire          rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [mm_clock_crossing_bridge_ddr3a:m0_reset, mm_interconnect_1:mem_if_ddr3a_soft_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_clock_crossing_bridge_ddr3a_m0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                                // rst_controller_003:reset_out -> [mm_clock_crossing_bridge_ddr3a:s0_reset, mm_clock_crossing_bridge_ddr3b:s0_reset, mm_interconnect_0:mm_clock_crossing_bridge_ddr3a_s0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_004_reset_out_reset;                                // rst_controller_004:reset_out -> [mm_clock_crossing_bridge_ddr3b:m0_reset, mm_interconnect_2:mem_if_ddr3b_soft_reset_reset_bridge_in_reset_reset, mm_interconnect_2:mm_clock_crossing_bridge_ddr3b_m0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_005_reset_out_reset;                                // rst_controller_005:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, mm_interconnect_3:pcie_256_dma_rd_dcm_master_translator_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, onchip_memory2_0:reset2, pio_button:reset_n, pio_led:reset_n, rst_translator:in_reset]
	wire          rst_controller_005_reset_out_reset_req;                            // rst_controller_005:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator:reset_req_in]

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (11),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (1),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),       //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_clk),                                               //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                        //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),          //      reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),             //                   .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),         //                   .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest),      //                   .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),            //                   .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),        //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr), //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (pcie_256_dma_reconfig_from_xcvr_reconfig_from_xcvr),    // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                      //        (terminated)
		.rx_cal_busy               (),                                                      //        (terminated)
		.cal_busy_in               (1'b0),                                                  //        (terminated)
		.reconfig_mif_address      (),                                                      //        (terminated)
		.reconfig_mif_read         (),                                                      //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                  //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                   //        (terminated)
	);

	top_ddr3a_status ddr3a_status (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_ddr3a_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ddr3a_status_s1_readdata), //                    .readdata
		.in_port  (ddr3a_status_external_connection_export)     // external_connection.export
	);

	top_ddr3a_status ddr3b_status (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_ddr3b_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ddr3b_status_s1_readdata), //                    .readdata
		.in_port  (ddr3b_status_external_connection_export)     // external_connection.export
	);

	top_mem_if_ddr3a mem_if_ddr3a (
		.pll_ref_clk               (mem_if_ddr3a_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n            (reset_reset_n),                                         //     global_reset.reset_n
		.soft_reset_n              (reset_reset_n),                                         //       soft_reset.reset_n
		.afi_clk                   (mem_if_ddr3a_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                                      //     afi_half_clk.clk
		.afi_reset_n               (),                                                      //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                      // afi_reset_export.reset_n
		.mem_a                     (mem_if_ddr3a_mem_mem_a),                                //           memory.mem_a
		.mem_ba                    (mem_if_ddr3a_mem_mem_ba),                               //                 .mem_ba
		.mem_ck                    (mem_if_ddr3a_mem_mem_ck),                               //                 .mem_ck
		.mem_ck_n                  (mem_if_ddr3a_mem_mem_ck_n),                             //                 .mem_ck_n
		.mem_cke                   (mem_if_ddr3a_mem_mem_cke),                              //                 .mem_cke
		.mem_cs_n                  (mem_if_ddr3a_mem_mem_cs_n),                             //                 .mem_cs_n
		.mem_dm                    (mem_if_ddr3a_mem_mem_dm),                               //                 .mem_dm
		.mem_ras_n                 (mem_if_ddr3a_mem_mem_ras_n),                            //                 .mem_ras_n
		.mem_cas_n                 (mem_if_ddr3a_mem_mem_cas_n),                            //                 .mem_cas_n
		.mem_we_n                  (mem_if_ddr3a_mem_mem_we_n),                             //                 .mem_we_n
		.mem_reset_n               (mem_if_ddr3a_mem_mem_reset_n),                          //                 .mem_reset_n
		.mem_dq                    (mem_if_ddr3a_mem_mem_dq),                               //                 .mem_dq
		.mem_dqs                   (mem_if_ddr3a_mem_mem_dqs),                              //                 .mem_dqs
		.mem_dqs_n                 (mem_if_ddr3a_mem_mem_dqs_n),                            //                 .mem_dqs_n
		.mem_odt                   (mem_if_ddr3a_mem_mem_odt),                              //                 .mem_odt
		.avl_ready                 (mm_interconnect_1_mem_if_ddr3a_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_1_mem_if_ddr3a_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_1_mem_if_ddr3a_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_1_mem_if_ddr3a_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_1_mem_if_ddr3a_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_1_mem_if_ddr3a_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_1_mem_if_ddr3a_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_1_mem_if_ddr3a_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_1_mem_if_ddr3a_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_1_mem_if_ddr3a_avl_burstcount),         //                 .burstcount
		.local_init_done           (mem_if_ddr3a_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (mem_if_ddr3a_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (mem_if_ddr3a_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rzqin                 (mem_if_ddr3a_oct_rzqin),                                //              oct.rzqin
		.pll_mem_clk               (),                                                      //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                                      //                 .pll_write_clk
		.pll_locked                (),                                                      //                 .pll_locked
		.pll_write_clk_pre_phy_clk (),                                                      //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                                      //                 .pll_addr_cmd_clk
		.pll_avl_clk               (),                                                      //                 .pll_avl_clk
		.pll_config_clk            (),                                                      //                 .pll_config_clk
		.pll_hr_clk                (),                                                      //                 .pll_hr_clk
		.pll_p2c_read_clk          (),                                                      //                 .pll_p2c_read_clk
		.pll_c2p_write_clk         ()                                                       //                 .pll_c2p_write_clk
	);

	top_mem_if_ddr3b mem_if_ddr3b (
		.pll_ref_clk               (mem_if_ddr3b_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n            (reset_reset_n),                                         //     global_reset.reset_n
		.soft_reset_n              (reset_reset_n),                                         //       soft_reset.reset_n
		.afi_clk                   (mem_if_ddr3b_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                                      //     afi_half_clk.clk
		.afi_reset_n               (),                                                      //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                      // afi_reset_export.reset_n
		.mem_a                     (mem_if_ddr3b_mem_mem_a),                                //           memory.mem_a
		.mem_ba                    (mem_if_ddr3b_mem_mem_ba),                               //                 .mem_ba
		.mem_ck                    (mem_if_ddr3b_mem_mem_ck),                               //                 .mem_ck
		.mem_ck_n                  (mem_if_ddr3b_mem_mem_ck_n),                             //                 .mem_ck_n
		.mem_cke                   (mem_if_ddr3b_mem_mem_cke),                              //                 .mem_cke
		.mem_cs_n                  (mem_if_ddr3b_mem_mem_cs_n),                             //                 .mem_cs_n
		.mem_dm                    (mem_if_ddr3b_mem_mem_dm),                               //                 .mem_dm
		.mem_ras_n                 (mem_if_ddr3b_mem_mem_ras_n),                            //                 .mem_ras_n
		.mem_cas_n                 (mem_if_ddr3b_mem_mem_cas_n),                            //                 .mem_cas_n
		.mem_we_n                  (mem_if_ddr3b_mem_mem_we_n),                             //                 .mem_we_n
		.mem_reset_n               (mem_if_ddr3b_mem_mem_reset_n),                          //                 .mem_reset_n
		.mem_dq                    (mem_if_ddr3b_mem_mem_dq),                               //                 .mem_dq
		.mem_dqs                   (mem_if_ddr3b_mem_mem_dqs),                              //                 .mem_dqs
		.mem_dqs_n                 (mem_if_ddr3b_mem_mem_dqs_n),                            //                 .mem_dqs_n
		.mem_odt                   (mem_if_ddr3b_mem_mem_odt),                              //                 .mem_odt
		.avl_ready                 (mm_interconnect_2_mem_if_ddr3b_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_2_mem_if_ddr3b_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_2_mem_if_ddr3b_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_2_mem_if_ddr3b_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_2_mem_if_ddr3b_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_2_mem_if_ddr3b_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_2_mem_if_ddr3b_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_2_mem_if_ddr3b_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_2_mem_if_ddr3b_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_2_mem_if_ddr3b_avl_burstcount),         //                 .burstcount
		.local_init_done           (mem_if_ddr3b_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (mem_if_ddr3b_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (mem_if_ddr3b_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rzqin                 (mem_if_ddr3b_oct_rzqin),                                //              oct.rzqin
		.pll_mem_clk               (),                                                      //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                                      //                 .pll_write_clk
		.pll_locked                (),                                                      //                 .pll_locked
		.pll_write_clk_pre_phy_clk (),                                                      //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                                      //                 .pll_addr_cmd_clk
		.pll_avl_clk               (),                                                      //                 .pll_avl_clk
		.pll_config_clk            (),                                                      //                 .pll_config_clk
		.pll_hr_clk                (),                                                      //                 .pll_hr_clk
		.pll_p2c_read_clk          (),                                                      //                 .pll_p2c_read_clk
		.pll_c2p_write_clk         ()                                                       //                 .pll_c2p_write_clk
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (512),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (31),
		.BURSTCOUNT_WIDTH    (8),
		.COMMAND_FIFO_DEPTH  (512),
		.RESPONSE_FIFO_DEPTH (512),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_ddr3a (
		.m0_clk           (mem_if_ddr3a_afi_clk_clk),                                          //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                                // m0_reset.reset
		.s0_clk           (pcie_256_dma_coreclkout_clk),                                       //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                                // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_ddr3a_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_ddr3a_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_ddr3a_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_ddr3a_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_ddr3a_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_ddr3a_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_ddr3a_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_ddr3a_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_ddr3a_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_ddr3a_m0_debugaccess)                      //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (512),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (31),
		.BURSTCOUNT_WIDTH    (8),
		.COMMAND_FIFO_DEPTH  (512),
		.RESPONSE_FIFO_DEPTH (512),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_ddr3b (
		.m0_clk           (mem_if_ddr3b_afi_clk_clk),                                          //   m0_clk.clk
		.m0_reset         (rst_controller_004_reset_out_reset),                                // m0_reset.reset
		.s0_clk           (pcie_256_dma_coreclkout_clk),                                       //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                                // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_ddr3b_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_ddr3b_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_ddr3b_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_ddr3b_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_ddr3b_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_ddr3b_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_ddr3b_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_ddr3b_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_ddr3b_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_ddr3b_m0_debugaccess)                      //         .debugaccess
	);

	top_onchip_memory2_0 onchip_memory2_0 (
		.clk         (pcie_256_dma_coreclkout_clk),                      //   clk1.clk
		.address     (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset       (rst_controller_005_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_005_reset_out_reset_req),           //       .reset_req
		.address2    (mm_interconnect_0_onchip_memory2_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory2_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory2_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory2_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory2_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory2_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory2_0_s2_byteenable), //       .byteenable
		.clk2        (pcie_256_dma_coreclkout_clk),                      //   clk2.clk
		.reset2      (rst_controller_005_reset_out_reset),               // reset2.reset
		.reset_req2  (rst_controller_005_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	altpcie_256_hip_avmm_hwtcl #(
		.INTENDED_DEVICE_FAMILY                   ("Stratix V"),
		.lane_mask_hwtcl                          ("x8"),
		.gen123_lane_rate_mode_hwtcl              ("Gen3 (8.0 Gbps)"),
		.DMA_WIDTH                                (256),
		.DMA_BE_WIDTH                             (32),
		.DMA_BRST_CNT_W                           (5),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("3.0"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.internal_controller_hwtcl                (1),
		.enable_cra_hwtcl                         (1),
		.enable_rxm_burst_hwtcl                   (0),
		.in_cvp_mode_hwtcl                        (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.use_atx_pll_hwtcl                        (0),
		.dma_use_scfifo_ext_hwtcl                 (0),
		.bar0_type_hwtcl                          (64),
		.bar0_size_mask_hwtcl                     (9),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Enabled"),
		.bar0_prefetchable_hwtcl                  ("Enabled"),
		.bar1_type_hwtcl                          (1),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_type_hwtcl                          (1),
		.bar2_size_mask_hwtcl                     (0),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_type_hwtcl                          (1),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_type_hwtcl                          (64),
		.bar4_size_mask_hwtcl                     (27),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Enabled"),
		.bar4_prefetchable_hwtcl                  ("Enabled"),
		.bar5_type_hwtcl                          (1),
		.bar5_size_mask_hwtcl                     (0),
		.rd_dma_size_mask_hwtcl                   (34),
		.wr_dma_size_mask_hwtcl                   (34),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.vendor_id_hwtcl                          (4466),
		.device_id_hwtcl                          (57347),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (0),
		.subsystem_vendor_id_hwtcl                (4369),
		.subsystem_device_id_hwtcl                (13409),
		.max_payload_size_hwtcl                   (256),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("1"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.avmm_width_hwtcl                         (256),
		.avmm_burst_width_hwtcl                   (7),
		.TX_S_ADDR_WIDTH                          (64),
		.ast_width_hwtcl                          ("Avalon-ST 256-bit"),
		.use_ast_parity                           (0),
		.millisecond_cycle_count_hwtcl            (248500),
		.set_pll_coreclkout_cout_hwtcl            ("NA"),
		.set_pll_coreclkout_cin_hwtcl             ("NA"),
		.port_width_be_hwtcl                      (32),
		.port_width_data_hwtcl                    (256),
		.hip_reconfig_hwtcl                       (0),
		.vsec_id_hwtcl                            (40960),
		.vsec_rev_hwtcl                           (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("true"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (195),
		.cpl_spc_data_hwtcl                       (781),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (770),
		.reconfig_from_xcvr_width                 (506),
		.single_rx_detect_hwtcl                   (0),
		.hip_hard_reset_hwtcl                     (0),
		.use_cvp_update_core_pof_hwtcl            (0),
		.pcie_inspector_hwtcl                     (0),
		.tlp_inspector_hwtcl                      (0),
		.tlp_inspector_use_signal_probe_hwtcl     (0),
		.tlp_insp_trg_dw0_hwtcl                   (2049),
		.tlp_insp_trg_dw1_hwtcl                   (0),
		.tlp_insp_trg_dw2_hwtcl                   (0),
		.tlp_insp_trg_dw3_hwtcl                   (0),
		.use_tl_cfg_sync_hwtcl                    (1),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15),
		.av_rpre_emph_a_val_hwtcl                 (12),
		.av_rpre_emph_b_val_hwtcl                 (0),
		.av_rpre_emph_c_val_hwtcl                 (19),
		.av_rpre_emph_d_val_hwtcl                 (13),
		.av_rpre_emph_e_val_hwtcl                 (21),
		.av_rvod_sel_a_val_hwtcl                  (42),
		.av_rvod_sel_b_val_hwtcl                  (30),
		.av_rvod_sel_c_val_hwtcl                  (43),
		.av_rvod_sel_d_val_hwtcl                  (43),
		.av_rvod_sel_e_val_hwtcl                  (9),
		.cv_rpre_emph_a_val_hwtcl                 (11),
		.cv_rpre_emph_b_val_hwtcl                 (0),
		.cv_rpre_emph_c_val_hwtcl                 (22),
		.cv_rpre_emph_d_val_hwtcl                 (12),
		.cv_rpre_emph_e_val_hwtcl                 (21),
		.cv_rvod_sel_a_val_hwtcl                  (50),
		.cv_rvod_sel_b_val_hwtcl                  (34),
		.cv_rvod_sel_c_val_hwtcl                  (50),
		.cv_rvod_sel_d_val_hwtcl                  (50),
		.cv_rvod_sel_e_val_hwtcl                  (9)
	) pcie_256_dma (
		.coreclkout           (pcie_256_dma_coreclkout_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //          coreclkout.clk
		.refclk               (refclk_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //              refclk.clk
		.npor                 (pcie_rstn_npor),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                npor.npor
		.pin_perst            (pcie_rstn_pin_perst),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .pin_perst
		.reset_status         (pcie_256_dma_nreset_status_reset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //       nreset_status.reset_n
		.RxmAddress_4_o       (pcie_256_dma_rxm_bar4_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //            Rxm_BAR4.address
		.RxmRead_4_o          (pcie_256_dma_rxm_bar4_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                    .read
		.RxmWaitRequest_4_i   (pcie_256_dma_rxm_bar4_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .waitrequest
		.RxmWrite_4_o         (pcie_256_dma_rxm_bar4_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .write
		.RxmReadDataValid_4_i (pcie_256_dma_rxm_bar4_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .readdatavalid
		.RxmReadData_4_i      (pcie_256_dma_rxm_bar4_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .readdata
		.RxmWriteData_4_o     (pcie_256_dma_rxm_bar4_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .writedata
		.RxmByteEnable_4_o    (pcie_256_dma_rxm_bar4_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .byteenable
		.TxsAddress_i         (mm_interconnect_3_pcie_256_dma_txs_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                 Txs.address
		.TxsChipSelect_i      (mm_interconnect_3_pcie_256_dma_txs_chipselect),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                    .chipselect
		.TxsByteEnable_i      (mm_interconnect_3_pcie_256_dma_txs_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                    .byteenable
		.TxsReadData_o        (mm_interconnect_3_pcie_256_dma_txs_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .readdata
		.TxsWriteData_i       (mm_interconnect_3_pcie_256_dma_txs_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                    .writedata
		.TxsRead_i            (mm_interconnect_3_pcie_256_dma_txs_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .read
		.TxsWrite_i           (mm_interconnect_3_pcie_256_dma_txs_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .write
		.TxsReadDataValid_o   (mm_interconnect_3_pcie_256_dma_txs_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .readdatavalid
		.TxsWaitRequest_o     (mm_interconnect_3_pcie_256_dma_txs_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .waitrequest
		.CraChipSelect_i      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                 Cra.chipselect
		.CraAddress_i         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .address
		.CraByteEnable_i      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .byteenable
		.CraRead              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .read
		.CraReadData_o        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .readdata
		.CraWrite             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .write
		.CraWriteData_i       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .writedata
		.CraWaitRequest_o     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .waitrequest
		.RdDmaAddress_o       (pcie_256_dma_dma_rd_master_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //       dma_rd_master.address
		.RdDmaWrite_o         (pcie_256_dma_dma_rd_master_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .write
		.RdDmaWriteData_o     (pcie_256_dma_dma_rd_master_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .writedata
		.RdDmaWaitRequest_i   (pcie_256_dma_dma_rd_master_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .waitrequest
		.RdDmaBurstCount_o    (pcie_256_dma_dma_rd_master_burstcount),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .burstcount
		.RdDmaWriteEnable_o   (pcie_256_dma_dma_rd_master_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .byteenable
		.WrDmaAddress_o       (pcie_256_dma_dma_wr_master_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //       dma_wr_master.address
		.WrDmaRead_o          (pcie_256_dma_dma_wr_master_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .read
		.WrDmaWaitRequest_i   (pcie_256_dma_dma_wr_master_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .waitrequest
		.WrDmaBurstCount_o    (pcie_256_dma_dma_wr_master_burstcount),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .burstcount
		.WrDmaReadDataValid_i (pcie_256_dma_dma_wr_master_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .readdatavalid
		.WrDmaReadData_i      (pcie_256_dma_dma_wr_master_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .readdata
		.WrDmaByteEnable_o    (pcie_256_dma_dma_wr_master_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .byteenable
		.WrDTSChipSelect_i    (mm_interconnect_0_pcie_256_dma_wr_dts_slave_chipselect),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        wr_dts_slave.chipselect
		.WrDTSWrite_i         (mm_interconnect_0_pcie_256_dma_wr_dts_slave_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .write
		.WrDTSBurstCount_i    (mm_interconnect_0_pcie_256_dma_wr_dts_slave_burstcount),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .burstcount
		.WrDTSAddress_i       (mm_interconnect_0_pcie_256_dma_wr_dts_slave_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .address
		.WrDTSWriteData_i     (mm_interconnect_0_pcie_256_dma_wr_dts_slave_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .writedata
		.WrDTSWaitRequest_o   (mm_interconnect_0_pcie_256_dma_wr_dts_slave_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .waitrequest
		.RdDTSChipSelect_i    (mm_interconnect_0_pcie_256_dma_rd_dts_slave_chipselect),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        rd_dts_slave.chipselect
		.RdDTSWrite_i         (mm_interconnect_0_pcie_256_dma_rd_dts_slave_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .write
		.RdDTSBurstCount_i    (mm_interconnect_0_pcie_256_dma_rd_dts_slave_burstcount),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .burstcount
		.RdDTSAddress_i       (mm_interconnect_0_pcie_256_dma_rd_dts_slave_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .address
		.RdDTSWriteData_i     (mm_interconnect_0_pcie_256_dma_rd_dts_slave_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .writedata
		.RdDTSWaitRequest_o   (mm_interconnect_0_pcie_256_dma_rd_dts_slave_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .waitrequest
		.WrDCMAddress_o       (pcie_256_dma_wr_dcm_master_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //       wr_dcm_master.address
		.WrDCMWrite_o         (pcie_256_dma_wr_dcm_master_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .write
		.WrDCMWriteData_o     (pcie_256_dma_wr_dcm_master_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .writedata
		.WrDCMRead_o          (pcie_256_dma_wr_dcm_master_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .read
		.WrDCMByteEnable_o    (pcie_256_dma_wr_dcm_master_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .byteenable
		.WrDCMWaitRequest_i   (pcie_256_dma_wr_dcm_master_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .waitrequest
		.WrDCMReadData_i      (pcie_256_dma_wr_dcm_master_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .readdata
		.WrDCMReadDataValid_i (pcie_256_dma_wr_dcm_master_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .readdatavalid
		.RdDCMAddress_o       (pcie_256_dma_rd_dcm_master_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //       rd_dcm_master.address
		.RdDCMWrite_o         (pcie_256_dma_rd_dcm_master_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .write
		.RdDCMWriteData_o     (pcie_256_dma_rd_dcm_master_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .writedata
		.RdDCMRead_o          (pcie_256_dma_rd_dcm_master_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .read
		.RdDCMByteEnable_o    (pcie_256_dma_rd_dcm_master_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .byteenable
		.RdDCMWaitRequest_i   (pcie_256_dma_rd_dcm_master_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .waitrequest
		.RdDCMReadData_i      (pcie_256_dma_rd_dcm_master_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .readdata
		.RdDCMReadDataValid_i (pcie_256_dma_rd_dcm_master_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .readdatavalid
		.IntxReq_i            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //      INTX_Interface.intx_req
		.IntxAck_o            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .intx_ack
		.MsiIntfc_o           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //       MSI_Interface.msi_intfc
		.MsixIntfc_o          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //      MSIX_Interface.msix_intfc
		.reconfig_to_xcvr     (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr   (pcie_256_dma_reconfig_from_xcvr_reconfig_from_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (pcie_256_hip_avmm_0_reconfig_clk_locked_fixedclk_locked),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (hip_serial_rx_in0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //          hip_serial.rx_in0
		.rx_in1               (hip_serial_rx_in1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in1
		.rx_in2               (hip_serial_rx_in2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in2
		.rx_in3               (hip_serial_rx_in3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in3
		.rx_in4               (hip_serial_rx_in4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in4
		.rx_in5               (hip_serial_rx_in5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in5
		.rx_in6               (hip_serial_rx_in6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in6
		.rx_in7               (hip_serial_rx_in7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in7
		.tx_out0              (hip_serial_tx_out0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out0
		.tx_out1              (hip_serial_tx_out1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out1
		.tx_out2              (hip_serial_tx_out2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out2
		.tx_out3              (hip_serial_tx_out3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out3
		.tx_out4              (hip_serial_tx_out4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out4
		.tx_out5              (hip_serial_tx_out5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out5
		.tx_out6              (hip_serial_tx_out6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out6
		.tx_out7              (hip_serial_tx_out7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out7
		.sim_pipe_pclk_in     (hip_pipe_sim_pipe_pclk_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (hip_pipe_sim_pipe_rate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .sim_pipe_rate
		.sim_ltssmstate       (hip_pipe_sim_ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .sim_ltssmstate
		.eidleinfersel0       (hip_pipe_eidleinfersel0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel0
		.eidleinfersel1       (hip_pipe_eidleinfersel1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel1
		.eidleinfersel2       (hip_pipe_eidleinfersel2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel2
		.eidleinfersel3       (hip_pipe_eidleinfersel3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel3
		.eidleinfersel4       (hip_pipe_eidleinfersel4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel4
		.eidleinfersel5       (hip_pipe_eidleinfersel5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel5
		.eidleinfersel6       (hip_pipe_eidleinfersel6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel6
		.eidleinfersel7       (hip_pipe_eidleinfersel7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel7
		.powerdown0           (hip_pipe_powerdown0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown0
		.powerdown1           (hip_pipe_powerdown1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown1
		.powerdown2           (hip_pipe_powerdown2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown2
		.powerdown3           (hip_pipe_powerdown3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown3
		.powerdown4           (hip_pipe_powerdown4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown4
		.powerdown5           (hip_pipe_powerdown5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown5
		.powerdown6           (hip_pipe_powerdown6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown6
		.powerdown7           (hip_pipe_powerdown7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown7
		.rxpolarity0          (hip_pipe_rxpolarity0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity0
		.rxpolarity1          (hip_pipe_rxpolarity1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity1
		.rxpolarity2          (hip_pipe_rxpolarity2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity2
		.rxpolarity3          (hip_pipe_rxpolarity3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity3
		.rxpolarity4          (hip_pipe_rxpolarity4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity4
		.rxpolarity5          (hip_pipe_rxpolarity5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity5
		.rxpolarity6          (hip_pipe_rxpolarity6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity6
		.rxpolarity7          (hip_pipe_rxpolarity7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity7
		.txcompl0             (hip_pipe_txcompl0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl0
		.txcompl1             (hip_pipe_txcompl1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl1
		.txcompl2             (hip_pipe_txcompl2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl2
		.txcompl3             (hip_pipe_txcompl3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl3
		.txcompl4             (hip_pipe_txcompl4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl4
		.txcompl5             (hip_pipe_txcompl5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl5
		.txcompl6             (hip_pipe_txcompl6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl6
		.txcompl7             (hip_pipe_txcompl7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl7
		.txdata0              (hip_pipe_txdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata0
		.txdata1              (hip_pipe_txdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata1
		.txdata2              (hip_pipe_txdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata2
		.txdata3              (hip_pipe_txdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata3
		.txdata4              (hip_pipe_txdata4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata4
		.txdata5              (hip_pipe_txdata5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata5
		.txdata6              (hip_pipe_txdata6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata6
		.txdata7              (hip_pipe_txdata7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata7
		.txdatak0             (hip_pipe_txdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak0
		.txdatak1             (hip_pipe_txdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak1
		.txdatak2             (hip_pipe_txdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak2
		.txdatak3             (hip_pipe_txdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak3
		.txdatak4             (hip_pipe_txdatak4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak4
		.txdatak5             (hip_pipe_txdatak5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak5
		.txdatak6             (hip_pipe_txdatak6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak6
		.txdatak7             (hip_pipe_txdatak7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak7
		.txdetectrx0          (hip_pipe_txdetectrx0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx0
		.txdetectrx1          (hip_pipe_txdetectrx1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx1
		.txdetectrx2          (hip_pipe_txdetectrx2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx2
		.txdetectrx3          (hip_pipe_txdetectrx3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx3
		.txdetectrx4          (hip_pipe_txdetectrx4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx4
		.txdetectrx5          (hip_pipe_txdetectrx5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx5
		.txdetectrx6          (hip_pipe_txdetectrx6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx6
		.txdetectrx7          (hip_pipe_txdetectrx7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx7
		.txelecidle0          (hip_pipe_txelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle0
		.txelecidle1          (hip_pipe_txelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle1
		.txelecidle2          (hip_pipe_txelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle2
		.txelecidle3          (hip_pipe_txelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle3
		.txelecidle4          (hip_pipe_txelecidle4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle4
		.txelecidle5          (hip_pipe_txelecidle5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle5
		.txelecidle6          (hip_pipe_txelecidle6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle6
		.txelecidle7          (hip_pipe_txelecidle7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle7
		.txdeemph0            (hip_pipe_txdeemph0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph0
		.txdeemph1            (hip_pipe_txdeemph1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph1
		.txdeemph2            (hip_pipe_txdeemph2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph2
		.txdeemph3            (hip_pipe_txdeemph3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph3
		.txdeemph4            (hip_pipe_txdeemph4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph4
		.txdeemph5            (hip_pipe_txdeemph5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph5
		.txdeemph6            (hip_pipe_txdeemph6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph6
		.txdeemph7            (hip_pipe_txdeemph7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph7
		.txmargin0            (hip_pipe_txmargin0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin0
		.txmargin1            (hip_pipe_txmargin1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin1
		.txmargin2            (hip_pipe_txmargin2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin2
		.txmargin3            (hip_pipe_txmargin3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin3
		.txmargin4            (hip_pipe_txmargin4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin4
		.txmargin5            (hip_pipe_txmargin5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin5
		.txmargin6            (hip_pipe_txmargin6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin6
		.txmargin7            (hip_pipe_txmargin7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin7
		.txswing0             (hip_pipe_txswing0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing0
		.txswing1             (hip_pipe_txswing1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing1
		.txswing2             (hip_pipe_txswing2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing2
		.txswing3             (hip_pipe_txswing3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing3
		.txswing4             (hip_pipe_txswing4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing4
		.txswing5             (hip_pipe_txswing5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing5
		.txswing6             (hip_pipe_txswing6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing6
		.txswing7             (hip_pipe_txswing7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing7
		.phystatus0           (hip_pipe_phystatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus0
		.phystatus1           (hip_pipe_phystatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus1
		.phystatus2           (hip_pipe_phystatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus2
		.phystatus3           (hip_pipe_phystatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus3
		.phystatus4           (hip_pipe_phystatus4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus4
		.phystatus5           (hip_pipe_phystatus5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus5
		.phystatus6           (hip_pipe_phystatus6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus6
		.phystatus7           (hip_pipe_phystatus7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus7
		.rxdata0              (hip_pipe_rxdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata0
		.rxdata1              (hip_pipe_rxdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata1
		.rxdata2              (hip_pipe_rxdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata2
		.rxdata3              (hip_pipe_rxdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata3
		.rxdata4              (hip_pipe_rxdata4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata4
		.rxdata5              (hip_pipe_rxdata5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata5
		.rxdata6              (hip_pipe_rxdata6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata6
		.rxdata7              (hip_pipe_rxdata7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata7
		.rxdatak0             (hip_pipe_rxdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak0
		.rxdatak1             (hip_pipe_rxdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak1
		.rxdatak2             (hip_pipe_rxdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak2
		.rxdatak3             (hip_pipe_rxdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak3
		.rxdatak4             (hip_pipe_rxdatak4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak4
		.rxdatak5             (hip_pipe_rxdatak5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak5
		.rxdatak6             (hip_pipe_rxdatak6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak6
		.rxdatak7             (hip_pipe_rxdatak7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak7
		.rxelecidle0          (hip_pipe_rxelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle0
		.rxelecidle1          (hip_pipe_rxelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle1
		.rxelecidle2          (hip_pipe_rxelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle2
		.rxelecidle3          (hip_pipe_rxelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle3
		.rxelecidle4          (hip_pipe_rxelecidle4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle4
		.rxelecidle5          (hip_pipe_rxelecidle5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle5
		.rxelecidle6          (hip_pipe_rxelecidle6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle6
		.rxelecidle7          (hip_pipe_rxelecidle7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle7
		.rxstatus0            (hip_pipe_rxstatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus0
		.rxstatus1            (hip_pipe_rxstatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus1
		.rxstatus2            (hip_pipe_rxstatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus2
		.rxstatus3            (hip_pipe_rxstatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus3
		.rxstatus4            (hip_pipe_rxstatus4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus4
		.rxstatus5            (hip_pipe_rxstatus5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus5
		.rxstatus6            (hip_pipe_rxstatus6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus6
		.rxstatus7            (hip_pipe_rxstatus7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus7
		.rxvalid0             (hip_pipe_rxvalid0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid0
		.rxvalid1             (hip_pipe_rxvalid1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid1
		.rxvalid2             (hip_pipe_rxvalid2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid2
		.rxvalid3             (hip_pipe_rxvalid3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid3
		.rxvalid4             (hip_pipe_rxvalid4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid4
		.rxvalid5             (hip_pipe_rxvalid5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid5
		.rxvalid6             (hip_pipe_rxvalid6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid6
		.rxvalid7             (hip_pipe_rxvalid7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid7
		.test_in              (hip_ctrl_test_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //            hip_ctrl.test_in
		.simu_mode_pipe       (hip_ctrl_simu_mode_pipe),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .simu_mode_pipe
		.derr_cor_ext_rcv     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //          hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .derr_cor_ext_rpl
		.derr_rpl             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .derr_rpl
		.dlup_exit            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .dlup_exit
		.ev128ns              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ev128ns
		.ev1us                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ev1us
		.hotrst_exit          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .hotrst_exit
		.int_status           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .int_status
		.l2_exit              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .l2_exit
		.lane_act             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .lane_act
		.ltssmstate           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ltssmstate
		.dlup                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .dlup
		.rx_par_err           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rx_par_err
		.tx_par_err           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .tx_par_err
		.cfg_par_err          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .cfg_par_err
		.ko_cpl_spc_header    (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ko_cpl_spc_header
		.ko_cpl_spc_data      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ko_cpl_spc_data
		.currentspeed         (pcie_256_dma_hip_currentspeed_currentspeed),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //    hip_currentspeed.currentspeed
		.tl_cfg_add           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           config_tl.tl_cfg_add
		.tl_cfg_ctl           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .tl_cfg_ctl
		.tl_cfg_sts           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .tl_cfg_sts
		.RdDmaRxValid_i       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.RdDmaRxData_i        (160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.RdDmaRxReady_o       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.RdDmaTxData_o        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.RdDmaTxValid_o       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.WrDmaRxValid_i       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.WrDmaRxData_i        (160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.WrDmaRxReady_o       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.WrDmaTxData_o        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.WrDmaTxValid_o       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rxdataskip0          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip1          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip2          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip3          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip4          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip5          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip6          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip7          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst0             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst1             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst2             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst3             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst4             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst5             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst6             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst7             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxsynchd0            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd1            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd2            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd3            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd4            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd5            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd6            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd7            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxfreqlocked0        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked1        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked2        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked3        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked4        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked5        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked6        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked7        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.currentcoeff0        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff1        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff2        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff3        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff4        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff5        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff6        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff7        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset0     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset1     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset2     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset3     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset4     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset5     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset6     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset7     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd0            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd1            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd2            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd3            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd4            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd5            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd6            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd7            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst0             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst1             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst2             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst3             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst4             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst5             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst6             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst7             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.tlbfm_in             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.tlbfm_out            (1001'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000)  //         (terminated)
	);

	altpcie_reconfig_driver #(
		.INTENDED_DEVICE_FAMILY        ("Stratix V"),
		.gen123_lane_rate_mode_hwtcl   ("Gen3 (8.0 Gbps)"),
		.number_of_reconfig_interfaces (11)
	) pcie_reconfig_driver_0 (
		.reconfig_xcvr_clk         (clk_clk),                                          // reconfig_xcvr_clk.clk
		.reconfig_xcvr_rst         (rst_controller_reset_out_reset),                   // reconfig_xcvr_rst.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),     //     reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),        //                  .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),    //                  .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest), //                  .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),       //                  .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),   //                  .writedata
		.currentspeed              (pcie_256_dma_hip_currentspeed_currentspeed),       //  hip_currentspeed.currentspeed
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),  //     reconfig_busy.reconfig_busy
		.pld_clk                   (pcie_256_dma_coreclkout_clk),                      //           pld_clk.clk
		.derr_cor_ext_rcv_drv      (),                                                 //    hip_status_drv.derr_cor_ext_rcv
		.derr_cor_ext_rpl_drv      (),                                                 //                  .derr_cor_ext_rpl
		.derr_rpl_drv              (),                                                 //                  .derr_rpl
		.dlup_exit_drv             (),                                                 //                  .dlup_exit
		.ev128ns_drv               (),                                                 //                  .ev128ns
		.ev1us_drv                 (),                                                 //                  .ev1us
		.hotrst_exit_drv           (),                                                 //                  .hotrst_exit
		.int_status_drv            (),                                                 //                  .int_status
		.l2_exit_drv               (),                                                 //                  .l2_exit
		.lane_act_drv              (),                                                 //                  .lane_act
		.ltssmstate_drv            (),                                                 //                  .ltssmstate
		.dlup_drv                  (),                                                 //                  .dlup
		.rx_par_err_drv            (),                                                 //                  .rx_par_err
		.tx_par_err_drv            (),                                                 //                  .tx_par_err
		.cfg_par_err_drv           (),                                                 //                  .cfg_par_err
		.ko_cpl_spc_header_drv     (),                                                 //                  .ko_cpl_spc_header
		.ko_cpl_spc_data_drv       (),                                                 //                  .ko_cpl_spc_data
		.cal_busy_in               ()                                                  //       (terminated)
	);

	top_pio_button pio_button (
		.clk      (pcie_256_dma_coreclkout_clk),              //                 clk.clk
		.reset_n  (~rst_controller_005_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_pio_button_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_button_s1_readdata), //                    .readdata
		.in_port  (pio_button_external_connection_export)     // external_connection.export
	);

	top_pio_led pio_led (
		.clk        (pcie_256_dma_coreclkout_clk),             //                 clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_external_connection_export)       // external_connection.export
	);

	top_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                       (clk_clk),                                                           //                                                     clk_0_clk.clk
		.pcie_256_dma_coreclkout_clk                                         (pcie_256_dma_coreclkout_clk),                                       //                                       pcie_256_dma_coreclkout.clk
		.ddr3a_status_reset_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),                                //                      ddr3a_status_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_ddr3a_s0_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                                // mm_clock_crossing_bridge_ddr3a_s0_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset                 (rst_controller_005_reset_out_reset),                                //                 onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.pcie_256_dma_dma_rd_master_address                                  (pcie_256_dma_dma_rd_master_address),                                //                                    pcie_256_dma_dma_rd_master.address
		.pcie_256_dma_dma_rd_master_waitrequest                              (pcie_256_dma_dma_rd_master_waitrequest),                            //                                                              .waitrequest
		.pcie_256_dma_dma_rd_master_burstcount                               (pcie_256_dma_dma_rd_master_burstcount),                             //                                                              .burstcount
		.pcie_256_dma_dma_rd_master_byteenable                               (pcie_256_dma_dma_rd_master_byteenable),                             //                                                              .byteenable
		.pcie_256_dma_dma_rd_master_write                                    (pcie_256_dma_dma_rd_master_write),                                  //                                                              .write
		.pcie_256_dma_dma_rd_master_writedata                                (pcie_256_dma_dma_rd_master_writedata),                              //                                                              .writedata
		.pcie_256_dma_dma_wr_master_address                                  (pcie_256_dma_dma_wr_master_address),                                //                                    pcie_256_dma_dma_wr_master.address
		.pcie_256_dma_dma_wr_master_waitrequest                              (pcie_256_dma_dma_wr_master_waitrequest),                            //                                                              .waitrequest
		.pcie_256_dma_dma_wr_master_burstcount                               (pcie_256_dma_dma_wr_master_burstcount),                             //                                                              .burstcount
		.pcie_256_dma_dma_wr_master_byteenable                               (pcie_256_dma_dma_wr_master_byteenable),                             //                                                              .byteenable
		.pcie_256_dma_dma_wr_master_read                                     (pcie_256_dma_dma_wr_master_read),                                   //                                                              .read
		.pcie_256_dma_dma_wr_master_readdata                                 (pcie_256_dma_dma_wr_master_readdata),                               //                                                              .readdata
		.pcie_256_dma_dma_wr_master_readdatavalid                            (pcie_256_dma_dma_wr_master_readdatavalid),                          //                                                              .readdatavalid
		.pcie_256_dma_Rxm_BAR4_address                                       (pcie_256_dma_rxm_bar4_address),                                     //                                         pcie_256_dma_Rxm_BAR4.address
		.pcie_256_dma_Rxm_BAR4_waitrequest                                   (pcie_256_dma_rxm_bar4_waitrequest),                                 //                                                              .waitrequest
		.pcie_256_dma_Rxm_BAR4_byteenable                                    (pcie_256_dma_rxm_bar4_byteenable),                                  //                                                              .byteenable
		.pcie_256_dma_Rxm_BAR4_read                                          (pcie_256_dma_rxm_bar4_read),                                        //                                                              .read
		.pcie_256_dma_Rxm_BAR4_readdata                                      (pcie_256_dma_rxm_bar4_readdata),                                    //                                                              .readdata
		.pcie_256_dma_Rxm_BAR4_readdatavalid                                 (pcie_256_dma_rxm_bar4_readdatavalid),                               //                                                              .readdatavalid
		.pcie_256_dma_Rxm_BAR4_write                                         (pcie_256_dma_rxm_bar4_write),                                       //                                                              .write
		.pcie_256_dma_Rxm_BAR4_writedata                                     (pcie_256_dma_rxm_bar4_writedata),                                   //                                                              .writedata
		.ddr3a_status_s1_address                                             (mm_interconnect_0_ddr3a_status_s1_address),                         //                                               ddr3a_status_s1.address
		.ddr3a_status_s1_readdata                                            (mm_interconnect_0_ddr3a_status_s1_readdata),                        //                                                              .readdata
		.ddr3b_status_s1_address                                             (mm_interconnect_0_ddr3b_status_s1_address),                         //                                               ddr3b_status_s1.address
		.ddr3b_status_s1_readdata                                            (mm_interconnect_0_ddr3b_status_s1_readdata),                        //                                                              .readdata
		.mm_clock_crossing_bridge_ddr3a_s0_address                           (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_address),       //                             mm_clock_crossing_bridge_ddr3a_s0.address
		.mm_clock_crossing_bridge_ddr3a_s0_write                             (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_write),         //                                                              .write
		.mm_clock_crossing_bridge_ddr3a_s0_read                              (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_read),          //                                                              .read
		.mm_clock_crossing_bridge_ddr3a_s0_readdata                          (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_readdata),      //                                                              .readdata
		.mm_clock_crossing_bridge_ddr3a_s0_writedata                         (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_writedata),     //                                                              .writedata
		.mm_clock_crossing_bridge_ddr3a_s0_burstcount                        (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_burstcount),    //                                                              .burstcount
		.mm_clock_crossing_bridge_ddr3a_s0_byteenable                        (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_byteenable),    //                                                              .byteenable
		.mm_clock_crossing_bridge_ddr3a_s0_readdatavalid                     (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_readdatavalid), //                                                              .readdatavalid
		.mm_clock_crossing_bridge_ddr3a_s0_waitrequest                       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_waitrequest),   //                                                              .waitrequest
		.mm_clock_crossing_bridge_ddr3a_s0_debugaccess                       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3a_s0_debugaccess),   //                                                              .debugaccess
		.mm_clock_crossing_bridge_ddr3b_s0_address                           (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_address),       //                             mm_clock_crossing_bridge_ddr3b_s0.address
		.mm_clock_crossing_bridge_ddr3b_s0_write                             (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_write),         //                                                              .write
		.mm_clock_crossing_bridge_ddr3b_s0_read                              (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_read),          //                                                              .read
		.mm_clock_crossing_bridge_ddr3b_s0_readdata                          (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_readdata),      //                                                              .readdata
		.mm_clock_crossing_bridge_ddr3b_s0_writedata                         (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_writedata),     //                                                              .writedata
		.mm_clock_crossing_bridge_ddr3b_s0_burstcount                        (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_burstcount),    //                                                              .burstcount
		.mm_clock_crossing_bridge_ddr3b_s0_byteenable                        (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_byteenable),    //                                                              .byteenable
		.mm_clock_crossing_bridge_ddr3b_s0_readdatavalid                     (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_readdatavalid), //                                                              .readdatavalid
		.mm_clock_crossing_bridge_ddr3b_s0_waitrequest                       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_waitrequest),   //                                                              .waitrequest
		.mm_clock_crossing_bridge_ddr3b_s0_debugaccess                       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3b_s0_debugaccess),   //                                                              .debugaccess
		.onchip_memory2_0_s1_address                                         (mm_interconnect_0_onchip_memory2_0_s1_address),                     //                                           onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                           (mm_interconnect_0_onchip_memory2_0_s1_write),                       //                                                              .write
		.onchip_memory2_0_s1_readdata                                        (mm_interconnect_0_onchip_memory2_0_s1_readdata),                    //                                                              .readdata
		.onchip_memory2_0_s1_writedata                                       (mm_interconnect_0_onchip_memory2_0_s1_writedata),                   //                                                              .writedata
		.onchip_memory2_0_s1_byteenable                                      (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                  //                                                              .byteenable
		.onchip_memory2_0_s1_chipselect                                      (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                  //                                                              .chipselect
		.onchip_memory2_0_s1_clken                                           (mm_interconnect_0_onchip_memory2_0_s1_clken),                       //                                                              .clken
		.onchip_memory2_0_s2_address                                         (mm_interconnect_0_onchip_memory2_0_s2_address),                     //                                           onchip_memory2_0_s2.address
		.onchip_memory2_0_s2_write                                           (mm_interconnect_0_onchip_memory2_0_s2_write),                       //                                                              .write
		.onchip_memory2_0_s2_readdata                                        (mm_interconnect_0_onchip_memory2_0_s2_readdata),                    //                                                              .readdata
		.onchip_memory2_0_s2_writedata                                       (mm_interconnect_0_onchip_memory2_0_s2_writedata),                   //                                                              .writedata
		.onchip_memory2_0_s2_byteenable                                      (mm_interconnect_0_onchip_memory2_0_s2_byteenable),                  //                                                              .byteenable
		.onchip_memory2_0_s2_chipselect                                      (mm_interconnect_0_onchip_memory2_0_s2_chipselect),                  //                                                              .chipselect
		.onchip_memory2_0_s2_clken                                           (mm_interconnect_0_onchip_memory2_0_s2_clken),                       //                                                              .clken
		.pcie_256_dma_rd_dts_slave_address                                   (mm_interconnect_0_pcie_256_dma_rd_dts_slave_address),               //                                     pcie_256_dma_rd_dts_slave.address
		.pcie_256_dma_rd_dts_slave_write                                     (mm_interconnect_0_pcie_256_dma_rd_dts_slave_write),                 //                                                              .write
		.pcie_256_dma_rd_dts_slave_writedata                                 (mm_interconnect_0_pcie_256_dma_rd_dts_slave_writedata),             //                                                              .writedata
		.pcie_256_dma_rd_dts_slave_burstcount                                (mm_interconnect_0_pcie_256_dma_rd_dts_slave_burstcount),            //                                                              .burstcount
		.pcie_256_dma_rd_dts_slave_waitrequest                               (mm_interconnect_0_pcie_256_dma_rd_dts_slave_waitrequest),           //                                                              .waitrequest
		.pcie_256_dma_rd_dts_slave_chipselect                                (mm_interconnect_0_pcie_256_dma_rd_dts_slave_chipselect),            //                                                              .chipselect
		.pcie_256_dma_wr_dts_slave_address                                   (mm_interconnect_0_pcie_256_dma_wr_dts_slave_address),               //                                     pcie_256_dma_wr_dts_slave.address
		.pcie_256_dma_wr_dts_slave_write                                     (mm_interconnect_0_pcie_256_dma_wr_dts_slave_write),                 //                                                              .write
		.pcie_256_dma_wr_dts_slave_writedata                                 (mm_interconnect_0_pcie_256_dma_wr_dts_slave_writedata),             //                                                              .writedata
		.pcie_256_dma_wr_dts_slave_burstcount                                (mm_interconnect_0_pcie_256_dma_wr_dts_slave_burstcount),            //                                                              .burstcount
		.pcie_256_dma_wr_dts_slave_waitrequest                               (mm_interconnect_0_pcie_256_dma_wr_dts_slave_waitrequest),           //                                                              .waitrequest
		.pcie_256_dma_wr_dts_slave_chipselect                                (mm_interconnect_0_pcie_256_dma_wr_dts_slave_chipselect),            //                                                              .chipselect
		.pio_button_s1_address                                               (mm_interconnect_0_pio_button_s1_address),                           //                                                 pio_button_s1.address
		.pio_button_s1_readdata                                              (mm_interconnect_0_pio_button_s1_readdata),                          //                                                              .readdata
		.pio_led_s1_address                                                  (mm_interconnect_0_pio_led_s1_address),                              //                                                    pio_led_s1.address
		.pio_led_s1_write                                                    (mm_interconnect_0_pio_led_s1_write),                                //                                                              .write
		.pio_led_s1_readdata                                                 (mm_interconnect_0_pio_led_s1_readdata),                             //                                                              .readdata
		.pio_led_s1_writedata                                                (mm_interconnect_0_pio_led_s1_writedata),                            //                                                              .writedata
		.pio_led_s1_chipselect                                               (mm_interconnect_0_pio_led_s1_chipselect)                            //                                                              .chipselect
	);

	top_mm_interconnect_1 mm_interconnect_1 (
		.mem_if_ddr3a_afi_clk_clk                                            (mem_if_ddr3a_afi_clk_clk),                              //                                          mem_if_ddr3a_afi_clk.clk
		.mem_if_ddr3a_soft_reset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                    //                 mem_if_ddr3a_soft_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_ddr3a_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                    // mm_clock_crossing_bridge_ddr3a_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_ddr3a_m0_address                           (mm_clock_crossing_bridge_ddr3a_m0_address),             //                             mm_clock_crossing_bridge_ddr3a_m0.address
		.mm_clock_crossing_bridge_ddr3a_m0_waitrequest                       (mm_clock_crossing_bridge_ddr3a_m0_waitrequest),         //                                                              .waitrequest
		.mm_clock_crossing_bridge_ddr3a_m0_burstcount                        (mm_clock_crossing_bridge_ddr3a_m0_burstcount),          //                                                              .burstcount
		.mm_clock_crossing_bridge_ddr3a_m0_byteenable                        (mm_clock_crossing_bridge_ddr3a_m0_byteenable),          //                                                              .byteenable
		.mm_clock_crossing_bridge_ddr3a_m0_read                              (mm_clock_crossing_bridge_ddr3a_m0_read),                //                                                              .read
		.mm_clock_crossing_bridge_ddr3a_m0_readdata                          (mm_clock_crossing_bridge_ddr3a_m0_readdata),            //                                                              .readdata
		.mm_clock_crossing_bridge_ddr3a_m0_readdatavalid                     (mm_clock_crossing_bridge_ddr3a_m0_readdatavalid),       //                                                              .readdatavalid
		.mm_clock_crossing_bridge_ddr3a_m0_write                             (mm_clock_crossing_bridge_ddr3a_m0_write),               //                                                              .write
		.mm_clock_crossing_bridge_ddr3a_m0_writedata                         (mm_clock_crossing_bridge_ddr3a_m0_writedata),           //                                                              .writedata
		.mm_clock_crossing_bridge_ddr3a_m0_debugaccess                       (mm_clock_crossing_bridge_ddr3a_m0_debugaccess),         //                                                              .debugaccess
		.mem_if_ddr3a_avl_address                                            (mm_interconnect_1_mem_if_ddr3a_avl_address),            //                                              mem_if_ddr3a_avl.address
		.mem_if_ddr3a_avl_write                                              (mm_interconnect_1_mem_if_ddr3a_avl_write),              //                                                              .write
		.mem_if_ddr3a_avl_read                                               (mm_interconnect_1_mem_if_ddr3a_avl_read),               //                                                              .read
		.mem_if_ddr3a_avl_readdata                                           (mm_interconnect_1_mem_if_ddr3a_avl_readdata),           //                                                              .readdata
		.mem_if_ddr3a_avl_writedata                                          (mm_interconnect_1_mem_if_ddr3a_avl_writedata),          //                                                              .writedata
		.mem_if_ddr3a_avl_beginbursttransfer                                 (mm_interconnect_1_mem_if_ddr3a_avl_beginbursttransfer), //                                                              .beginbursttransfer
		.mem_if_ddr3a_avl_burstcount                                         (mm_interconnect_1_mem_if_ddr3a_avl_burstcount),         //                                                              .burstcount
		.mem_if_ddr3a_avl_byteenable                                         (mm_interconnect_1_mem_if_ddr3a_avl_byteenable),         //                                                              .byteenable
		.mem_if_ddr3a_avl_readdatavalid                                      (mm_interconnect_1_mem_if_ddr3a_avl_readdatavalid),      //                                                              .readdatavalid
		.mem_if_ddr3a_avl_waitrequest                                        (~mm_interconnect_1_mem_if_ddr3a_avl_waitrequest)        //                                                              .waitrequest
	);

	top_mm_interconnect_2 mm_interconnect_2 (
		.mem_if_ddr3b_afi_clk_clk                                            (mem_if_ddr3b_afi_clk_clk),                              //                                          mem_if_ddr3b_afi_clk.clk
		.mem_if_ddr3b_soft_reset_reset_bridge_in_reset_reset                 (rst_controller_004_reset_out_reset),                    //                 mem_if_ddr3b_soft_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_ddr3b_m0_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                    // mm_clock_crossing_bridge_ddr3b_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_ddr3b_m0_address                           (mm_clock_crossing_bridge_ddr3b_m0_address),             //                             mm_clock_crossing_bridge_ddr3b_m0.address
		.mm_clock_crossing_bridge_ddr3b_m0_waitrequest                       (mm_clock_crossing_bridge_ddr3b_m0_waitrequest),         //                                                              .waitrequest
		.mm_clock_crossing_bridge_ddr3b_m0_burstcount                        (mm_clock_crossing_bridge_ddr3b_m0_burstcount),          //                                                              .burstcount
		.mm_clock_crossing_bridge_ddr3b_m0_byteenable                        (mm_clock_crossing_bridge_ddr3b_m0_byteenable),          //                                                              .byteenable
		.mm_clock_crossing_bridge_ddr3b_m0_read                              (mm_clock_crossing_bridge_ddr3b_m0_read),                //                                                              .read
		.mm_clock_crossing_bridge_ddr3b_m0_readdata                          (mm_clock_crossing_bridge_ddr3b_m0_readdata),            //                                                              .readdata
		.mm_clock_crossing_bridge_ddr3b_m0_readdatavalid                     (mm_clock_crossing_bridge_ddr3b_m0_readdatavalid),       //                                                              .readdatavalid
		.mm_clock_crossing_bridge_ddr3b_m0_write                             (mm_clock_crossing_bridge_ddr3b_m0_write),               //                                                              .write
		.mm_clock_crossing_bridge_ddr3b_m0_writedata                         (mm_clock_crossing_bridge_ddr3b_m0_writedata),           //                                                              .writedata
		.mm_clock_crossing_bridge_ddr3b_m0_debugaccess                       (mm_clock_crossing_bridge_ddr3b_m0_debugaccess),         //                                                              .debugaccess
		.mem_if_ddr3b_avl_address                                            (mm_interconnect_2_mem_if_ddr3b_avl_address),            //                                              mem_if_ddr3b_avl.address
		.mem_if_ddr3b_avl_write                                              (mm_interconnect_2_mem_if_ddr3b_avl_write),              //                                                              .write
		.mem_if_ddr3b_avl_read                                               (mm_interconnect_2_mem_if_ddr3b_avl_read),               //                                                              .read
		.mem_if_ddr3b_avl_readdata                                           (mm_interconnect_2_mem_if_ddr3b_avl_readdata),           //                                                              .readdata
		.mem_if_ddr3b_avl_writedata                                          (mm_interconnect_2_mem_if_ddr3b_avl_writedata),          //                                                              .writedata
		.mem_if_ddr3b_avl_beginbursttransfer                                 (mm_interconnect_2_mem_if_ddr3b_avl_beginbursttransfer), //                                                              .beginbursttransfer
		.mem_if_ddr3b_avl_burstcount                                         (mm_interconnect_2_mem_if_ddr3b_avl_burstcount),         //                                                              .burstcount
		.mem_if_ddr3b_avl_byteenable                                         (mm_interconnect_2_mem_if_ddr3b_avl_byteenable),         //                                                              .byteenable
		.mem_if_ddr3b_avl_readdatavalid                                      (mm_interconnect_2_mem_if_ddr3b_avl_readdatavalid),      //                                                              .readdatavalid
		.mem_if_ddr3b_avl_waitrequest                                        (~mm_interconnect_2_mem_if_ddr3b_avl_waitrequest)        //                                                              .waitrequest
	);

	top_mm_interconnect_3 mm_interconnect_3 (
		.pcie_256_dma_coreclkout_clk                                             (pcie_256_dma_coreclkout_clk),                      //                                           pcie_256_dma_coreclkout.clk
		.pcie_256_dma_rd_dcm_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),               // pcie_256_dma_rd_dcm_master_translator_reset_reset_bridge_in_reset.reset
		.pcie_256_dma_rd_dcm_master_address                                      (pcie_256_dma_rd_dcm_master_address),               //                                        pcie_256_dma_rd_dcm_master.address
		.pcie_256_dma_rd_dcm_master_waitrequest                                  (pcie_256_dma_rd_dcm_master_waitrequest),           //                                                                  .waitrequest
		.pcie_256_dma_rd_dcm_master_byteenable                                   (pcie_256_dma_rd_dcm_master_byteenable),            //                                                                  .byteenable
		.pcie_256_dma_rd_dcm_master_read                                         (pcie_256_dma_rd_dcm_master_read),                  //                                                                  .read
		.pcie_256_dma_rd_dcm_master_readdata                                     (pcie_256_dma_rd_dcm_master_readdata),              //                                                                  .readdata
		.pcie_256_dma_rd_dcm_master_readdatavalid                                (pcie_256_dma_rd_dcm_master_readdatavalid),         //                                                                  .readdatavalid
		.pcie_256_dma_rd_dcm_master_write                                        (pcie_256_dma_rd_dcm_master_write),                 //                                                                  .write
		.pcie_256_dma_rd_dcm_master_writedata                                    (pcie_256_dma_rd_dcm_master_writedata),             //                                                                  .writedata
		.pcie_256_dma_wr_dcm_master_address                                      (pcie_256_dma_wr_dcm_master_address),               //                                        pcie_256_dma_wr_dcm_master.address
		.pcie_256_dma_wr_dcm_master_waitrequest                                  (pcie_256_dma_wr_dcm_master_waitrequest),           //                                                                  .waitrequest
		.pcie_256_dma_wr_dcm_master_byteenable                                   (pcie_256_dma_wr_dcm_master_byteenable),            //                                                                  .byteenable
		.pcie_256_dma_wr_dcm_master_read                                         (pcie_256_dma_wr_dcm_master_read),                  //                                                                  .read
		.pcie_256_dma_wr_dcm_master_readdata                                     (pcie_256_dma_wr_dcm_master_readdata),              //                                                                  .readdata
		.pcie_256_dma_wr_dcm_master_readdatavalid                                (pcie_256_dma_wr_dcm_master_readdatavalid),         //                                                                  .readdatavalid
		.pcie_256_dma_wr_dcm_master_write                                        (pcie_256_dma_wr_dcm_master_write),                 //                                                                  .write
		.pcie_256_dma_wr_dcm_master_writedata                                    (pcie_256_dma_wr_dcm_master_writedata),             //                                                                  .writedata
		.pcie_256_dma_Txs_address                                                (mm_interconnect_3_pcie_256_dma_txs_address),       //                                                  pcie_256_dma_Txs.address
		.pcie_256_dma_Txs_write                                                  (mm_interconnect_3_pcie_256_dma_txs_write),         //                                                                  .write
		.pcie_256_dma_Txs_read                                                   (mm_interconnect_3_pcie_256_dma_txs_read),          //                                                                  .read
		.pcie_256_dma_Txs_readdata                                               (mm_interconnect_3_pcie_256_dma_txs_readdata),      //                                                                  .readdata
		.pcie_256_dma_Txs_writedata                                              (mm_interconnect_3_pcie_256_dma_txs_writedata),     //                                                                  .writedata
		.pcie_256_dma_Txs_byteenable                                             (mm_interconnect_3_pcie_256_dma_txs_byteenable),    //                                                                  .byteenable
		.pcie_256_dma_Txs_readdatavalid                                          (mm_interconnect_3_pcie_256_dma_txs_readdatavalid), //                                                                  .readdatavalid
		.pcie_256_dma_Txs_waitrequest                                            (mm_interconnect_3_pcie_256_dma_txs_waitrequest),   //                                                                  .waitrequest
		.pcie_256_dma_Txs_chipselect                                             (mm_interconnect_3_pcie_256_dma_txs_chipselect)     //                                                                  .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~pcie_256_dma_nreset_status_reset),  // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (mem_if_ddr3a_afi_clk_clk),           //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pcie_256_dma_coreclkout_clk),        //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (mem_if_ddr3b_afi_clk_clk),           //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~pcie_256_dma_nreset_status_reset),      // reset_in0.reset
		.clk            (pcie_256_dma_coreclkout_clk),            //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_005_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
