// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
koMuDDr73Z01h9QNxhqmm4MoHH7c5bci9wx0yufT64nyBwmK8cVCZ7wBFWzKl7iq
CS0zh5HKGAIbpKcRO3gXkzs0JxQqvkniTR/1gye8MwHVnbdxF6jveiaoT3tDtFTO
+m3uJGRkg0npAVTbXsAuTtHfxf2OvSdqilZRE0tn+/8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28800)
8gJU3vY597EFG9kAHFxupYM6c2pkn0pA4UcSEPB2WOWdSN/cT0DyGD085BdKXkcD
GDR2tytwiuOJy5Vbrxzgq0rFqoZyvSjigDLiNkiyCtreL6V1fPSPtheCIxKfCBKH
74uN8wgkNhKv1JOE6lbXAUXy+Obd6D5aB0RmOYCaYTkXkruTSrXTtL+4rCaAAJzh
xDfTMtBU/4CtclLR+G/lKMibzYgx6Q3eHwB9sxcZk7nFjeXETRtL1jC6PaN00kOf
4NnZLaM/0qyidE3bMb+C6meZWobi5Zvd8Zpli9tADPq3iqud6Yv3afneq/8xYtIX
3UBv3isRm52AeJSzag4zHAoB8zigTN709ozVydEOAXRebzus4WTa2euRagFJLOv3
hapvsZpdw61TILXr0ogjIDRNoK8kVj14whNLa0ccelFuT4WySOFadZmsL4vp3H2A
/cGKZS5e7rGiTpQXQ0uEaZPaFaAKw2xuNr9ofu88Ou+WfBa5OofiGUbbJTSF5VWn
HX7gXccBvBBDks1PogmeC3BZsIOwQzjVg7wTzViV+TaH2+zamLiAK80CJ+ksHQfq
qMbNg5L21r3j9CAxh5bWuyK3krqCXBBsY/GWwv5GZla9VlxNKj9T9TH3iRwSl7tG
YC8dzvwetzerkMLZRR9jccamhvs/qc9Am+lQsfLNIrl8SCys4z8LsmMnsQ4qH5rk
hyRJbee8qgGwOtNog1biYXLHCft5IUD6WNAU1qwpeQdmdMmqDA3RkLrtRqaefuhO
G/gJufxAxA2fr7hg9RGgUqLuK+ESuJ01WS6xgcPHsF3Ak6TQ7NHlyuK/BACtEq0h
5rZUY1qcncJyabSyt+TPLvUVFkJgiuAOlMQUlAIQLJMKsPhIp5sdSCrLRmPaiNLk
dmRZTfHmx6P6WiA71BnSmxOQRAzfnv/+2f586TCnVstATTcr4pOW//1OkoXu+GRc
7vTnHyYljyBX/ZEzx0Zc2sNQVL1G/VtK+zYZiKbQQzCccijsLbf5iYyRlsRJHhAZ
ta6KySekIgkkGApCdL/ojeBcBJUeaSohBrvCOTAixOcI1+rhsz0C6K9Fs0HATYUN
RG0n4vEMGCB6KUyQCpiCr1zWDDfgB2DZQ0I2Hm8DvKqHXuUMKNir/KKrSTuJMlke
QHDRdTJsNlYyVUP6tiu9tXQVGU9uF9oDfq4Wgp8zbbelGeBFAMc7/cz3jUkhah4T
uIrcmq+mftolOgD2h5J/yBmiKFJuLfswmkv4Gu0W47s+4Pl9T+KabllISHrxaq7K
mqikVdT9+yE0AiF+T/u2vn+Ne/Mf8VP0n+U7/2L2IcnhKwHWu+bjZdyr/U64ddjG
M5GNz5AxUkxC/3y0M884mqf2ziTq40y2kHGx8dXZ5aJEAKwaxUdfjDIr/AS0ptRt
5r4m/2F7gv85LoQrSbpNsqnJh5wzYlS1jj9B7ft0i7a3bdLhN0tifjDsiZXamWzG
Q9ADWf4L55khu3W1m7OoViaTx2IjmV5RaGTqbHCFxte/vjNFXbE/yp8BKd2F5WnZ
3kl5adKebcTKNieyUhwuhhuS5IXSad6KpxtfbKac7Vfw+tn6YhjVF9Zi5wHgRAu7
zvPx/OCOwPcfjPbc6lWHptHeTm/6Mavx/R8u3/dDAqPu/6jvFD2Su+slruGHzB+r
xBjdxPUm+f9eRxtJ+zxtbRBcEc15SF+e5xXpeeTOFSJjsm+Cz8YScIdvKnilNzct
ihag4d+grjxQl5mqeOBwggs8Z/2FZytl5++F90TWEZ1ALCvko0p1rSBfN3oazGw6
PEu5SYoxgKv5+w/XrVphtn80H/8+Urxb0RSFVax/ciMW7blP6mUPWsPhXgUlpooD
zsI1J1le8A/MKhG0tBgCckGG7GWHGiDutr6g6mu/8wpW8l5JkFK0nleQCykCHSqc
usec2Ur/UegrvCmxEoq4sbfiiFnANF0zVpn2qg3Wkb6PNjqGo88uN2WneXBkNJF2
J0+ZMB1TgT866U7wwc7szsPAENfQl/Bh2JSajTZPrtZInWhKn/kmIETlp3K2HDFP
XdMa0CeTMq7j29ji1y7Dk8a34458wOGAFDaxtSw/iHFUb+EjWaVnM0jQaDBAJDAj
6b5ddnUJ44656q6GKwfaObUIqTIcKe7Jz9Rvkv6y2iBHHCk3uiFeJHFdy068GFW0
jnGEe7w2q10NQOQBHOWwcNe8Vf2R8tdYa2/mpFe8Wx8Wp/8KnIkNE7409kyf+gtv
7cQ+2E9mqvR3L2EBVKjOZLsi/9uIfW2/vFDUoJ+0K6FemO063130mrzMQfnzEbsp
qkV1xAlLjayWRCdWWkRy4sHe6eDqDPuWbEM/7Be24mbBEecD+SoTgjEWK1h20xDi
H1dUgHfN7GRyO9tMefkZeInzlTrhhZ2IPHEhCGDWWHiPwBup5iP5mMlxRVS89jdT
XsNQ3LkiNS3Oi0PJR5LIdo+wY9VbuxKAuZda5iZHG7NhZ5Vp1rfXDFtNwzuxxssu
kqWoI8IRjVegIjU0+Cowd9SCGrS+O0kQIpW+qQeWMtHq1onY7WlGA7BP/s1akZ8i
ZEnaxgadnvuE/V7RvcIyfJOWeNTRcMnQ9J30Czkv1dXHhV3clpQyEUrPlaldMbNg
QPA2w3jrvUNpFyTWYiytw+JwEpeAEGmWf6JcWqYiKpBOXNFkNs9JxT4cSKNm60Tu
0zANpBXSBZbr7BKPrc2BpmyN+6ge4XC+aIAt5Evk8/eG+pUTDgunzJAqSNpJPVuJ
SXFfJUh1N4mRTF9zoAboUgkRpu5xsLB1RC3S+suH7qdjrXgpyGvi+Wn06Tp4lhm1
KHkfNDH9LAAYmXHTvGGOnOrfiE0zotKS6uWglWKxngQrXNCXPKzXLVsTBhWt+i0n
L4Qpk+VIT4r5T270KMmoMHDTbvL3MEkFqnYwGL7iTwYPRGsOYfjJ/vewNbrzs8g7
NtHqYmolAJ99aEltvHWM3eqN3EoOhuln5js3wmqHjCd5Xc0+xMYC7SvIp77Ytcd8
yr6bClngLoJxFrhCBtaghK2XTNHINNABTnYLylW9UgPw4A8atIPX1qQ0As7r1m9Z
H4LPIk0BIPk8fTBvLiTG3UdXFq3k7S8e15EuTSJaadRjmJUNNbuYC7GupUZkOyIG
cRCYHzmPGggrdCmNKx91vJa+UzV6gnbZ4HP4CgdrlMr6P2AOUytL7x154QN2DA5r
FxuxEkaHrlw5YCVrb+FGfCBNXXpcbAs6ycR3T2pu4a2rBwI9aHSAjm46fnMlI7GS
2PgAhbDoKsNQ6KiXfoJ3bw50C1n7z4yiFklezqxuFikOplcQb798XVyZUyg+50Kb
HzDlhf7EASVkatciPOZJeMIlFKZ2aUThiTuHhZB2dGSx9CHrLz3gDG45rQ86behO
wtMG6HJ9tgqCZucje0SvzANAfV8h4BTCcME4EkeGI77Elo09q+4YXSnihG8vLL4K
10N0vVEhZmsML1IzMLSt9sQ1JcFG1M8XrlbIVscHO71Ll9idhH1q2IrqMhkpznis
niU9B0mn+mBWRIySxOAb1Aqi6s9YmChbwZdyVImJk30GXhLlwDBHG0Y3gcwkR+Uy
xixHB1jvRucO759eoDSuS8SchTZcSxhGD+/VDtE6BSXx8pMQ6nCDTcMJ4boqm8oy
W5IAmurCk7K5OJcI4HCzOmn7HRr0sBvq40+Z3FwNunmRY2O58xRC5tAA8+nJGBab
y/zVreSYiDv45jC+5OBZRCN2Yc9zLfYdJzPiZEzI8KN2ySoAdgLAwFkbp2YUxujJ
SwEQ2k/KSgq5az6L3pnWRpxomH6TKjyZjFuLdR7tgP1A7JKh5ltpDBGc+QckvqEO
Z9xEVEbE3JdpPZURng8kQfZ9fPfcfuu1KB9B7wkZRcpXQbMkRwtNmAMjYyRuRUen
iI3C8LdJTByThUHdUTphgTSrDjWX7WU7XTisr4zO1kmjcsgJexK4AtBxYSZxjCnd
R5X6ZiWWfYJ9Kku4lYKR95AkRG7DCgzWkTa9Pr1EXANuuTmqp8x44X83bL6G3/bG
D1y3wlwredcfk7Ch7YbbVpKL3AUCdTecmF/TfvyGK2GvFQeBdN/zNmS+k41AL0ZM
KPspspGFsmFxc1C2Nl3CTDN5+ui0QAGnrBAIxs04FfNpUccNsBhFEplY/N60cpJf
hdh3DUSj9rFU2c6VJxYRNIFK4XWMafg1awefd9duIpsqiysIqoKkPCkeB6jdy7CM
Bf7MuzSMljIVJ1MoZywUoBBp+NkYzNWx9NUHE6TGDuGG06sPBZikqt4alEHFeugt
+KK1vpNpZf5/6lp5dpoVlCLWzjrWoaxrPpdiZA8myjeTZuxe0bIY5TLACzT5EFs7
GbSDHFgx7T608q9SHkLUYHcoHE/Far7MC0FWvjEEz+pHVKV3PUKQ1nX/A320C9Yy
B0Y1wngU1KwhCn4Hi4LsKL94JlGaO78JPnaaBwMb2ViCYmo00vZqvJ5H6qrV3+WD
XkNUFRTQH58qR7aWjTfjIf3z9uaZXXkNyWAVc53UZhIIVhmypaZSyFG2patm7VyI
8YBpICEfVvgNpP0DqYW+Xz3nu16/WepJfNjRrsZM2WhF+XV9zaotltROGAkmHPqN
OphWvDfF7OqceBnFw8BE46SVr7UvLNgGMQsagy0rGRzdV+9Qv6kOH4junsooO2+d
aYHQ5ekHtEZZrux3sQdRkF4ka/AvB+CJrd4/LQLnshpCvgtBV6i27+kUK9+gFDjn
XG7RIYPZmYf5FtXuMbnthhn/xPgqsjYwpqWXdGZ5/1tp6eqE+LcESDCnfR4dybV7
5Ngpv9ni7LXboOLcNX3IdWGEg6H0MJomRQ0o3P4xaZe5Zpa/qH2gSbyIovmlEyh8
XbHYnd6ymoUtbeqM2WMH5r0dq7jblWIJ2Ig7T6btFn0P5thu/KsdvUwAh+cKzXN9
yoDmFQxFwswXLU1AsXrIIarxp51KwLWz/633TL7cqxyCfHWdTjX/LCyRDzgEzC0q
k6GZnHiAP2CjW282EevuHSkdF0w3Nyd9jXw1nPVmGuquMs77PslSVl3agA1TOaaH
B01ti0GS7pH3bWey6hE7axWfAGji5pbz3uyVY8x58cnhB3P84XOzr0EadqfYw7iv
kFhFt+kyXtlQGa6nobfHWNCkChxjNXleVOw6OiF6n3W3m3+accdEgMbsn+UnIDGs
o5srhDk3/qsMuhZR8n9CIfpNBMIVisTzfaPrbngqXkyrEdoQZJ6NG2iBnFyJbTjx
MfsfEQasR46wiWjl3jBGPoc4aDkzPg0njZa8f47N0x7CjqWGbT7fVUWzFt51W5aF
eoheS2SgMFyGUiskSpgvs2kCM/UTc26mf2c5c6mtt7ep4rAsb84P5yCluiegN/SB
8xSZsJQ5x0F6nUvD9Dv0E8DBe6ARGvHRY3aMxNtZ8LsQwmXyqNGATRbMt4hIpN2M
GHUOPOVFtivYh2tp+4xbmNDXaEVDai2xKkhDWcQnSGWfgsjHrNEsKLaoTCW6T1Gn
7EQFyrDuaBQ23LJFpQ11espq+Lu/GWw6FKDZKr/KbHt48OhghrAB62CJSojjuKqI
r8B2thPhYtExQIm3i/8z7wcq0WrgzhgjyU63mKk8YCNTct/pUoHb3mSiD/o17n9v
MndLY+FUBMpiW/YZKuaGQW59Xj7yG+Gch1qLO7Zurn2iaIVGPW1tPGGV1uRnoAHx
TM773X8p8Oqq3fcL1BtDpXNXRAaRjNO2EQ3kW9GkPI2JD3jzQWU4I+1tjUE/1asE
kRjyfG0nHKPAQwCVYnYUN08z65DLh9JJEX6UWi8J/mdE+irmOmVcS1U8I2rakW6D
pmhCvIc8DXSoFFGS37v0FV6OSVqfKTQBThUf8pXjRvHlZVCl5msbNCKBAiPjAwOR
C10TwPSXufrPX1g1l4xi/pwaW/e6C6TPNC2V7Fk0xx3HjEFS4OJNS5u12Ql20FqD
XXynefK4rolN5Uk0r12JhEQNeXu4ycoNrnniYQBnExf2uuUTVtY8SFsqsX5lLggw
dqTLV6hVsD8LcCz9ldyEx2F49LWHr09QAdUgPx4AoT24WEyUe1uVjILFygrLAP7a
sjEjWRVaWpNbQAA/9vAFwifQ/8wWphPPvnoT2kBBxOvCUB0eZCs0m5WgwD8Bgm0n
SGfXR5mfFMxgr7EwedVUEUk/HMkG2rGn58EtgLaqo8Dxd3uzWK4FjXZGaeBfwOO+
HwdXNiB0IVTM4BEd1tozWWcUQi61olfyB5YYvIq+vu3PtwuBoxElIKSa0qB3slBq
r0FqQL9V3SVftFQwCuMyx8v5YlYRlfxjHTFsl1tI6vwyLebcrhQxRsxtebTw1yFQ
tMkS8rfohY70sD+CmNq4LpqO84drZ/JOet2Wz3L4H0YcxPUpLbmDLBp9VINzgCN2
ljt1DdtC+hYq75lDnQHWJ52Z6WHNIpbzAUkU7L3kLD1SlVGhIcAb0erQjXcPIkvM
uD1jMmoG/c64td05wzUi+AbSA47MRD0fB4368v6NAQw9HjulL19tNrRU5Q4o2q58
E2XrvVXvgldIGziQqF7gf0d4NWn2PAAngrLzb6m743heRw142H8uWsh6Wsl9JYk7
qJkly/QVg0XSpRG8r2/8qb9ZOsEij96f4mk3KsAbYaYyCYo52tbGdKsCuKmSjQop
lQRLdHZKDpVUbhfjjHD6vsWYtQUQyctW38Rkj+MTwqJEnSxzCH+wwC5Hmz/oBPEt
u9oS4cnrNvdS93SY5WtcLmn2Y6t5N+PU1SAZ5nbpRqed65g5MfkoxcNIdbvTm3u9
F55w+rdiBShdtORcHm6B2/z2dBQVT3AGEdlqyl2qVpRJpzwU58Fjcml88JPu+mNW
cQigjD9exVXHFBs2pHZlgo5a+NwFOS8Ab0g5cfbb6Am5BWzaoPUYUXE8goDmYsTK
eT2l/O13xHgei6xxCOcqP475EmY9BS8u+XWm5Dzw7wZfyhKWfky71t1br/QCuUA0
PIXnSA/KKo+22NeBquucrFgptiQDozT6e6IkalGUw2qIdYHHiCKVcPnQ7D8uZdVM
qHrTSvQwUJ0jPMWcWQ4tR9FWM4R6GUWE8h5XFhvIvCAoE4kQdHDUqd+6HxCmJHQP
YNmGnudc5m28wfS8upx11KXzciZYyzpx0C1ck5Cq6EGFunU7n4YrVebY1j1RgPdo
sWRiCPsaYSDeF32zvjcbxAM25Fx9COsvoFpOxT+SfThJpDD6FnqB0RETyDFE68dN
gUNQb3fWA0V2Xs9H/i73dWiXyUl/ByA4ioDh8359ejAwLaA5/j416Mz0vr42235k
NfVIur55FLJQBR2oSiPsVDbPhCj0XHbpURqFssLWDa3M+aSIv/aPhzyFtxBwli4p
UoEfI0VXBzC4u2qUpguURFEIBQ0jdpUDMhunvryYhiJ2fzycrOdKbYIBvISqTuCV
dp2dhDdwT3wiJ/7nbJkZYhX5hpy5gycyNvzQOkhwcddCkg/NgQWSc6R6J2QngwY/
EUvuQBQE+cDZfHZjSCsGR08Hr7pi90ZzwBuwfmmBAZvOAk+rdRrKCWAiR9RW9t7R
2PYdlYBqL1EKCtALzjhn8oCm+yWeX1c6SU6Qmi1sQ6K0DuH+Ve3qC7I2HHH6VfPu
anZX0xg6JTX0/WGR6XRYc3h4OrA8mCsicnqiQLlUgLYyej0qdJKNvxNzDUI5VjOt
vuwb7/gLyVOF4bLdpOKoaHjn8zEZV5OmeZRXeb/pTAahUkrdmX5XlU829SpD+Vxv
BpnSRdLS1CVgCb7jnFHHB8fmOhK9lry7PSi+NMmHqsJK1P5OezkuQWVMBvbB7u6n
CyAxoIATQ0U1dGlOOr592BzqUcq6UU7k9a9jE9nxqSj2deJEoKQdj4oICzFPOHLU
e+LguTIWItcWD/49sxMPF8tl6spBcM2NMTdN6ijOk48AvBF2qHTeHcFldy5Gkp1o
ZEfKHggWgneOkr9eRxwHmXMgYppwY2vANyGA2JKaddRZ0X/CoUYyxdOGwN/KtcQ0
suHvHG5CSjGzy8iYeYYy644PLrHXs8lew/u64Tu/QG/ehBVMjCyXUbrgFBtpTy91
UeIf/lsRdvQ4TJ3rfEKUCVZZq+s6WbOSgWvCCXQfehTQNOt1azbSMjT7rPgSP5Zv
T3qYlPLmIsrVfxm5o8JH9hmPRDUG96j6THnfavekzPRkYmRTlKim0Gy65mMaZ2wZ
6OYPNxr4b6NUI28XT49IM7eC+vTfCDVMPQva0HHmNSk5AfBCXpmWuFGJMMhmDa6N
a/MfEQ07m5S+8TrInBDZSlpkRgKYh4AWYoJNpTXECgpl6sI4ku6Z12nSXytaX2LN
wKCZb5e1ExV7u+becj2IUrnCrDvPqwNn03FE15r/1HEX1JZ5ueAUHyaUOB9AJ1pU
j7DEqZQR1AK+PFQ32Ngw+UxqCvBySMzQ6Lpow1/9XVh+s3qD7k+5L8KUHFL7V6ap
goY1nZnGxDxRvO5mdWf1JnyHnjnXVNi9JMuNM5T+qKTgV40r3bcwIMcjGalzfWKx
zV1pFSBHnjT3/Q/OzjcIru186HbETg6WF/5OHW+txEHcG6NrczhGXxdvd/VNLIxS
J4uBlXC9W5BzsJRAq/nOuOftgiRcfcKKGH7NWvo1yHZUaiQdv4P4Gs1gbJt33vbp
MrYXDPw3tUQpPkzs/coLD4YyMoet+KPMgoYZynjhT7lAD3KlqV6djeBadr6HXK1F
45tWvrKlY939qXr9ks1bn94nmVK4QsX7mpmlpvG23rXihU9sXk6USj8XrMtfSKlC
kFDqDYQrat6PFXnYJJ6LiiccaHFh2jKJRLte7vS5l8Vp7zVFElf9lmRjRDa9VQgC
upwovfE716lB++pVt3bM4nK86MKj7Vksp4vPSFFlF6sS3hjLqml6xYTodCSfvTkT
YNT7KDfRV+N+5CafCP3aBftxTEGzh/dO1xeZz4O/oWUZX73NA+iDNb8lAUgi/B7g
HWi1LXfg05kuLFrl9V9/1HF7RcaHjkzVfWzngWyvGgP0HzRyH1v41Gxhdm/dSmqm
4XTmwoZCioC9/MA29+ZYRE3s2DLRndn1+pcA+ypJS/8BfLv/vhqkNXjA0xjWtxSe
e1xDuI5FI90VN8yVp2EqIvh9XU94MpYHnOP43KrzGfjuQrz6MfDn3xSe3iTHLdum
8Qxg1j07DCP7y3fCrkwZCh6ANYOIAZV3sD3x87jOvs/X8WE1NtIXT0Mee2QQaCko
ANlW99BSt+vx51gK1irhlbdFQ6sLKJAZB9BAtxOfhsL0t/1WftvTXh20ZHyrBCvK
e3kZuULc9Nq7momBAr9cK+OoKfEaGd5juW+J5DixyoJ8Cj31n70PWng6SEZQR0w9
wmyUE3rVxL66KrVx0UDlkSqtuwj3Fe7Q3sA/mTqATpRW+mVIjm1J/kRr7YHys/bZ
bqs3e2U8BGZFOK+ahl0dr7V8qov+DZDjMyfhc6i6+LrvowqAlALk12fSjjxoIYVy
Uoktvbxb7LEp6esHH8gZynIVfPMv28sffhojiUVWcXDfogKH1a/9axKaMeD4gvWQ
AkwjGuvQ571F1+KRnMIQFbYfu7vU7Qmas2RIFqKaVQGeK918l0Wnk5QAXMPYwkbf
qXgJSBPfxn36ZyKaQYodBGorP0m2FvDcx5EnHaZx4ocbYYvLguwPlbXFko1Airjv
xDGs4JcjZNtJyjuie+LiLtJSLYuEfk5pA9wNQOqyRosYHD4a7AosrKt9LrCcVMf8
ItiSlOP+aAFR/bXGCLPsjyGNfsZzxeaC17CXkGGq1CtIikXA+f5Qz8FEaIwyU87B
wKVstlkJFeAWwjbv2TBYNlU3wAGr3dmAk4p+XwO2MBZtYO4DdiqwH3aeZ7T9izj7
hgo7jIoF/8EOUImxYtObA/Tl1IMAdBjdVil1NmJ+EvTQYBrLFFKpKjdXZICQJdrV
EVhvSVZVUIJzlOrXnYRtqNO8nHA7ki6i4d+zxTR6ecLvqNbUCMLxe1oQhyZh7PDR
3IO7rkbtZj5yvtUOZBLCVCN7fp5bC2DqFeptrvS7VW+XVOo37H7XrL04rRM2A2vw
vPN8xOL+lFLc2dcic0fkIKw3Ts/uKfyx1aYaWqr13usiMJGNlCFTnpapXvKv/2db
oCOlFvYUsJqmSnnkq22W0WetLtjRoyqR0VxUSqF+cXWDnzDUvjGhepZRAy0cfhy4
hf3TecciuXFWVDIOiCEMLZSTLfCaxmn3xmTLe32lqsFEYCczjDepbQGdzrClVLJd
zPhaqLPGJi5KKAMEmPY3L5Ra+xX5xJyOtrfvCHRaaShvnA1tLbYAIzQJBAl47TGG
/Vl5bKK5+0i0rm/cBzawvIcIlJXLC7ur+A3fNWwUar1UdZrVGG8RYGnKt+mwMSGW
YmoSTrAUOHRIQuslQRI5hWDNMy4mAkDhEYtI095vGIw5tUBUmCw6MmSay/cPjqRq
BHyAKsBWeNMsGcvmpSCm3YGXSPJaz0pfF5BvKQ+XlMTTK0MVEsdHPjsABDfn/DwW
HCzZUnzWojWZkHltNqukCH7YOoucAX0jWoK+rla6UkGKO9nK29ovLfZ9+0/Tf9x4
6Rxrnp1PromvBn24xbMEk5OGenjTy/5Pogz/TEqXnbuI7IsZf5BCO6+iCQ21uwYg
CwpQQxOxR1nEcrQ8ouZ5VnGqn7yLaSKPwYKSLyaYhRNT/7acCnVYylSCbqewCEgh
586EOCpIgKRGLhu1W01oRmCcHf+n5Mg1Yj2BPhU6S9yKyppWUuLEwKzt7DsiHzI+
YRUAvJML7aTFc6uWFg71xV/s9dA8nqdFI2wRbzyP0sjpj9kznaXhpEHDPCfQ7ynQ
UBCKbli4MhNtS8HGAR2+O4O/5ZEf8WkablVAWg1K/5v7n32WBD3nsFvADpxuu3/B
rLCjfrcB7pb0jNB4U59bq498xJgCwGD2fpFxTOzcl6S+/aRvDGB2rT51ueLlTqfT
JJKIoRu5igiOHsPXrtSQsw4/aCPPePlllW+Upy/q0C0texbyJx0pZimxx6oXaOWQ
MDk9M1CrmWNwIAXrjiiDhnl+/70AKZKyvJe3B8fQEz3G/5NGesunUbiGI2OA9s6z
FvjthJFln8uSH0sWXfIlMqlrQk3ptCmL3J8zOlWijhCqF+7SZYQl07aOOqxDCkgc
n9e74m/k5w84BaPhd27RkQz+SS1qfc2Q/xsBPRnw8pzKJtJQkNWhvY3WjJHLUiQh
+AIRAB9vmsSPR9ENAJcW14Zzmwjx3jq+q69XPQ24w0hnQFfT0BDhPaiKTQw1IzD4
6rZjTSRo72S+bwnIGc71zmFeD8YLqhUIfeGQIKr5bP1+9Oa+LE7bbSvHvDe7659U
U+N27R1czP4Of5JOwd0vj6xdaS9F7ZJFZs6ahj7at42ZZ9lsv+mduj8rkPeJAWRe
9GM/mZL+IV8LfYzNKjBxPkZfFuGI1lN+4oWT12IQ8xHvrV9CxSzsxeLgyjjHUJeZ
KWRVK30oZfxV5JjYq/kdsiqU+1n7LkAtvSEAUSqxFmHFs1OdjGOpjAALMxdN11Zx
jlA2r9BY3T/hPLBteKnfI002Dv1J8SBQSea2b1/XnFalH2lcsfSetSb9MT5F/S5h
i1pszp/Qw9okbEufu4s7CKyYa97xT+TATjhsSo59XkIs1pZGtnB79gJ6r3B89uFn
1XqT1c+/0CYiuiVykUY6SgsHWG0CgbpCxAsDE8jJEAxWNL8wQRph2VwmvjjFUKNw
VvMk4/zckdGkGiaMwYI9tUwwIHaIm8MrW2b+LOAnjZl3EqfoZ0LxmUcoz9rByRzm
3KLhF/1esSSTWdfDPruNrrDTvLs8373NpY/fTbATvBQOHQ/+/2Nm3cqCqbedTkdg
yBVMxT44RKngQksLVJvzOZQHgA+DK+dRct+76WfY9hK+IVaiH/RenAj2PVdJuZxG
fspAc9yhGXVluc5lZw5F4Vlo4mNxXYEORgKcj0Q/tdup1QCX/9Hju+21/CIgqgqZ
NnnWYN0I68YD2gEVWfSeGmSCwN8zldT1ifd7JvarEaJxkPZ1MSICZzrfuDrZAi5g
4BDpJykvmiuETBVXw3SdKrHUzzeS1HUVGW+9H898JQo0SP1i59Zt270WAdfCtPYR
QbAUZYEIqZ8DvPgq0PlfmpPrTWtpeOfoOYX9dX+d4nhUzEiyu6oDfkiB2BkoN6eM
G5VLlp6Sr0JyLBuDkTSffQ6dNffp2cEYb1/T1qNlY7OAYTnW+coVlteMtklLEiEg
6QEHjvNmkx+czIuCJHwG7zEC22evNp04d3KOcZRFo/BZSE6K7te5J5MEkymFeAqy
eT/GAmkVYI2H4rmhjxBWeBUTTCOpc2XElD2kDH012BLJKf2vQMvLZmfb8S1XN044
ieQcEL8G1d1/nTqZkh9oswBpJ7KXLSfZJ+mTlCVRQm36+kvQ0QRh+JF/VJfNgQ4C
RNBXKOTpxB3JLE5P4T6zv3BwiEp9mKagj62RLGUtPoEi34+YxhAcq1IfWuFrQBvQ
+GwQdg6KcuFU+/AjHU31XYYEOxrdr2L/NCeA8eRwyiSlaxZsNq4xjrzcljL9eWrL
x0OHLee0IjTvwRgTSTtHnSsfoa0i2yUfbOXLuV521frTel+xNoZ8VMDmrclMRXDm
y2LfoGnI8xDzBkuF5+ZxrqpUX9FsRyKKAVJZARTtplZuvAZQxQHQSpFUzjNtcqmx
A8m4/CS9Tjf85oUbCdZPqo4xXS9EdovXDVydLqG54uQuiMm3fTv+DN4tVKmPT8dx
HR341as5SZBwDxKJBO8hbKiW2BwkXK9xlu59QhCiyTTt7XeRgOtWxnOI9zD4MS7C
DnMJF1UOXKuF2b3xTwdwSL7l02ldd/X+ddDCI1OOxDPSd3UKMB2JVRdo0na1XlJS
7kD+ytbQARPSZa3yo2fd9aseHOYWEDGLYkOfspHxhoxtM7ZHoVGY7nU8S+IgxQNT
Mjr/oU5MCeHU368wbZE4pWVBG5IbngFRCZ1BHyBfZi0A+5PLA7WYprpAEKnMyOPz
i/Zz0hYuOzE/mpcAlwhGktVyJIK2GW5aNzi+Rs0w2cbwcanl48QLIUd7UPV604BY
nPXet+/mfITrcf4zgwwbDly93XVMYxgaBH88MF5//eBNlofSrY61akpHNUVDkp2j
zYLYffJxryGtK++aC7es6mCu+qkmBLlFRDp22+RILgBYxd9XKixkPVooGkoNQ71H
20FUV7eUfiNkCAzk3q4USgeEeJSjLRfhSIjHM+9pkjOS/q2TOaUl6C+yTjfAAxs1
4FVeeM/F1EN5h4Fxw7YEc9hmahgoV3lal4qKAoVXQgTlN6rUQWSNhQmBItjRramJ
/jMw9Oyb+wM9ngq8P+geiBBVSWPdlZJ25JiXOEZronY5wL01vu62/CLD2W6mKwXV
bfwrI6IPI6c1+R05X2KtdTXt8zKNJxhPDfTfPREdTnqPNRo6eoOkLZk9VFGuZfUt
r1gBccM7+Bj+kbZxx1wX5veU3C1zmokj3+YDtRxZHF5bNhwnaYtBaAyDpBfPd+a5
9GeC4Vs3c3GWw9hpF7rB3E182Q0Lal29PUry3lmhTm58F05cnTLEhrMoRMTkPC+L
21K30eLty/CPFrf30rCvTvPA4O4tGFdLd1CJphfY6YLfJxHnrpFwXkIrT9RYHDoq
xRSWweyL14hiiRV+ALPjCcgarvHGcXrQWCW7rrY5XhDea/sRudcgm1kPTdfPGrsP
EPcuqZ6h4rOrEV8mfILHWLW4WBhl99Z/dc4LApn0BymEEyVWsTSvxZUns7UGx68W
U5rKGj04BQFgd3AD5uSH+LUrZ7Q6NCBo3osjhK9ZDpCAGQAjYhu+53j2gWpN2V5N
DsMYZzrGkwjXfttJYA9o6t0MiVGhS/xkFMM0GBGMIdaCklLqfjVgJSxHy4/KS7e0
c1jisl/jE9ukBvCj6gw5i8/XH831ys88mKHO4UoKuuwwjixmPdyZajVepRHAYiti
YtUDGb2wE73IGh9yZ4Hc5oHD+Hkrc+uPy5TYM5okIBTbdhpUzrXUKhuHfNNCdepO
Mxc30tEvC9P8gpgP3JzRbGz/0C8QUzV+cj2Ab39XcVVPWDKa7O6wBjtzaAtA7ACG
sg3Vjdzc1HXGNfbnMd43QhxT+/Hi45Wl+7vFoV3HU0fPtuJuqEibEwQEMhfYn4aj
6yHv2aNC86tebLCg5JljhdEZXA4j919AkDuLl2zA4C2LvL8hvoLghC/AEa70OKqo
9y/6+aRDPoplxD1yiZesJGKEWR0hG8tatU445JqRudAOWmR4vJUSxkED2cWEKCZ0
bOV63FxOp3KGu6R9/2YiAQu5K4/1CvIpm4ce2XQc0bK49gL7IACtoRdcgDSt0lcX
G1kJ1OFHh5j7Kh2svUcy7Ftg29xunQQU/kdT24xhlOUXg9ezYhNI+3D1tSjbCmYR
z+z2y7ojgw5kZptH8/CNNsZvOfqGt4nSAc9ICkINwO8QGAZipKl8KSrB3lMwVHsN
FefCMUgXb88GoMOMOAF2RMIEM66nd+EfiM6FeY9DZySUzjSdCgVJP3IcucgT3MwJ
bKW3NkboTh7NRiAEjUFQV3YIYikJdT5GQgNMHLj+umD2CGoPwPIhNWsA2I3+tF/T
nCo2AetZptglS3IB31LwTS+mlfFPivfBP77rnvwBYXnaW8zMb1qs+Iw9An4Egf5w
pNyKIMzQpAUWD2AXmIGnAWKd1VccjiI+JPSaxcwGnjluUCfxMVbzP3LIgGWhAiwl
aDBi0Jt7Y3nm//FdttP9uHjyN551IA69Uun9aLwH2LiXEIs/KT1roElavhxITh2G
HXHq2/S+4Z1zMn5zeSmy/+NyVTWvs8LMjI4gK3z4aTXpinI3bP1IFRqn0xVjDAcD
L0faiW2Wuw18a5cCPWPqS5y/yLyGweWLhMbIcx/9hsEz+jXFOCmG3Emb1TvWUvvm
IHBTe3zC3X7ZAMsSAUcgkkdc+WRsqosI4uGJNQMGmbY8JG0T7iMQk1IyBxH7hU2O
uixVQ5gm0TaHA7mAO8QwSug5SvVEJKdWyj0dkP8IcHor8LYcgNcDx8e8CxeuPCbv
k5K/rd6b4Lejp3b30OZAcqePv7sap3MEgRbv55tB8rRyBz1dBjx8eIcY4RlSY3Vg
WClfPkCBFZ8adhMW1D6z2qSfb2tqQcchzSRcuG8e53/NJ6PMCpr4jnno4tSiDGFl
3ptQq33GxyVqPvBNfme9Pib357k6lq2MUqjh/494LTMpqRl0UkBoiMLPjDhiHo//
HtY4KH0MKtgv6Wg+XmfXI/5X/wEG2aHcz288LmOwh8F1gS5D8TKH3U6h9ffapDjM
LEyFeKo3vScqzSfgxwYtObwhnR1a9dyV6Z6q1iO/kIPKlAYIXrAKBHahBAxblO5j
rRwpZGlJrqywHHZsOxcJ3mHtm3xA/RM5NFqcsC/2Sr7l3eSzF/51HhaTr9wOwEPX
X0vzqlkKwXTy3epL6t4z4u5FZr2+2rvIlD0naG9XfMv979iX0rp1kw2ZvusjMH/X
J0lqRa4nkreSctkm9ssU3lX29XlQifkMFF31fHWbHWwvJRiKo6Ru2yd9uZMg7RLR
KsOHseJKiaahAWMfc4Q+PJ769jOG2DDx9R03xMYAIkuo9qeEbt6a4XZYxzaEiLVC
j+qniILW8JI8rXaIzNmV4q39Aobej/xpsMHYNdSN0LXQArQ/h6zP1gDG4XkZOm3+
vVCA7hl0Jo06twJR3NN/2lNuO8EHZq+4oI6HsYVs0XZ35TkOs1C62TSeiPRo6H7k
4jdckK19n2H/Wxzhq0pSBkR4ozagRtWuRxIXnSNCc8k2SNDhOPjN11f7t1aOq2GY
OdGqvHy7bbWwgEj52PQwA+Da1FoNU24PsWKOrvSGRk5X9ey38CHJXnhjy6N1C2df
4G44smb42fhEe5kUWSZbWetH0ly1c24WVGbwiuEFY4BnGQgrFN6HW4TLvQLTJ09H
bQtUAoLbMDdeQtEnHm068fvI7cAD0FRkYp9B4DARoonEtC/AKOvSeMT/tKdylZf5
woNJCiLDJtGhwvoFtD3gbGVB2N4ewyJ0lIf7MwfLAR1jJmIGLceaQbd9QBOqT/YF
F4tynbxkBmwdkbC1n711SLbpzcST1mKQj0nOtOt3edKd70gPAj7eJjnNGHrf3tJ7
59oe2Fe1QC7ZBsrJ7qVjGYvccKvUfXejizgjvVWb3hyNg6dOxmu/uasMpcCEz4ki
TggoJuTS211mxr+EsLZaJiskcXgWi/P73iWe5hKLq7g89JTsE26xVnNpvlMJLcC/
FMDtqmj0fqdPDx8OcdNbpJAqq6AhgFXRRjlFZvd2jmyFFpaynlrQQX0agaCcACnS
fPUGdQoOr+xTtF4lJ0huDtxOyESrOIbwz1AVD3n9yD1ykLtwmuJ+cyewVuAE26px
Xj+xYNTBpIumsmrGtV2fQx+JBQHz+KdoAPgXGYSoHg+shU/rpTNRc1wbI0Q2Ioq4
LFkLHW5FT+5YKci9o+uqUXVSRO6tkz1Mx+zcFKpOjl8/lBIYlLGQtACZS1l8df4A
ujpp2REGTXZXM+TXz9xe73DcwSW5ozeJ5ZG+tRCQPyxWIgmvQ/sRJbc90uJEY3Lb
wxrgDZZVXloTAwLBwQBLRtWbtByhs8nc6Y+rFMozfhYisWpFCvB/N1K2sxXtrXgA
SaJOviwSyEPQbyQdfLLwwKI6bvZMwtrcMhb60h/8gPc5JegqIImWL8M49SryLbfS
c4IU2TgLRwKOb2EMblj2tZZbtgr+kfqEHuY+2/mujOYl4bebM+Id8q36J8HKYRp5
qY+IO3WJkneTI4DfpFY7yz/NR877m+LevSzqho7w/D9EChl/qde8QMfDGnQCiIVk
ROTgw0MnZ+ZlmhZcwqTfB+b8qxuKPZYaK5QeHwU+AMiRMu1f39TyZYcBVmLDOg5k
0JY9flo0V0Z1PuwWdQV0fYSIekL8W3SmY0190Ds6DcoyuYfUqE6OWTw8ijKm+EGr
gzOiDkq0z/2HMSdBbB/qa7Na2+Ibm2WrqGRVFdMfPSCdSn7TtAyv3X68xiDywq8v
qJy4Fk3fu5NomHIGZ7YUtLc3SL24M+avLdQoWdqTYwcwy6psBY1BNOeQci49jwjU
PMG/5YRDBIg9gxyryY1pr/K+vlvu06k/3Fp6FlkIGlnQK3DNoiO1oCBMD723Grhh
NRVAcm7ria6tJ7Yg2P1dkemYprjyugsfQAaNzWMSWboOmaNOMQ0jnIXgy+Myiuz7
JPljtBLRx10pX58XdBJyMWF8noU+yBi5W2r3uAf3GkqfCOLg/E3p7CK8k8l/14q/
3hYtq3znWER6Lun3qXOoFCRIxcDqUXDNaI23gg6ohaNBKf/7FESOBI3iUEhwXQZI
3eXEP9VLry4+MhliooJ+wZPVmJ2D/WjzlkEiNn8WBLQ8vV57J4lbYA48UEbOv4v5
Jk8Vw63MFYHLp0I63Jiku0CrEm9T5+pfPIeXeq96XYGcjHYFQ18NsWWPD7wuywoa
IpwjTmpGrQK+JGaYQo4Tv96ZFNL486tx0uMd0thcvnXp3FEXWRLNIlsIGeDkLi6/
bIg2/5G2RHCJRygq+RX24GMs1DW7KNVgSleSueA1GAn6eADX8xnT38K85fpjaoyt
yzVVC34DK4p7wSj5bN7L6bmuLgby37Iou6A3j7oTW00CQAusKf+M0zMtDusACpvZ
s3HX2lUEA63HfomHg8GukTwBX42vmCwZxtJRmcJCrqphr0SWDWh8bkPEDSxf9gCa
RORZ+6zftJD5ran1sW5mOcoME74eO8POEbwwiMHMoudb/Vi72E5KLxXODENhktJk
r6Qj2EhhYx77RYp/8PYXiQpuiQers2rjPCk9BKu3+vKkHyC2AMmrdIoltua2DWSe
UxFbTKJZnbTJyE99YoT6LxBiMr8i7rXUEcHzwYmDx2hJiAvyAXTXYj/ijedcicuN
b8WezUCGunrJ2XKrKQw4CBBQjWe0flcFhhdsWHwEwtYm7RA6U2fnaJ+5k54UckbP
7mEZR035/UD0w08JoEg6aB04aNCbSpJjA30++7i9yMPRnY51Ir+RRm4pnyFRtKk+
5CxehF7whdzO992K8snJe8fTsXKptlWQg86jP4nFIHk3SbPypyTHxIo39Bdn/Rbu
wOnOWCG5S+wy6O6UJn0/vHJDQ65fvSIm26Fe9NqVe0+VTQryqLpnJ1K297tUDsn5
xj7UiEphiBJn0tuM5kuu7nAq9Yex7rtIGCXZxuzzTlLjDKAhtUdf+f46YMnKmC9F
+rJjjVHs7R0wwT0bDmpLxl80b5ug9vYV8PL8koENT6ff3+tJjt0YIIZtQv7WgDdL
BqeAyuoYeMDY8PirIjSfinVJT7UPCOM/mx+NZdbV76VybtqlRIFhzO1dMX0hjPFS
P45w7kccdMo6VB6E8WxYDXMM8FFtCz6OX5pnU8KVzpzXQob6reiqH1b+HLRakc5O
50O1DxmB+cbDwQFcz/CboUv0wNlvnBYE2x5mRUJKBfSICBwndTghm3u4QGzyj2cR
GTniKITpsTHYFPOUSQJix+sSzfYbOohNugPbrT0IVIy4xxN4h7iFm8K+O0cqlhJW
BeCrEmUnOVZ2mAu19FOdFcLkX0P56BXKnlw2NZ+Um83++O1gUhk/VeUo+yiKCVMq
p1LkPgxRRkBYOSq6VZDThgSiFpfXfecrVcVXXj+q3vo3Ebea8ILMXWLFnY0WU/Kr
kcqSlWMYkHxHxuEETJncqigRvXoTvh8+lGiU63dKLLD6n6+k1+Jx4wznJeFbNSXD
yyo9+PSgFOPHO88r0gvKCIRacPStEo08Rs/UuCBYMIttZmcWx/oHNrup2exjW2K7
PYkqCtK/p7g42l/7FdNdB/G5y2KthaA6r8WWNo2+BDfIBW/2AESxRatVG+xhLClR
AXt9YsBgIWMqFGIxOPjQ27cqVgmNi81vRC96CiWZZtiBRnPC12d5ldPQeHzEM2Zl
eWykOvhVG0iONjAaZcQG/G5gsp15QYnynDwiYLF1Jiw7pAd9Lus6I2uaeVv+xeZo
qA3+R8UNXr8xyBqcwSguBZSk5NEKlAWRzAbL+mrdwpDEeeiDnZJVoJ8TN/KWlvu/
2hZji4GvKmFsOPbkEIdDVGzTMlGubFTVwCrUUgjw850PFKWyst3Xfnd4J6qkx60Z
i9qeL0TSf6PDjq+Uy71uxNw0S/mGAxgJL0Rrd0YscbYTQZhQyyfncyUlEyEUvtjO
JlZ+BboMLKxTS7x84iHr+g8hh2DDkL/lM6PfYCaf2LUWjr1Ss66cNXhNVo9JC3y3
deLZBZxvVje4dG2CMoMtSdaJLQZP3uTVIoL0B1ZFIrxCi5u0gePVp2C9ey/OQjwk
3nSfzYE+vFPHeivqTkNtsex7pnbGarhVFCsTaTycnSUOMMBaeBSnj9zDCjrBx41M
zjf/ee9aG2XwNt62BQor87LvzxDaJkp6xjOhTRtpCX5DEKN3TZfmlhZ/yCEkcLTi
8xJTyeVVBm7r9nMXPMeNvFT5vMxQ3W6vQ4LPJrUS6Rqm6XYvpilofzSEseztm5au
O0a7Xhqglwbgbrf3VE3O4cb9/ymu0WlDthl14Nj3FRZD2ch0L01338pTUGMnW2xd
IsIJtTs8TypBVrvyH8uVs1FxWhytqQH8mkgr5aWqjAWaQXPvV/2+zHamQI2qUoIb
e3oONSlXJE8bNVfugCmRWwA9cG1P19lVq40mxVV94hpGTTiWBqlw4srqX9vfs+Ux
sZkrXuISxGhKjPXJYqTku07p6kd8JaxhoHf8uo/Ao078/IMc+yECGh0R5ODFTatm
3UEab01FkQsjp4OBSYN4PCj3YfYUM9H67Mpd7I3FgbCjw4LV3ZVthrVaxCevOFgd
00dXz07EkygeB6pa8p0URC8kIyoa/MuR12opUGY2mAd+Z+v4OOHWhY1cNb6iSKT7
T8kQgmH5irb7tIowgmWS6tMSdzW7WiN0sHtnQjoB3rwgOAxGnbKGhiMa/rXFBGyQ
HvPxKbb18p7E0fyXA1F6v5P/iUkG8sO20kLShzBsPCdiRFqQB0YR+dMzhZ3JOMhx
BNQKhCcSL4JEQLciKzhdgdt7h7xry8d1Gf6p3BCYDF3ba/bWXOS558dYF4C58mJl
bFlwT7FSjIDtROwyJcIHaHiYHtPB7F7ps9BYUyS4LiNoMY35cGNuI9fus9/aWHLK
eQitkNJak1Mh6PpLRyongJWpx+t/7xQP+eUDDDp0NuuJammdxlUWYJt2dgoNHxlf
9+4JAFMCl3YgFAxPIW9Tqy0lDYUrmh/CGA+6nEsLTChxIltBpsJF//hypNS72WNY
m57PgrlH7ubHTgKJAFgGGWOAu+lWSaHHn+ZZfKYRlTF81EsWo9gdgCWUFVywQwGO
8ZDWH/Wnup2zMoOEUF1dfdu2n5pUU41YoOU83riUAuxRGFZQgn17HI20bNrn84ty
/tckyc1IpplaK7eSv+QDBGJQfABC1uLB1If+gsIr3/G7l6rjIgvzLo3AJZL8dOgD
5E68j/y3KhwuJoSOhleE0dkcM+dfK04An/PA7L0TcgxMM2R4VFdrnbwF3CqILHCZ
gj3QfUFdihS8cBVHKJGLoB16bM4wH+UQrTCao9nHXGHGmk3xcwTtGIW+lfAu1L0J
Ug71kJOXw2gLfn9j2SQhEprOC+xBoAD4rQ+y8xTwngcNJCNySTsafLSZf1LwJnEZ
rTiM+FDejuuw2Yk3bGTrR8Jbstzikgb4DwExP6pWYh3ZuzwiAH2L3R5ckwmSGZQm
tstwCkg6zjlIKF3lYFv9r4zY4OIMUiBmC/KjD4411zR7f8v6dIthQGg2VyFlBuPK
x5SpspZtnD8wwLrUPsf71sDuFGk5lF4Ey1gVCD2HeHXiHkrufgxc+9axcsOUO+pS
D4VFgQ+lcbypcDxwZ6+mCA7JS2AoKv0TpuaSgE6clijq6H0+HmxJzzKkaIZZcxao
x6qHM68e+uHVJytR0/m2Pflw5rNp32R4hWxatuZu7V35XivdmugNFQM5RegOJVDX
IQO5z3p6WFz8GIpCt+M4n1SnD3juBG68DEC2TfYzeWJcV3m/7taRw7aH1M7BWdxx
BYFCnd+1UKgjevox6DhdN5aUpKLzU8pwmjPv5q2gZNCtI18yCgd51FnxjWiS1UKo
/KdKWWxI084yfLb+ro+UPdU2C+sq8KRtP80cQJGP8ELBLSvzQtmpseD+HOEs9lJG
Jyh01Dxeo9WPcQkAs88rmwmimeH4V9RiFHUicEv88qEiHJcBzuVHguvgN4S2wAaB
gwaoRC9lEye6xFDs3K99qzMaW4TAtm/hXVbxJctGMLKQoGmoC+hdH8QGLS4Bc2QK
yXmTgWldl5hUYXbzYJH9lIjeCucD6Hr/ALynlo6MP6nj4vO2ETli6BLnDF+IH1h4
HX7XvxPV0Z6t8NsyPiQysUjbLX+ZW567mFdKtBh2vvTNKhBQoqkWd9GQJI4yV3n4
xOMHxchrehEkJlrqtCUrIX+Vxh3/sqC1AfX56LibL3ayGsHCecXZnjVaHvinskHF
98Rgb2sbnRWR7PSfMpUdsVV1BGmk7VdiV6xHtlINHGaBsq5aYWUTgUq/U5xg4cGR
Y8jB1DkQjiUpqTAtJqzp5n8n6O3gcKGX0V6I3JZ3aUMVYfuJltKdUOgcEhvwHpwt
bT75dkLhoZpDBbRedbQV/musodFiRaegIufyXizju+/KRnWQRHZyA+ZutTvB8vLv
N8bVtHfNYw9sHyqZ7TP9lBoCpnlrA3JZfO+C8j8Yy5xVGVWkujroN9T87PIUGpmF
b7VjvJW6EpbQgHENpgEZnP6PvQ3y37Q4TzFj/wszkqXKI3uSmW90uYchIFoFXwrs
4HJU6uOjRgl7n+sCB9q42S33xev1KDywyb6FhIDon77V6YroXDjxcEnV1kpO8bE6
I22jrZ9FY2NlmPuzFa0Z0mX1mhMG81s6aN9BKsGfVSqJCmKoKNHt3CFA9ma9TMcV
wZnsHOnEPO3PHEQOHF8MlvV7ZANKEL2Meja79i25jkJ0CvPSw6k8nHg6GZNieQ83
ze3tbUdkxYqr6BR6obZnQAav5myBRIbpQ/+Mt3eL6sHhvbBmOLk8+iQtZY8HWwx4
98g9mDrAVZzmE2C+ks8bgwtl4cCxTitkeH9jwJ7uUBU4LTinp0v3lAjk1LFZUJS/
tNWq41aXExf8cuE089U0m2d6MVvX7PL3XapnJiQ/G9+DGdyYw17Bs32WmS8JuovC
XsuIPH9KmFlwd6bUtu2YZk3l904995N0cC/JP0PmYEoj98667u1kKVF3Ga/nLnzR
8Mwk1NfGqkaEPyjIwWu2pN0VpmCzwlAP/y4RNeHVol3YadBVrjC/J6IhdGpw2cd5
wb+KFuHpb5KBM86Z667r3VLSmP6im9dOeKF0bKOy7exUzoUdl08pGxupy9UzMxVY
3mVmm8fS/GZUq7NBFy2Oy+SdWxzLYc9VvISpAPoxh4hobiArZz4nIfKaHwJCpcs/
Nk1qcfH5dQ2zQHmvsyOD1k3bJMdjfSSAzGn3VHbXjqVS+1rDc904i2sSF75l40JN
Y6XoU/JSZWNNFrS4HJjWIRYdzy/PBCkItykWCovHm19pgqr9HKnEx6hHPrq0VoBI
uqQhZ6GrUL0JbVQ1lvXgMFEEfssr1RTTxUpVlDPPEqT7fC87mOJ+Hbmfu0OliE/a
GTd2bH5xYXMjpVTP73PbwioHz4m+VnnrcnDrugDKIW9aMtb7pg3BfLy+13yY5AGk
pfKA6t+p+Z8T95Kn4wjzhZVezOvzHYS1AZp0ueilHB+G5nn8OBaFiT/yJF6nFpc7
w/3ZaldpHtYMmWx5WL26IdL6nBWBf9dY2NCaMr+RpXq25Xea7HwrLJXSCkkztM2I
s4nfEp5YpHiTAVw0a4RKLRUZfn1A6XglzZlRXxmdrzSRYmS5wKOuNKPwI/N2+OtG
NQHk1Hkt01Vp3zULIqLLOfw0E5Mak9v/HDXWx7ivKafcOB+Edvl2HrVyFPd/Bx2p
AXH6OHujssq4Z6cGdzXVMaqt/IJVlYH8itUNfesCiJdUfK0TSYcbfTXWZwQQUhq8
DKDY6yKpiQgiK53zM+lZ9rUoUJk0btFOAtzBmOEwfnOQTWq+QNIs7hCbXjQOWfpk
jN55Yai0XIf8uFHp2s7Qup3s21P0iRwo9g0wUy2k9+xjU7Hjr2GkY1nCW6UGiY+g
I61aDCLEPbpG5TuTiLOgOvEBgMcU41vl3VgdlpoyQ8JT5EZEJtH1cjw0HZ8tbyTd
egc/sWpNN/hMHZNLPljq6u7IUk5o5S7xE1qEfCS4o++QOpq+R0S+zwn5lKMZbBf5
dEe5zO8P53eENW2bfBDoVqQpN8nUjr0qO5z1kTnKCwLygQ3IFb+zA1bJYPBH4ZMQ
Qx2wqMRj3SgTch8+mWLVoNxvUvDmcQS2LUTi7HVrAfe9ZQyglSW62q2VoD3+PgpA
zvZz1P02T/uM6aoXcRc0bQx4PYOJNfRrglBnUnIexgkROXkzyq2c5e3+ntlSQRXu
OfRkJYYSZzOQOtj4Hun3nxIIXMKg897fWGs2vlVCjNh/iDECv1iJXr+FMctRycMQ
p8yQoK9yvnkJW95INUt9ahU0R1t3SiaOgQxICdQO710Y/fg+UemKVIPt1EPqQNGw
nWiSYNlNM75+Bd5T01kmL9VxjH77U51lZWG3jbZCrb2FQuRsSLPro+BGkuvNbb7d
0DAKzv/w5S8zfZU6WrfX/tFTZ+1sVWuK/P/fJU+rf/gSIimpAPcnI6LuUEpJM6x5
IQPjz89gpR+kjDW1m9KolbeSxEij49jAza3TawShUYjAYq9w5SQwuBQQH9kXbA2v
T6DCp53C7o5B7/CwBrbZcKBfPQxbPeN5uFMijIe9bXFGLOS0Z+AMIWFMoib4kpP2
BqcTtrbz8Gy6URX1fEEvCdhoYLyAXGCWtEzX7FRgkCYx0pcrG2G1Xt1K5vLnQMiM
bOw+rbClLF4p5f/In7N60ovnC2F1yvPLEWCX5YZ6V3stz27Fxzr97pmd7bcK/tTJ
mnX1r5vQW0zXmrfCBE7CiA12ocVRwdr0pnCIkgub476bQCi/LQ18w+IjkptIbcYQ
SDxdhwG4/aB/DTQwoGLS3PHc4ilbVZXVz+Oh2CGJp4MaLukiKsUuGiDGdLcT05P7
VJzEeQERQn4UhcKWWzT6ec+Ifo0vOoTUGiOfjl7qbtNnJASEo216aciMcedSVTwM
nF5LVLdCFXXeql79dKD41EWcdETj2J3X4okqXSdXSUxOvQM59KEIkech6nkVhrPk
ahCq5FE8L4WbzaPP+MWWc9sZpn0iKl67ZtPw17u8ije/QsxQaqvxJ+1VvdOY6sIo
u7p2MDxdtO6ylU6V80gjnaKAzRm0eXCjH5NORlNJqUXv7djXTU3gj7GLsCq7pYen
AoLVT2LIrvxS4Rzay/FRXd4YBdufZni0V/dyM0hVkJZsIpg9uanIN0M/tvDXKKyZ
8VHV54u/f12t1f5jDoAVA3oR1XCW47FxqT/67VyEEc5R7x8AQQW3/cMLQMBkev6T
Ey2PRgCEIizEkDhKkbEmO32T6Evhjt2aewhfhxIc3JkOK+pYD8x5AutevVFZMeMe
4UvFCbXWVcMLuh/fkh92e7P/Y7V9xs8Zbu2s1NEXH7th7n69XSXMHqwLbHKHKQA9
nVrruOKXbooK+7LQhM5OUhcqHli4QChiH5lUve223ZJcdk0EazQhFv6V24zhGuqX
F+eBwvx7oJ7uc8kmwTfPmBFAHbrXQGCN7bIfvN5lh4hzGVAWLl4xxwUEuASv9E4p
L9BE6Tyh7z9j38SwfntESiI4x2g0uE6+cuFtlnFVcl5bty1rA/YnaS4k6ml80jy4
wLkF3xNCkw1bfjfbnXG1Hp8DuFCirz5Rc0ubTox4NjcUmjVeaU1XZo+300gckaB0
3UPfpS+8gmFudvs7HNjVknwdOPm7p0Q/Q3J768Hs010v6VyhvXLnefWGyBo05rsx
lH8+WzSY01lWDHiElxB+ktIgK/8M1Da2DJCAp0ZhIsYO8txAiUxXXkcAdJzClIA4
ZwLyZc2BS/D9/q+h7Vdb1zrsx9H+DdOae9ZJczZVcBO2RmYxUKXP17gHCkJPphwR
v/D34klazxX4BrvxMEIDdVYJ4Z6d+//tul38TA4DMuZ/V57CbmxMW5XKNN4umrel
bIhz9xQtO2i+JxgwHIw+T3o5nMIKfiaF1HF3CwKHy0Z92H8UO9ggaMcRuv81TcmS
rPEhKYKuPmXYmKciQrr18YUp0dAUY6mF1JV7770AD2gtWNJ54o7fxYfh7qj3NM+l
kTwdUMlJqAgGu9l6SU0QytbjN2Zzd6AKid0U+NBGOD7YfQkBR+DbxGIiB5cTLvxW
WAqOA1yiCmaRswfFeR5zuCwcxLi+Pz/HonrFo6tH6c0qjzYsVl9O1Lrk02U9zgUG
vm3SphWpy10WquEF+xRnoGrw7ucPaJN2cBWNQ/8ADaeXurYBF3LAFyKsH6kYQv1a
8ow4+d/ghJeD9rHernBnCeRr1TzjmrnV2IigDyRDsO384ic/W0Cz+lHU2XF+13/I
v98p1e+vvZu464w2KtPgV/BD/yuED7rBFs7oi8s86YQzu6uLWiiMAUtdXHL+oY00
CUEVlJSFCX4Cq4Gf2sbCBb8pck9PSuc0cAXnI5S4XzKygnFOc8WMIDWL8YIrA2Rf
URHRCN5DeQsEi/HV4hk/gEKS3KWigbtTLl99dF9OqyqizPfCvrfj+AQ4nC/DZGAM
xZtL2PpGNLVxn2vZ/KH+IYxTk4UQHI+7ZWwNtV/JMjbNGl2iY7ZoSwwxx3Jg8s8X
DYe+Nhfk2u1D9/XIxgSWhQSvI92pcX7EDrrKhor9U3Sn/VrLm1NasnH/oe7/q174
DPZvWcaCCDlhKrDEu9VYLr/LK9QkmzMCrUx3DzqEO8zJ7i/YHYwT4VMROTvvmxXG
ZA3csEkx1tMPpOBAE21g3Gr4bG/rHPtYdDF6SngSlRRTcd8el3D5HlBpHGpG8tM/
cOJLv/Ud83ocM33QG+Cso4vzgnhWGC6U5p+5kUI3Zbq46a1pdVFZr9RVBZ1cCM8Y
qiz1n+86H0TkZcEzby1kKUo/8aTd4i++Rb0gVbyjMUfjnDNMLn6TbpXQV5SQgjTX
H3upTrK9aQPZWBXRc2YE7Xh2CBY10rc+CFGC8NPBj+6vEkCu1aiq41SpIKsphHGA
eHE31WBqTCytleBjV6FbhP4L77Bn+8I3eRGTm20M4uPtQ60gCueVm6lttWSqvXwO
8sHLrYkE0A1jQZr6yplo5vAlALtqMy37orH/LuKq9IyQiG2pTnQy6Gk3hoZM7unM
pn4d9fm7knv4b53E0vLLo1TAJ5/u1Xu40vyiPOScIwCLQkABKJN93xTVy9gdZoog
XGYx+HfbEdHK/geNMUZxgc5JbGpZkXbjWKIqkfp6HnrIGR1cUFMhhHsYqOL0qv+B
F842dVmJ+QNPF0z0jvAFiKgN8kuDwX16R80OWulHiDZ6Qzk+VU1fplG2Ec1CZdKP
+3+ncvwISsUmZnZ1pqXfL2PWMVYYj4eER3tWfWa3rS1md+kCvs6JyjyQkBQ6wtsj
+EY/mtkFdllIQBTTfegE3IZXo8dGPGuzJfOG/Y/9B+vmt3HPtD1SrraHOHT8RMyN
kVMmX9fwgu6BKLCBOVDiHF1KwMWhM5pXyCE04mYxzcnFESYxSLRoQTNqwKUaB/sY
jwAw0FVEbKigeuFvW8AlWlX5gQ+yrIwpYc098bjJ+EJzf7kjxQxKGzVCl+x4BFQt
h+EyYI2jBA0Hvwz2Nd3KiffOO9JG5tmTcmqc/FJNBkW7ZBAhPnNMqUE8OwFuNgNq
3be1B8AUzYA+ChbCJUI3K72GomJ2sXum9wnNd/OcJwBPXZJoX2yn3N4ygcWTUH90
duvuNZin1ppaUm9LSr9LSIzmjwa7blC8xgxdHAcI+0uZy2B8AbdKOsllT66Vk4hJ
PMSffjX5amWJm57TSVvjzhW2lOFeYpHe3gnBxEkVx97MhafNaCWAYQoByUCKWwwq
5Q8YNcDbbMDTDFdS/cGyDFOCiG4r3EuGL5kCx9Wc0KRAppaurnrp5ujxGZsW3y6X
/3giPF8PUM8E0mlpkUQYZGm9CnFEunI0gB2B9KAxfFdIIbXxDlKdBmtapxbUvx7h
dhgY1LeDYHl/KCk1qrqzjEcibaaYI46BP0BCrhBWxOP1t3NjgrqMtrpDrCeSBb+U
FVwV5Yw1r9T0BBoULco7bR9lM4Yx91BBNGDNxxJ/QBJ19Ik5sGND0scCh7VFZIjZ
0EsxnQAn82QXdz3IqSuVH9ZhHxiJ/ApRjs4utKKpOZoZnxlfJhWF+sd0Q2xx48KM
xGt+ACuWtRwtwA/ABrkMlFZAlXwQhfQDnEaS52yW7oF+QfnB7rKr1Y3MvZbjsvWv
ONRLdE10hYiGnVvLWToLYs1G8FmDRKJjCe+pR897Jdq7O76n1P6ub2hjaDOjY5wk
K/BMjaPx6V+KYfynTUP8AFU9Cc3AZ8b9HAwuc3OzQmLTz4BlCwaQIIuj2LG5yokg
/ORUO9uJfvZBn/S9B140xzz12+GQTiHRogRtEVixJ384kIrU7wQOj4PIlRlBDDTy
DQDfmvKOSGwLeNvWHJwg7KEUb8m6hGS/z9wUGZysUU3453X8ugM4BMU1ZCCShwnj
vL2zo+fm76EtO2HxS73kHgnrZ23cOWaw9lxgsuZPylY4yk8wsGqgGLakLNCxJ9Xg
Ul+u6NAP8PmjoW0OMlYcV3vjQ0DF+g8xfMdOotOP9zV9ENfqZAwBgPo5yVf+QZk/
8DBV3U/RfbWjkDi50GC5542ZCrA0JapU2lU/njdEwjjxFnC1RKH7UKE43vEHqPWY
mUTUDe/KMsak+1n/g3d6TUE7X168+gjn4Sb6UsFaCy9O/m2KGgvT0HyL1x7mDQyl
jLCMFCml3e5uCBbza/x4ZRHIeQcChkQp5QfKwrF1X5CW04kY1iZ5p4FojM2Ufb5r
7VzYN4KpTaWADSsRWvdODKYvs5qIJgWJ1FkM0ZIyYuoswIZpwUGiuGVNw5d4Ii3Q
tK0IUTRQgrqX8SZWJrOecEeAyPav2mjbqh0Qv6/mQBcwV56cv/jzUU4aOg0k2qMn
4wGJGA5zdR+UhHsssxOEqWXAiGlauY//ACfYytIwfpwj+TNfJnaxbkCpW1fMi8FX
v+4p9ar7H47mro6Q7+ZyLLTUViWybBUNXXRUIO1uo9IfwPecCn/rKSO8dQKXzjzl
Pl8rJv1gMlAog7Y/LD5L9W75m1IJ+xMMLX5vWjvQqyLJr6ggc1tZCV5GpBe0+YAo
Lj37FvyG24wLmBiBIVHIIUbJMe2tRblHx4TmAwIewhPLE79zT6KqWGer7APGJsID
vTMUa+ZXH0ApZxlwvLcFyDKHI1CQUllPf7NUWsKNmWdNZ0G6wytfs/ybWlHXk3eF
e8SVc15Ug5mqngD1/20dq44K4tx1dSk+8r5zhWaLPwhS1F6YL7smKqEgU6jiy+Ol
cd9jJRls64UuZqvWu5NR/YDWsB32UTCg5xysuuwdG+Ck5XmzYJVWgjITw3lP8JvQ
JnKygtMFJJEccd/rB+W1kH1Oia8LKBcZbn7gYab84sPv+FqNkB1/deYm+uDfVi5v
6U2Z76rRjC7Hwm6ZS4U51sB4MXy0UwU/YxjGAN81ATjz/2EBhMVPcpr6iecG5n3p
jtrqjOplY37lfKtyL4eSA4Q7lYyR7R7br9rvxJsdyZt8xtRBg+NYAiOPQxkDg+LA
djQpxklHw25RScqYYx5eZoWGnBSZP3mHbxM1eko5nsFc8c4Q3mZBQ8QgYKNAYUpt
xCBcBpiVTOztgwxADT8ONsJswFFjk9RvdPa/GmKE1k8HuG3NZWHV4E8faPG6C2bD
K1N1sXT0MvPDcBH9xGcZ3tF4qIntXfd52n8TVc/3JsVBZozRsoAp2tG6IzVWqz9G
RwcJjBlR2Dju7uXIhEP23mMMMDpeDf63Ne62weXXerbcpx1o34M7R4CSg6nxiSIi
5IdvVvGuIH9VvNgDRR8NS1BA4kriYjhOulmj5kEdxm0xilFAYT/ckddACvevxO6O
KqSb+ukhQyofmuIFx0ZYOr9Apxpavi5s3xzUbzNTrFTC+wACoJ+Aqdwp3OrPEuQO
4hjDXVAr254YrpWh5U71ybfa1ffjbgBFcNIkPpfYAH0e4fDNmOiyznr0cvFN27YC
tKtcFp54+G0+/5pMf0a4MJmw+QHFWKzvO74e7bY4mErhSL0CN3B9R3obraesj+dX
5rgKpxHvt+9M4DOgOKpQAmCxoGAN+3aD7Pb+rdIhUk04nmB+O1Tuba0PHmhdRY0c
oozExShxY/zGFP/qgUoDPm9gSJuwMQS3c6nWPPWpRGWnuryboHT0yiQSajcchNaS
kgxhsZ9Cb2/tkS2Aq2Msr5rqsBvL0f11ut9erVySfmJOJQ8psXVjnfn3yK1+Qiw0
k9lbByWphdmXj9+RlMqM+6yWVNuI3ikKrPgzmH3u2eoIr9Ujt7IDxg9Xh/mwJaNF
Gn/NBpL7jbabOMoP64ZojYUCy/kguOmsxt+a/v7jQeicv0t1K784KW7+HCAigcop
gJZw+zdJc7RymGuMk5N9PYRq3kTN9KVrWTYNjPKg02m56muDVrGp4meuy7eVqo8u
fowuGD6MAt3v7W/uKYTV2ut07C7D7dKI5vk4OTr0fxh/p4oZhi83H1pJrAV1F9Ec
Pyp/4TvHrboVI8auE3pm2AX6EJF5NL2blapR3yKp8+zgGqxpCyJ5pPohEeWKkXUO
hDF4Twxtd3ZpVJf9wTTIFJxN4Oddpw2SRjeVBQWSExcERSnmYKx6ZlG2kUc1ZLg3
VkiTIHvr2OqGT3kexJATihFbrOWewJOA2cQYRPCpgPXTAPL0hfoiHGXDZ8QaPyb5
hJmNr7XrufSnIyjtJrIYNH8FNPZ15/oE7ahNe3Y0W+ttLm7GyHI7eXZS0AUgV3hp
Jng9Wq8wM4Di++kL22gXdl/ht49hGpDtgRasP5YhKmoaA3sKVj8N1Uvag7bj0+xq
0Z8+aCK+bYQ349zAK69qpKzCl4fEC/NshVC6CIFmHx7Wt1fHj8oN78dero1bB31k
N7BBq+tx2rQWpyDKg6PV+hM3Hj53znQz+C3JRNSqsc1PqBzMOzFsTgpP25ZJNSmv
7PBqpkdtP7c13wK9i2inDIn/+9lAOMXYW7UOhBzwy8FPRgrhi4KucxP8iLGtf00s
c1enO9wgreaQVwLOaLrnAUpqH/X2H1wnsurdy/b3JtewXb0qhopjjVqQe61X/AJn
3FG4Xa49EJkD3czCyLjQC5uIIUfzlImWKI+KzHXJppq6CcG07xnnb5sSZ0kaSdi6
aW5/ZjNT4NR6xFhZtNP7CSUGDV7Ff5QJIcAEOcxWExg8YZyjZRj/iB7f20oW9qqD
dcKJKRlZ0tvt8xKeoor/P+XVIZTgojkezeI9K6Ejzv9KLvjFgcf17WyDDYdRQUDK
zuMtVlkVdGpjJRrDK4yq/6x110YQoiEI79Ys5HKsui2xDNYoccqWoqYRzR8TNJ8F
xCY5sdrqFZBxFQl5DFkghxX37tkv2ADyPfm2ilLtLcoeRBxrXNP96H6GbH3RKBsT
rBuJ1QTOEvl20XxxURdE8Aqtq208yDPce8LUd6OCw0cAE3RoTi+52B4lI4vdlTJL
kx5EH1JVczNjwKedU+7fMaJMhcPChllYwOx2CDWE1gMa7DsZichr3NbJlsQwYLHI
r1XhiqcOaGozD+cBmQODR/5bp3tfho3GX7xF2Vw5Hf0AA+sditAb19TjuFPWNF54
dEPo8JcaHIE/XU3CWMyiG0dyPzH0Hz6XyJI4kRfgLiVi8IllztUn2/IszCc6JyQa
LeUp4YyJpoGDuXgWdkcybcv5y95FylecIlX5XasI3ZhZb+0hXvzFxyuJejQtorgR
cyf8o7zZDHZFZamhhsT5Ku21m7ZXRNogdMeFtxu5mk4unWAzKE+rWIUQCN//MPC9
pkQ/ugQ5XPQR0HGUPa9YsqnwGR3m2aSXuFAiU/c//+A/piWdJg217wnu3PHJwY6R
bFwq4kRdDyS8QMY9FvLrewFez376M436tgkqPcIrc87z/EISjmMlbVtoDnvrBxuZ
teJFFroz0ZnX2iXmEcIzzcOGDa6RwOpAf+r3LeqmaLs1chzPKKXRGyf1tf/6jiJ+
FBJDrmbHoaNRWrudk2Bp1ZE4HfILByOVrQ72fB6WAJi8TCwA8muxh2yPhfyYOIxf
cUivcFriMPtNS4PUCXKepVLGusq8u2kMqBWLfjIAWqHAK1rZm1mcSxMwPNXHQwDA
qfK8kvSrqK4rxx/mBIwG7kNE5v1zYL+J7+mcU4r/PuidHOyWsOkBYOX1bypjhvsh
LX4tfstyWTYOgi6w4FobWzD2R2NF6g9CDMmcghNagpxDwJ+gG3z30vZxLPYp4OMe
lTA+WHBlMYm+wPVMQc3JKPj0PewZfjC7jxL2n7cL1xU8jTO1SMy/mm8rDO+RuJ89
JO/zAOMUNOyQkFyOO2Stz0etSWWu4uMayZGteVl/7jT1VY9z9SLldjoHHUmehBX0
qdYh6yni8xlhs/DqeiBLOHnA4KQgup/KKj7h7wJYQo95VwgwsSj9ig/bgwcYsSff
5CLQvlbzKSglWghorQENpioqE8aHsXrZraaS8mlZCYFdwyVT5aj+CpCsYiOFJ+Yl
p/IQk53YcXfwSm63xvL91lxzRY/zElYkscff2KByL7e+njnlsBfOQSBrVYA8hHYq
0LyRC3MeBgshjWOVBvbOW+yL+BfXr5G9GKakqwv5kTPZplD3fRXbeLR1ICfes5gf
V9W9fyRBBt4JsB21Aui1Q2sUC2ykKfOR8TMUUGynJRuev+QYM1VjEK0lnK8uFqGf
mXy266G3XjGGyvXsSBYdiH1dG8k9cb17WeiBke97ekoSvauQoOKwMiEnFW0t/aIZ
MGr7eowl+kJJKpMRnWL9Ljr3dGUQOWCUme/3sw//2O5q11pOdGjXthzrSgH81CYG
QUTGo0NdX/+tbvkAygbXRZB3OF00lM2MCMoU6Xrlpf5xAm/YcplTuF+Bt2HFxkl/
P8Wvyqtt1n+nkb/Mj77bclrYuz7Le41wlX+6zGl6joYcU/wU+26GVF9FqeEgbneh
exw4pzoxXxgGZeeUsn4awUldZ9CS/6WqcIBjPLdww5VWTF1Vlm47gLF3G+gDZarr
r36mEezNbN5VkuZProuC7un0/+D+1Xy18TYQDUy9fm3JNa6tgZWgqdy6QWQ1W3iE
evzhv46ALxtjQ4rG+rPXvyY/0ZkbZOy4aDa9RTJYMr7FzhPaA/AOart0TMXrvh6a
O2trkgdsxL2hWBMKh64y2w7N8AJY0K6r9qALu9TWbuXkPe1DICnBFUve4yDwSdig
QuXw+6h9u7EpPrSVUodyAAcV7aygShp2FaTYmQcR9M7wt0O1qRHfC3DWEIMvQsql
+IZSZz/4JHPilgWqoTEcz2otFQ2w5H8VLUdgT4yybQaZ+BEoUFrK+0ERE03SYXP+
Vye4SIzAf3cL7LssMqUsCqHga97TVTMnB3ZBAqtJLl+kHFkyv2VHYpWZYm0iIacl
iCxTnxuD/GbTkakeqpfWtLyZIqpmlNBsQ8Zn68vOA7Or1JCKneFSMBbLKSX70h5H
amLVWgV53qn74j9OVmjrGnVkZLkMTKqqILCXNVcdgQMRbgJcY/KSaKnhQY66jy4c
lO5yEsXaSViNt6nubLwCBDFz0h62op/ipmAtT4YO1yT5bwG05/k1NVqsBaeWJ1VJ
kcz8MQxf9tufyp0bB1pPjA+o6o1KjxZkgvgSb4gMGN39Cn+4NB7vD2OSIxLioPrd
npmhYg1BWW8q61P1gWF4GWz0A5Mt04Nal1hpiMmoc2UrOT8g/oJ8h0TuRYTizzBy
3tclH57o5olW+qpVdnZLCjzx2A8uUonyGMdzlMTtuWEImHHMiT4z8kArL2oyIJMq
9/fsymS1CPaWOOSEAJAuUGz2Z7Li6CF+biSAQHNJJ3ODOkMFQUB1kbbKtztnTB+/
zbwmjONb0ENhP97m8tWsJBilPv1t/zVFs02AGuwnoFhUixspkPK1HScgLQ7uQBNd
ju3cf7SRkwjKlIWZ9h2uQ+kFpTIZmCTXfy677E/z5qmdsrwAIpB8spqBU1GGr5NO
Tlsv33RD9X2abv9alggTcCjcFg5kqWEci50Qt25+py0QWiVTbw52h6H87E4fXN0Q
bgnQ47m//QpmLmlEFF+ana+z6DjHoiXxplz8fQ5zpMTKxLPCndySY3UXLrRxLviz
uuEYQ32ROrCGZTBHjanoUlsdPmQEhz3C0G0mo/YE/TtBJgHRJt+ZI6bBgKXUSa9/
9/X+ofXz0sdrqQU6b534b6nPFiRF8Srj24EP3Bl3PnJDQ2U01rLt93mLqSD4QD4Z
v1/lZaDi3Tz0sBptruRamkLBPfv1Jin/rEijGFO20qSa4ntemGx3QiEhrVrs9TCA
8r20S/yKEz9pBOkIIfd26NnSjOudP7pDj/MxbMNUhKA0aYL6wdHCaX9Zjg/0EkSw
P37Vzz6OiIjvqqyWqTPeySKEQKW8lIPwKTXkGGXofppWcS/n5XKlf/HE7OVOnYYR
0PlCsgXNDSJTD0w7KhSolrMEZeb3DrMELJ98vtfAhviUjlbGj6ykHwACfGhMqU73
09Ff8O0uRBzBQ8uRKBoQJutLmOOMgFxM4iKvxwY6NsqlUnECn9MocXMZpbnX5pK/
70u/t8AyIVpkMOgTxWdGK5txrPcXhaipor2aolxLzpNZ4Y2Yr5yAoh2nR7JuJ/Jv
gPAg7pGIj7dudapkDw39nxrFLp3Mb+eZCl23XoanXznoZiNLxY/w/VEWn9iiAPKI
VKmlpc59JVgd1iUSaYhwHFtICmFF27VL/DCNO+h67yr/LQ8no9m9SGBr4b3nplYY
HfovqTd7bPaQKvE3wZAwyskD9JRcLBLcnJOHhh1Vpev1xEmZenNyao94t9qPEkNs
wVUQN4jPSAxUNyjor4+khERRxh6D29DeBUTwQSR4uzOuUNg7IVf7IYhIAE8uZpP6
ra3UVz/5M+C5ClEMT37qJek1uRIzXy1Q0EVvveFAnAvH/qEm0ytFw7kuZfowJ3tn
Z0jOWGvEyyhNAYMstnsfNgPITNPwX4G6iB81KdNOTdvMatSgMnECtUhdPnwgUa+8
fSfpPD1wUMff1oot/ndBJd77pGKVS+FQf1HXOXPCTtlfG6dQo0FdyCBRKrgNQiOd
y5c/wjQRHRS0Pjx9di5k9/kIkO2suIGozTpqukwx6bNN4yttG8ej9YpeHDWT+uHn
ZSDhFWt8gNQwgTokPne7wjj1UlqQXrZ1vSxX5gBkpxoONoiwcUYxThHxoxYoHKjE
BCDkp15K4wxZQXf0FwRxO8Ie1GK9Pzv7UZT4AfoI1vvks3b+Q/v+mUBwzNiXegsJ
1VMUzU96xVLuMaLiyTHW0fyJZAd+Q3c5G0deIBCo76JraxdXDHyt3ttVs0wjihKd
vulJM/W4iSnWYjt4uDRc2o7f9kXIsC+d2DPiVKnxlvbIOatVTEIqwY0RUUxFNpz4
n55G8XKgvt/rfMZsXYBk8uj+6gP340XC7ytwx0oQANMS2oE6UH4IEkc8pAhUmKEC
SOwf9VrvzC725nEDVOhl4yni8xjUbU82CxtNzc146ASqVeeUHSU42B/ChyX6RjcV
J+SgFlwp/rKiPKRZALCaUTe+Q+IK9OVMEd5oVgbx8YHRVa2TdLunR28ZsR3CDLLw
ahxKcvlQFHMSDsKZVFm21TFFR+B9dvGipCnghJE6P2HjYwAt2VXmQtVooTC3iQkz
WUyh+qfrzJ4uVsACyxjymn7Nw1qmlAGFMaAT9D2LN6auy/8wl9UN4PVavfTDxBHV
Ds/1GAfhu9Id06TYUbq0FjFJ1nBRXwOqCDk67cT9QGphdMuzYemgwmE7lLmDbisW
lij2x/KYH8I9hNDxV+B052thJB+QaToZDtzF7wZkp/HHLOVRGU3xLXxQ+JVApMcX
/sQD3wELF6gJcDxxmpA7HcZviQK7ufVteDtzKct8JwaTkBcw3sKRkeq+avSN5ux3
CQ0KX0LDkKYEMpr87Ottc1KbQ1hD2Hm3oe5owjWIcFPGwAO8LgJGjEdsEf1ZahkM
ywOPpl1/9M8GXkuFgI7emABAeHsVBY9DNah3jnKGscrvLVnhTpFfI4fdIdjhb9IH
gtUyLIfn+M9/StYFx/iafk7vh/Mi67pWKHJAChfDgl4fNex6JzdG3dklxREyGqMu
OzDU8CVSqYcesbhNcf3C00Ax5MQRQ2EWhmnz7vIAuW+IVoj8jnOGh6FfgUq7zulu
gTizXup/pALtCLYOBEkIcVGgoil4cwXJFqAInaLrVubqzHWhSw3yGqkqRvnTkuxQ
Vr+Kd6MmSPfKwqVGgfAoWL2OCm5rPn5hr3KWeiv/0yjYYF4dG6uwjLZZzf8tjGCT
vzKL/0eXqM+ZxfDwLHTwq5m3qPD6YnJAYQKbCwau2rH7O8stGPyUv4ux+O9dbLO0
kYG5lUru+rX250R+ABKDE2I6MKdMVKENMWCVDJ0jyQIrXpZz+5AW4Z1OGDcplWW/
IK1xa1pBEb7OipJ5U24NeJp3me2pzF00fXwydcqx5gU/KIp4Pra03v/3naeK0FMB
sTn40MEmKIkWOS1ABOrvF+eimQkjRYNLsMYzXFH6Kc2FyDih1QBFkXwS3tSj5bMy
xIXgYcAgqwTPZam/rGkJW/w2yvK9Y4CszQu7qcg/e1WaLKJv/B6bMwniIhCuLOUH
cnevNXoBbuvBGzvJnrD6rMTxqxlHSlLBkAG7GpPuVB3aI2m4t0hKzpja/wQc/cPh
WCS8RWTiT9W3TKn6zIrmKaKPbvkWK2kQHuHtdaF2/Elt/3/tjOfLT7DanH2bvFMX
BuQpHz7YTxfI2zI3m3LOUL7DJFAbTOPI5OnQdMMpa3akDVSDOYc9TlQuWj/8MC0t
J2mlXDgXOOtevpWq741Odp1EdWaYNATZhKw3eVTkpQuCG+SFKNt/OWaHnlzvf/YV
kgKbzgafHjkZFdL+5hgAjl2RaGUi37t4d5xrq0ttJ/0+cl9XrI1vXPxOn5ksdOFb
uvtbC/H2rdrSvmzjDGEPL2OpLTDkV5Fcti4D93xm1fv04oEDg1IAuUVTYVufKy+2
Iswiu8Ri6dxYMnVS5SXFnVcM/QnpimNdNn8ClaIj3x3yxABk+UoQNS99o94OonjA
6K2ajL7wOanMRR1R0TcvTZSaLHvOQVBBrd14//B2J1bPft9eAQYnuE1h6MGpgpCY
pRk7ICczSwl7DSThxVlMiJyQ7inxKL1AfhDydfKCkJyVZgvJgOHB8fCJYMA8nctP
vdc4zwTs5RWJDcCGMJB8u0UA9mkceT8xRy4H+0NlQF8PRIiJK4mFLo2FyFvxPVQP
Uvxwd/svapZ9wplGO/S4efaek4wTb/1r3ONvgvJjta79uKeN8K9IVCaFTEbv0wK1
nOIS5+QvgX4h4SlGotVxuHS5liUjWOrtJ2WBFv9m8i8YWChye0VLqDQzlDgVaJ9o
6Nb5S/c8OgOpafuMQCotS3m/sH7gPmOWMuV11LdYyMt8ap3UQRhE1gW7mkUSdEK9
f0HiYb9+vTl6Q2vS9y3S9UhaLnm4AxJVgVn9Rm8w+HyYN65MVhk/QJOoyzrec06u
gPbP0LQz8Jw2AZ20YKUIPIJ5ZLw9nJvBlCMC5Jcw7fiHyGBnDz04UanuBsWXNnck
dKhs5Q4ne9eboWuJMs8F1iSCV/9k59TWDsH29Oe/TdUHDpYCqR3KuKBPpfEzpF3N
KoltTOibShJe4f9EA/Pud5efQhSbXLIjilB5X6FX+ez/uUEyH2hMdIMh1IT+YAnM
isKB8cvsnGFV47POilOluRGvHTvU9tO8okaHfkyxTF5eW7RxT8D+Scb4DWG7ffaj
r/TTkV9yNCwvcmfU03zNOAYdLOOL8oqYSSYnTlQCmmYpS/m6hR5SCzuHueQZNvDP
7KGqxgFzlnlaDoah5ST12Dso4/feFX1fVAycNcaBF2WA149RiAAmQnNyK4RmzLUo
QRZTGNTblYFnaM7Gw3Ikt39glw2iClMaykG4VULWaXVD42b4393aQurBCC5urPyz
sYizGzYllCjZBvHDzUICzfZGmzMYXU+9261829OG67TBmYYHEqApd+J4lYJbo/GU
0a+ZhkDnts4CSN9Uh3OOTENxsZKSKIHZU7xkauBD8+OqNRhA/M6HHKWw9qbZLtAC
2lOMtOWAwOkxPnYH8VqSXn1GLXo0tgSGrfWaZ7n8JGco2gaq9AEJVp2iTghqAAK7
tsA06pJ/i3pagGmjeygkq1+PnBOk23z+Ymo/JrX/ynZ1D+0nznooqJqFOHqFUHwd
B3T0rZ4Y32dvDLYFgAaAtGHAmN8UDG1/CGGM9SS30vfaA/ygHykSqgXQrWN5tj4d
cjm3psqsZ0XeHUwiINkHB9MeOwYnujL15oAI9xdKAvIW09cDsNAxXYkLgTptqxtz
p35ktz2pKtY4y190qDJGU6/EpeE4m//YUwOkUUbjfJSZ5CX1i0KX4tLt489YyQkI
dCIqVGUDZof6THx3FL8OfZnsp7Qaw9wsy52SGGPcvY3Qf0UpH8xFOoHOXCV8NIGu
LAq6xUk/34yxAFthSpOtJR08O0FxrjCLSvIQhVuHJkmGT6Oarg0wEy1eERXm01cN
yiTn5cliEsNEZI+vBXeDY0ZRSEgX3ip9lSPhT6E8VZNCnaqSYuwRx+ZTNt6CX9hf
SXtUjqLbcs5pUGw2RudlCFtXk7qTX3Al0sch6ZNq2WApQv8y/H5wL4KSdJlNbo+q
1y2tUGoNLuPgUzkRBxWCD2Ts4TIqCrUq6fynwGY1P7ZKbOKzmIE4jUuMmZBqHyec
J6PxmJHUKxh6TEYEMSWSQk0818dryRqk4U/+kuWkvO4h3iWwonxitXmn92GA1Trm
96SQI2toFNBoNilIZIE64fzfxm1VbpR+rz6WxcAvjvkv6WKaEvUlN2eAsR0Znmpi
ALlUR6iGCePDcrr7BxGWceY+NtK/ViqG0hLhTBTM/JAlEhg93cfK7KhZPx9F0AES
vfMDN3jSNAaO3frP+y1wz+b/eCeV+bsTQa9uuZVkQk7SKnCSRy/oJDE4fHfFwxhZ
8a+DbIrzkWynGW2OLQDGQ+qvQ+CtwiXgxlZjNmiMLXbsCwa88LYy4MidxtrKFUai
XEvU7lO2CWSLGTXR3yjEG8MDMTnIHRZJsyPL6EDrHqCKh6nca+YO7WjjAdwOxLhI
T5r9b1FK19ijX9e93H0eNsT6c0JmDrs4sd3mU7230lUFycOi5WW7mJFHu3hgggXe
CXjwPsv9uJJClPjjmeVRYLA5qJRUrHkNQLMUlpPEgW/1sNR5Gw/fVPhbvBnHGB/J
`pragma protect end_protected
