// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:11 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LatHWCUQX/u/PYoY3y2kee93kiS7AHr3mudpXy/D/QdDfhtGO8oeqezxB0kBsKF5
5RQ/xChA/NbpbiXfqXVmI0XrVFysvD3RihD2MDxxlAIq8h7MTAik6cnW3znguE6p
4Xv7/XQqmxdofZvQ09I1IVTkVyuL9fCkTRx1OnFs+b8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 135008)
Buz2PVrbqr+QQy1QL1SLtLObTXsF0zGTVeilLBkInT6Cne7IxjqphPrKeoTHFm2n
d55SoCSwAxiSKythyDd5TQSXutIScbMpCYha1QFitIePswCGo/O24IsmMMPlhMEo
FF8bngNN8OszXX8eP54nxs7mrkAY4WxYUmmOlkiZygUdiyJDA3xTXbN5RcLqCzXJ
UVbN+HUgxu/qD1bv+x4dokxyuJEXs7fIphwvrEoZdctwNqU4BIe+4pLZFbYvkS/s
v9xHU/Rqwowq7Ljg/uE1MfBly+7GuEV5Jx8pvXlT5g5yTo1nFrAuJW6Ayv1b/KKd
q2WK+9qKeSxt1zS2cS0gTnElw8MhnV2zFnxO63LRs14L7buTzEM4xm4OHByrmijc
JRamZ5GKYrkdjFCAyHPj4mAwu1tQS3NuVkKdXrlq70lXANOmNn4bWr94JPf4te8C
U/ycM8+CX+1ySX6i9CEdvj/kbBcbB3R256+cjY8mMhTbPp025AlIY4LcN7y3z1D+
5KCSiRzEZxY8RvE1xC6UEOQUZ10o1+eQ0d/Gb5ZmD9mlZbVtn0Ugu+lOiuLun/78
SbHPOjTwjxMhB4+9dIOHKJfEBSbPKA3bxBWtZu8Ysq95DZpX6D6JrD0BxM2k+n6r
xZtFPNfiKsnuWKYYozt7zinrD040IEU7c+pm/IL/hEdK/N1IO22hMOiDguOS1VnR
XU/55Lbcfjb3jkGa9/Kpqq8gzrRgGW6E78UJNO+xu0lpU1JRi+ueh06wwJiZfOB2
w8LLGz6j2NASX5Y0HxfFoJQMum0oC2UnV7TAvjeoqu1F/8l4omnAeGCIq2im0Kja
qH9cTXYKNUucy6+YYKKQoOfr7xL21ERQaV6yOiCkq3a6VbbKehSsIYF9T6D9MFnw
2k846LZShm/5Fb/sOF1VSoJP+/xCTXuzMO4Dg/lU/9pJIg9MfzjeqDDAr4Xbk92J
Y7/wdsgtvPPnnEHAx32Ortd3kz5iPufysQ/mHoxJVpWbzzZhTm+fTWk3gqeFQQzu
WZ2yBgsaGAxaAnzLFbpaA31Zh8xHVsGp4NAwiWynjUFZPNvTM3S4deEnagy9UkTS
Fyio0WRUxiXLJgnnIWb0zXijpXqa2XHXcgipNceo+VKNwAg5ToxiZcttK+XQhGkE
PJLUOCd+f73/30TnWML3ZIQcG2eO3kyBDxS6cvAycFeM+LfqLw/5qZhWzLeqVD4N
9067snvodqyx9PHFUd9+/Xdv1xcM0JDKzE6ZEPfRZmCQogmWEx8FWJH+qkgm/sva
QW1kOU6TttlaMe8dop5K8TPqGpE820IItB5VwHNHuhDKZKk/FzBucpHrL/0mWlGF
z8x6eb6/cjh38s3G3rhho6zswYyvpxu0W8kuavvBLjPdKxgXrstMtwy25MJVakh8
uRRjfcDdnPbA/rpnuAtptf8x6SwauyUGlP2cfvPmBYyAzqCeulRq6NxLhkRg6+ks
IWa24WujwExwHJ0djV1oMUQfTceMmjNbn4NQKFrsQvYTGqegoDTpbFrVjD7JkFrO
HtBIHop3yG/70jjozL6c/weh37XaFYxCl/b/ay7HUai8J6o973RbqkbFWzKR8Nfj
F5dCeyMqvb75Co4tcMu9pP1Ha0T6tupQzD77A/7fImMHQO/oPGu6Ejn+SFCpd4Ja
1o/9JcNwDyCRmGdAXBb3Lb/Iw7dN+A2vCCKZKro1xFIY4A2DJpp22Fq9YBmA/3bC
ERGLviNkZ7rk9iopq91bVucehPiAJQEA6pomNvFLXinMx5s2goso0YtoY9sqse/Z
fS2Gg7IxlJ0U4WxIz1VtpYvPw6KxTGsI1EwMIvyseIO9pGB6Seo/zWQbvFvhS7OI
4sJ+J+vBYb1PPMfW4VWG/XInGrYHfcJYw2lZAQtbsCrfgCtTXugCYePihxCDuvcS
LLGSIa6BdIAGGZ9Rs7tHPRG4IOHjeeNSM39D25THbj0QZqokzqmBEWjT571nTWfY
Y0O9xa+FEOax7gkzAaVjYrXLkRXLQJ1VheLLKOQw9Mwi2FBpD0+rxA8eT63oNo8B
PCA1K+YZdzFQSf4TheZbORnzf6VyaVGBM5HtSku4YMmpxnTeofOA+dBpGzVc779H
LL9/nlozl0wUHC2+NnIulWOKyOpvOVMlDI1Lj1g4YTJpzQsaRNxi8bz53kj5z8yw
uvJqTdareugwiM+j/TSV0tta3FvabkwahuV2w24KI18ZG7Rlc5ZiuXA06JGuqVHx
j3H8aIU/hCoC0pdPdfSE9+SW9NSLo5Yj2V9EfUIWWBv6TcVe3hiubbB00XSUxMJa
Qu6qN49obsmcS7xmwYMiUn+XDCHfLAR+kx0/hDrwePDaCQsFcPwZdVRE55ekhxeX
3XoXI8qOq+ZDoWJ6v6+Pnfkju01CYMRkBIBQTX5KngoaAXqdtiAwOD0trI1oFqOL
C2paU6rzK3HPKYcGtzCrdZbMy3aNizi2wX4wgj46OHiVxeAFqy8COD2pxK/Py+FM
vzZaozrDw2VSqyZmpqgaTSSZyq6apT3zmPRGPx7awWjfoQaMfUBJQ2Ux56XbOUFf
suHlPRB2LOEVp+HZA3QWI+wLHJsVqFoedTfTS4dn6kETzCjA9MTU3droSpZwoXmO
S3xfdRpy2fTQBA1txQ+SqVwE15OUUUKN/8gENBnvNtJO2IsTECQYI5NgMfBPqgBE
sF5hBMS5l73dZ4oa9W8OffFDzqASlo0EpO/2sPw7FUZhnqSOQpyyvv45ECu96kKR
3YFEpYe3IwUs2KRHcAAi0Hsxl1VTzFCtGvIsFWZIguF+OULvdJZ6fcjRxOzIgsIN
s95w1Nu1+Kxid6q8DY2eKX610Ud4GwuVAUNKmGmnR/uHCX4wdhoQDr6KtB3pMKcY
3mSd+GwCJwhDSZSn89CJMHLXFZSoCu8O60aCzCqKlATZnANiLVG05L6Gr1U6JxNC
gsA4K1sY0FL7oXmoKLn98uTnycRZJ7Ek+s6RJd5jrebqIao7keHEpHmpEG6KzfFe
qA9GIebLsGuCYRxGaN8VKwFXK+MbNTx9IN2GmQZlO3L1igNTapKJjY3RovEEsCNM
0vvOxZ59kt7fqF2Cuc8jBUz+wQXmCxllUDtyBRxLo4bWFMN2YJhBKMhRkSgbl+zf
pNEv8rOhirYQGZNHAr5/33Ib1h+bUFCQRDE+de0RfqaFbRHChaAhFw30GQZ3oy/H
GYN1uv2Z+NrCG57z2CuPKGTOx6xVCa8g3QnE9Y19/o9bH96Lu5gJgXRt41gysSWa
EbCEiSPxZQQSDX2T87tmt4TCbkqs0IdUGWeQWhi2TKrPBSIvpT72EEBUVDtzKcMS
2KgdX/5sfsWZvU5m1Vyx/jhSE348OKrxcPFR0mlodo4xRLfATqev/HLzdImhZLTS
Toqdj46A5/2PBv2AyLFvvOk3ufa9tM0RtONNMrXkHB025Ue4tVURsKhDH1FLisE6
LVISAieE7Fdc/0JN4pv012JxZgLYwogPu2bSKcQDeWoRVYrgC8NToye/2HVyi2Wf
A3bqrxqnp4Xah3auMx6GGmS+LPbuUsIzQ74DAjp9sAPHy3AotZBjou3clHvI4AJK
KwYXySAR5MgwlE2hlZOa9Fx78O3A9+JKBpT5RPiA7blS13lTe30cBCehHemcnJ+u
ndFlahDMNnazPMIG4njHlenvCDn0tBva4ibEtLQX1yigY/hgwmY5NmUWup4hP9in
f3IbnaIvasl1x3nJk5SrdmROg6dOy21FpwvyllvowugCht0MZip972cBH/NM4uEV
PjXiY27gB+0B0kCk1KjfWyC5w5JA8DNYFK7Wl591eobi+lesbQXUPdRqdd08Vqsb
0JQEpy97pxfNGR7c0L/HxeQC5PwXZ0BAusUTzzbE7yesetSydN0m+hqdOrPqoVip
4/f5ZsQNTPYeJcEnd4uxS+YebAuAxG7/WR3zn9LH0NLAhnFfCvU86XrQfzARJBmG
lBg1WA56gbgaTdPHe4Sb0OjtjbXvJcVbKVmD30OVF5putMv7k9oq1qX+0gSJhBCH
pnnnsSUkdySkpXFSCCkJL92fDmrBs0cOY0GHbZJbS+fLAZpyLL7S43X2niB4Vm9W
kyuZ3xnv3DJZmh0oMyHPmyOK+yriWxlIClDqC8DoxwQrptOzxGuM2hu8fPV7CJkK
YeLsAvi93TA8vh5gfXDwwEOhSPf80MuLluxu/husZNSEfeuSxfPIFOz3TPoPejsi
Nz6dFdaruxr4JJLPS12nx85kRZK9seU15KxdNA1ZzlQvF6fHLy+MDpYo7qJ6kWMw
DR6fVlIx/1wyzF7grex1hHim5IgkG214oap7zy+QzktxHO3EBkVdZX1FSCwYwbll
L0EXSnlIEjcwz8gHq+WfeEqyDx2Jmep3LqdX9a12AuBr/QBKBuMXdHeiz7jocq7I
6kePbm6z/9sktJKXBR7fdpXMC5fN9BP7L/TTGayyvz5NrTV9XXQM/8h1eApDw7Tr
F/zhOnGd9ethNvBryuZXrbojggrbUlvR0AcIWboUIYSBGDUL5m6ULpElxj+HEw5k
sZwVtc/t2YPdob534FKb+JVG10zKi4+KIBPVG79p+maxXpiHD8I4T7HtS3Hm7pl8
H2nL6zpx1K3tNTHClJ9a2E7KNaqcJBvLVdNOmbEZjA44TzLkIosFQ4B/GwxNeZ7s
VS22QnJ4V1LxWKJWqIlkEeBg8KxQl8mpWidgrypHhTnFUFNg4T0XmD4rRxIwCvNG
V7+5u+SFHAz1IFIhdrR0t8LMSwsdEvhNkCdUEwe44rFZXR/GAErJ/bnknflbyJHe
IME6ZqZyzA3AAS4wMPd0tLjxEKBvi9OSI5LVixiHovEIRFUiwl5yWeRkXZyTEVxt
LquGrR0n5zlrBcUkzCtABkfggkSmwkefOsWUy6iWckcKxr0zvuJxBRIvJvbEowp+
oBil4+gIXw3YmhaXyKIq0bHJbdiuCQX0gal6AaoVKzRPlJzGqnOj27pNKheOzUps
fJI6x+NZCg1seofQO9gBv/e5Yh2EtvxvlVKxztMMp/T1o91xgHmOtdIwjfu8Xrbr
ajdewCdVqF1pSEprYVdr5KEUoydogDWW5riSuKca/mGKpWEymT9t6oTzZF7VmKSm
qRd4g60i/Z3G0JQCAtYv+kBSE4g+B3ikxhpt/Ys996nxjw0PoPE3U9TQelSF6i9w
EAY3gXYin7IGF/CPinJK+aoKbA3E+rd940ZRaduSk2JfhRrxArwcSZ/JOw3lEe7b
+QxyDXUKmMoZuHCk77B0arV2WMZOCbKuahyeabkwEHgNwqlJZtjIbt02vMC3SoU5
xw0MFomTAOEZ7PyADfi+X/neO5NfzHUf1AKfwt3qMbrFudIYqYfDHiR0ghoX2PGF
eWJLTuW0mfUaLE7ijjVhI3kT92Ayqi4BwV0mhCuZfwJHSVZYtIMTvzjoiVPlE2rq
x1ThrzhkjqEsdyjmVLWrMIGwMZJmUgqMX3cIr/DyPyFrXyPiz7x1oKxJEYMmbGD/
iINpYPx8In/TaY+l+9NFSj8ms/wX6ghWe3E26fj2zb/EKvQDUJPXw+cEN1Fq26yl
q+sERI+BKe8S29O7iZ/rOvugqpf2YEY8PxZe5Fh0QJQBRDhkTnVKOreZnM4jmbQx
4c46hDFcU6PZKo5gV+swra6r5ZZwFdcPfGg+rKdlPywwUE8koFsq2A6S4VPznXIa
cb4zBjMd8NpvcFDSdq5X57bOlaL7otsBHC00tZMvoaj6tIXVKVUV95ab1iK/bls7
4f+ROCKYEwQfGOmquRieY7rxAA884TYKyLYELdgWBrlQZuL7bf/Q157w7f5yDU1u
l+ytasvuth01eFp4gAnuSvzRzmkSNt5Le+k9ih1KWKuJObGV2G/967QItNe8niFz
AJBiV77AlLR96Ykvc6SqvO+yMTbhUt3IP00Z8moOtYrnDQZyVNAlXW9vgaN80dt2
9SWD2qxsiZVzNgNWMmb8tKGJcT/CfxtC9hwut8B/xeM+IwS+HUy9xp2xf56JdYJ/
3rK/qsVZDufKmmlsXTO/gwKdyQwvslYhGAj/sSw0EmMUvsU5I9CygzSOZsfIHMeg
4SOiNNQbxPlvqUuW8kxob00UWbNtg21acSw5YmkFlccyBuBUd2KXEADrXkbmA5oT
JUHGphlhtH2/g9tjfatzT2n1EO1kR7oZaBYzJYa9+cGjhc07WJLSqNPqaJZE0PyS
0ZVYtZ3bVo2tiW3ex6rqzds+jHo3qdLPOFvPv67/IwwkYpQLnL+NOqHUHIb0/8EU
b+dxUCknC1ikzSpz7j0nJJmqWl8KvU7+mkAjSfp7cvpNXzQT3ryH+n3mJ79NsjFy
tycEM2Sn6dyDWvXjhl6+WZktPBuKNybAoJvcd55fdAuXZsGLv+hHfjukZ8YKGwqt
xbBb87o2UoJr5M8UTYKOtI7K63Mj42XTvHJ+Y29X79ewm+TQ6bCCsA3XJ49f6WuC
+hDuWWXw30GU2UnZOkPmTGWJmD30GwT3FgipsGsJh+h2+uMjFiuNf6Tjtrs/S64J
AN2pggr+UNq12L0ofBEsX3Tg+gukpM7HtQ1jpd0W1WFDjRcNE6qcgTRnsJGAXjAd
5wHN2vriuKXx70GFFkeKYq4C1GO7tHW7fbuJ7AJdBmLCQGw27y7qnQdg4Uq0xdnL
a2+iyB917A/23Lm+N6SjtMTbiuFaeJQ5THyV3xHn+xQFIOn7xk4UVkgNJbruK+he
OVqIw2hNCJAWxh7klhdrjuauLLfyCm+OhfltrJIFharq02w5fK6BePC41LCjf0nl
Z/wXpEdBW9kthzRcqKl9hqz1x22gjrAJUnASLugWM5JqLeDwLHVPuIaF6HIlOb0h
1nzZlZzr5UzVGiq8Pyb5e9s1672WvORSltCVFsr7xGR0pyFDzEvOD3Ndzah8Eg2F
UBpebK+bz+w1SD95lZbfLR8Rxw1Ov/0vcDU0SYGpW7FebxXpn0TWvcYVdg1ZFxQ/
NPbP5QPU2zigKREj9e78lQjh+9ANHy0NJlBDeNvFdEKZkVnYTfMQFiKeLqIelgVH
QkxpJHGpntJZRAJdgTUDTPRWPUDNliylhEtUygYLuKU6ywHtGf2jT1eWksziojOO
97hG64+P5b3l5QHJ7KC/t7JcyLq9csAJWROg4/rk1dyLGOffUjOuXmjYO9dfV95k
r88vBT54pEMnhpunCdmG66PL6ce8CK99fN5HeSZmfqJwTbMnjfrR7BerWjA4gA04
41M83VAQU4e9VU2g0rbuAuyRqK1rKuUWVCQ7TZLbKxGkS3sJuPeHxNC2o+FRME0R
JOfea5Mvk27iRLEXVH63/saqrVeEn5TkoiNDN4+IgaM5jQixdGaL37LElsnhiA9u
O1tK0ltMzMDbWTW6vq41grIcoo7uIMlxTSlVMh/f46oHsyJnW16Vh+t7VmAEc+Et
1QfnDfrKiwedp7fKSNk/0JhUvg5P4dzfFAXCYChkEr4gJ1r6BFo9898Qy/T3f9MG
vKtmWBcU156iU0ooRFzNnQT/3d1q80NSsq7D95qU6p6eAPjzI2L0zqhyKetgXsx/
Ky/QT+t0JQygdnWJudN/3OrPG8ikoyd4Oq10RW0bIkubASLIf38oxV1nvRTJCBTG
lARrJMTGKkrrtaAv12INZHMGNZz/yNjOQQktswDQiduMljPV0YF5eOG9K1sgydPt
TyKYHJ+t+Kem/D9NGBsCRLpT++rC5DM9AaWtwglWGsjPpZN+nCbW6QWq2QPBMLBK
gc04eRjbP8PgR20kZ/1PvYuN9bEhDacx8d2UgD+oaCvpxpXdktaH3dR4BJBoVP8b
acd9lYTa2IHo6LtdE2YelWD9WQp4wnhBnTeWBbGF8odQoZc2Zslm6tdDXC9tMGJT
gVdXYW8+hAJQ4BiE+4/tAP0b1Oz4v/PesVsdG5dw7hzwtqjrK8Esj2JNNGeoBwkw
ovgyG0jkusSGozolDc7RsTWI98pcQB2iNal28Zhhd1BT8aMuEbP1oi70huyrbnZr
HzUBHBbhN7AUe5hhL+gm8SpFXnzrHx/lTHM675JO1w0WA29V8/ESqN3dBlrPwJwJ
Tgql3a6fGH0/a+CHUp54o3WtY9U4GMrUrz9qLdGzb1Cp/FzJDZkr/sn6cCRbsbSj
zzXuItiuqF8t9BSyIRDp4CxBfwRjXVVJknNHEZgTsxYJEraY411lwiPUTZEWaS9P
WLWgbIfReArpgcFkgPf+GOAsqZsO8RcNG9TiQCN7FHlj3h9/XLyJ0MmlMe7nSRMu
ZOhHlHBKPN23MmryoniqbN3YmWSC2ZS9UkLFVareLc338i6phUD6Bzmm5q99YNje
IR3/1EmwFDiRQo203LzBQdvbqBa9CV4wtXxN8lx9kWbOXCZk8/tIinB7JPn4CkZv
wmeEvbaSSGQfYIrtjLlo945Ir+UWRVQexKgp83Tzwj3bIBGvsohdwyV+5I53afk5
H0D7iY6IB2MjLfKHUT91M9CXQrZ81iPuh1IGEqSEkkbnphVE5yW8wdeb/Gah6NGR
w4AColWE7Dh0Jqg+SqcPjA1tSvb0lfw5mPRWx9yfnVQfX+23BlZTqIEgqWhNVi2o
8FxjVEEjAEN5Qm757MHejoH6TIKBEn8+GuNNXxixOyOz3T+zG+tjjkroKRHP45Ly
hMAhuau2jdHlWsrAerrlwZo1wgCQsvcIhtOThkAOP97yPqd98huNuPOdRK97at0N
yB9DWLcMIXhmFWUDncSIL/cJoXeE/smPVcK4CdG95PcrckhT3fBkOo+cBOnNtZpc
JQ4c12R9AfmNvY48UZeFF7h11qJlZ+K6hkS+tZRYMnEXE9Sh3hnBmsncVQLq2/bf
PjL5oKMkhJXZEmXiRa7llT9LO+ugsYbkI1XPtRuaGF7LiQI4dKKbN8KqCKgdWRzY
B0J6yNTxogsE+QS5In3/ZzcWMHmGdTIoIbpo1SDdpSAsbwNpbXEZqwqU6faRZcKX
majhBuSKx5n/Ugyh7NN5tgxmW5gcaVITDOHwpDpsZT70345Y0s2yA/grbxiL1p3K
WuADDvaupe0YfdTukxu5QDQXhDF+399Vkt3ZVC0+4NGmWax4rg0w4hPXvpMlpT2u
1icIYjwfYKNAQQgg0+fY4DLGC0RWwE2lchPDr/JCWqZlgJl1miEzUsid7rbS31a7
v16QR/YaFF48tFmO9YUbGL8eSiSCA6NyGmYO4vH3TSNsF8Qjom+k5ZShve8gMvEo
qi7CdsHO+HeGSErouedQsCkfw0wDpEAi3sJNZLusr1TMijPaEIANx1uAOQ3zahdK
vBl16sLM1sR8Y6GHgiMREM6SRq5TbHCEz7gDshjxpwZ0wAyaRSq7nqfD9Sv+CuNO
hKjrpHASawjGlLuK4180+RO8ZMuMD5meR4k/9Glvz7q/IAopFARbsLkSP05cOVTa
P5M+elGA+Gmcmt2hJ90pYK2wTeF2CKjuiLTg3kpabF5BXgApMs3NelcYw9WZ7kpH
DQgtQKuwcWEAWGJ86n9Wi/IDChn/eaUZ/fbZX3nCMZmStOIMSP4W4cPfDqDCzluP
5jdopYARua+5J6ibdBvXbPLfxEqGEZwRjRDeOD4X4EmVL/+8oaY7hwu1w/K/8DbE
NzUHDBEeRkY6S+Wshg6uN7vsWoOqv+aLgMriwelNKl8hBfOdHTh7GCRpv/3Gqrf8
v10C9RRBLWfGQt7/NqKgFWuUK7RxLqHh2EItHGbq04q41ACKSNwWFV0D4yLmgDVK
BK0ZqDg2/EDnB66Sq52vfobUu9UiNL6VDvl0HmqUmjwsGKglkf6bMPaGEWxtUGcI
2GuDp3UpENOEA3c0EOvm3asP3aC3m0kYz2lA0CnboKXU00p0fKkQTqAKDKC4Egkn
Qmxe5l17Elqhd9MJrKPYRVnRpCh2i6N0h5w/GAvJNbC7ZMUFAMD7BICv26yYPJJi
CQ2hh2KNfF670jRXP1bTVflfJo5Q8480OK0umpfRqrfXdpU96yP6/ZAls1s0mna7
gA6xdsGPiIcfz98pnqVr2tOk67aojcLBI8hc34PQiLEw+iEnR4Tn7RzaIur7yZJ0
zyc0tNobe+TWs9hJOqG6ei6zFm61dfwMDOziU+2CRvb3ZFjT5j9dCSSZm0ZOLzBS
T9z4Xt8dB3Uw+BVxVF2RIXD0a6ftFsFYDvdS9azqHqZqPntakCj4CYPv0fuyGZEY
sjTifmtSSePiSKOTs+vRtiG4jL8NedHM51LZSHag5TLWx1bqyu/W/w0Uj2QCtcdC
G1CuXp/2oK0QsG/n79FVmhju4Lluqk5YQMGuJEWtRc9moEcEMpjZQe6kb+/lHeBI
nInVh2wWKL9LPET+C8e3BoVNbZPBzlu+pCDN8hsrxoxfyyh6Jyn4lohUkMLjSQce
JOBwVXnT27wTEXgcibn5dcNQGEVZ/4yOrxX5HI4IItwkA04z7Yn1Gf2zTzvLPpbr
yyQxg/NAHISy0QNwZKgL6mWjDQEcBgDKqlaO7pAShOjOV7F+aUhGpu6m8AvHUFFY
Bb8MtlFZ6QWEjacDVGznuThH45UZ0gr1VU4ckohN2YHZ2ybkBJgkoMFrJJSem9J7
9mbimEOrn20d5G2QZXVTIbu1gDw8MKmm2br9d6938xol4vrJJLKziyognGHaxp70
BbF1jKKLRUJIdjKMmMe58/GrGFT8gVfSs+tz9imIX+A5JAh+Ue3zHjMfev5DA9yQ
OuW/Xn6pTQawz8ZXQrhzv5DwHhG4bkF0fhFATkecQ2s47GFK67AMef3akELocffW
HxC6D8dPt1xQUplcKkrMvAEvv2jQx89QcUZWZvhQqwFGm45yQeLtigPYXsstUBI3
1dbc19RqttAaJ/DF24moG2PJivEEwdGDT76XmYBKU6wyxzy5MdTs5MCs4WD9Lyk/
DiownwarBjc6hXYZOAGDKFZJfxQhc0w2KNzZ9y7lua4ZFF216dzbHb6CicDEtgcE
yFjmASCj78Cya082MeG76dd1pyFUCkmV6Fc4F3h6OOBTF+cOnQV9a6m+e/POKwSg
qqcxj+6z0R2hhQgH2zc0AcJPv9blVXc3B62TC4Y7bTthMh6jMWwI0AjI8NnxqgHr
hgqJ5Fpj/XA69nN79oyPtU8h5i3B2NtM2CJ/3cyfvcy+5HaWc/7VINZQmis2mtyb
tBHDDcy4gx1gyRhIf/sQUNkjFKnliwAJSjHWVyvL/PR3xhMHXtYJ3Tzw8XTf1XVx
AWJUJdwYYiyA3Bid82lkFFaBw7BMfbD5XyoAC+T4/WivJ3rHL4cWuASgpcy1G0JI
f2Tuen49xyPRGpPd1GIhtWCAWrsa0b/PJTD6mVcr/DTnFbP//LMeFXjAHi7i9WaX
fwxRn5PBibB6YD/pcKmBbZTglQ6oQF9SXnMhSTT5mgFi/eLZ0BaoMrDoDKOJEcWb
TfBimliAjgP0EjKJguGw7h1mlIuPzL0395bwv9FgdLes/aKnt24oW1LIXv4Z0DWh
d5ZuG2zid+rYPPazL03vTdmlt1L8SaGE8ln1UbyJC0vmG8GGhPF61Kbe2rWOT6M4
N0VtdTywM9yLcZ+Uyc4Lrt2v2sUFbZ6xNL2Zt31GSymLBJ4M7kuBspwlemMQbets
Iu6ZHLGCjsVUD9hT0wDc+1tU/7vB/VNdgrVgTD3tNQsCc1CfZFNrNCXOh6Dnk/GD
/Ejb+bePi/3NbdZpq5Pmvu4ptiHpNh+thTgikELwkUH28F16ptulAhxy1kjCcQzW
6dU8qOBx2wTLGzERPqRMCMCBxXKti9m4638RpNcpAo3d++VGIV81P5v+ezWtnjGa
BnoYkAlTI5l8E4VzdtH08+/YjTghojtI4GXvzzfgtlnafy020+sRmAS8jLZjAIWs
yLtB292fPBXXMtdIFHDmgbWRBVzeJnUeCfZVNzjtmJ4rRAZ/LDXf4Walf70HgMTw
ARnWqkm60qI51SlskuyuELCSutNri0QjLDErCfaYKApOebItfDG7Ia/tdlld7Eii
SlQlcK2aNQRJoINNpBsy7SMI4aKkorSekmGVyyil3wjZl7H8ZYs6nXbBgl/Qwx6s
G/gdolyqihLu+epWz13pDnun8uXol3Kyiz9g6IXP/UnNuXFtI3xpMrhf6zxxcx8g
D6QbvZopVW8C7Bvsoeo9q59qqj1A/LEl7PzmV2S3DEOY3ajMzyQPC6RQCi/0irfz
9kX2AyXlAIHxteOMeZE6+J1Wpv5FJvxZ1NLX82hR9GA7grs1ac1ayjpEK3fwHYbo
cHECcDZAGwXPQs4shQVA7xZfY+9Qf8d2HTIRIxR5ABi8aZ5uAL2DMi3GhwHfcmr9
tUKJLN/R5xGjb+gqk1POrt7N2avWcdDXztoElkMvLTMeq46JtjGZH4SSg2IGrApZ
+zZyyiNeyf8GebL8quYVLE8+Y2aLQ+GXLmaaCemDJsg+g75pKf6/3oCRGaeUHjIM
b/6vjRWHmE1ujUxo851PyTifq5a9pHptXAIgcYFvMN5NYtzYmmKs3XmLiJ2yf5Iq
4+oR2IHrnK60hYrnK56LGJe4cHE2jfWKSHoaHaNpQk1gSmRwNyVpNr/BI9BtT1if
p12p4jG6uH02vkeYib3aIrbnDuIkwjMuYCpxdGcPv6MTy1uicJsn0WJU9XteMWVY
JsvIMaiuA0P/UaQ138ZXFzaavjnweiangXa6bTyiKv6dCVs+DB5fVhmhbBbZWH5L
2c3q9+s41avqupKH2CSvNHQ8pfsz9KGAMWAAHLwXPEY9mK9FywLeVkMErc8Ry3GQ
v2ZO13wtEXIoE2CawA3c03NWS4sFhXVWyEiRw071f1a3HSLp7vh6OtDNO/YPDvVJ
e9RTw5JJCkZygV53osnOD+Hxd72iz9/WtwVpYcY7vHYNwN526WeWeY5hqyVzn7P9
7SJOVgQQcn9hdhnUYePsjTVy4knuErrMNRmenK0mfC8OULTrJjjfiNkuh30iFo6E
JlhoZVWP2OdSXGcN59G+7XDkFc85a56IYKgbxzNEHu+G0QcGqdckhoHd4D2C8va8
oOBe4PdszF2Z/j90pn+fkHgPPr1SAQHnctuU54S1KiRybOuuamfLkPikCmSxx97r
7b/uAA4SCASLoqoDFPzsHB34QIYjUp23kPctfcwo24G/VRdpuyC2UZsaKGrQHTt2
Ms5AAghSxMzBMKDaELPOhLsUGcCZ+t7yQ/eF9IhomjzFC0ocYtyF41f5/7Z+EDoh
ahGE9eMmMttbwum+/8R8ZtsfuguKrkQ2/mEb0/EQ8Bq7f1NweWSXNfJEFsEMxdcP
kVXAYE50H/hsqzB19bvQgIQgzkPdIphZfdW973Da9MCDSLk+HV4qoLELAzGG5EgO
GuJ4yvqoTeERbwqZsSwlf3m+P0bYu2wLKAQ61zjGlK7ta5jjjDQnfkJLiHKOnnnk
s4YQk3GPcHCNIRjFrJEYBXzEJ3pNAS+YBak66ya6wKS0Bs71CsDlBMbprUGZAInl
9bF0qRw8RlqzVIg+VFU5XPNXtt4Vr8G3jC03UNxxz4BYMHbOb5s5s/No3hUVjARz
dw1/LOHqeOdsVJyfzS9UBm/jCMdLiqGN36NNhiCjFOCCk0IIAIBIrH7o7YHGFCyn
EQDUXDyTu7AC4Oeh/StDZ1w2/5doqEktv3Qicx0aHyqeZDH2J3+8Sa1XXfdir91I
MmtJVNBnaLlSVtkIdW76bZp7lM77BwRpFNRNZ9W2rVYCXdP9Mw/dcCG5PKDR/Rur
tq8K9q9RWXodp0x5rcfaas5dTGhbvelarj7j6m5u2wIJ+P+E3HhA9QPoDO83xCXm
0pTjCCIbX8TBpt0PTvzRJaLY5yPz03919JQj9TDb4njPo2u/b6jC9KGCmr5VonAA
Q0vnLIttBuH/QvqllCEq0Xrv9kAoJtnW+wOC5g+dNr9tfQQbL4MiWhgDgOQHElZj
sNjVwErVyp3pov3LYbLUtcIdvM6GXlC1h+VxRw/WpFLkMwH0L2pGl6ecJ0kfReS7
7Q87adzEGoT6WzwPcz2zp6aZVMiWyLIqdQ6G2EIv66oWf1VRcG2Zm7DvEaY4r63E
1Lmtz0IbJYtewSZdWj59vi1FLJbKK7CiUMTDU+FY7zn8geIjfmqxan0mAyMfUklx
BSjhlUjSOol0PIlW1AcsSG89C1dSZs6VXxQ/cNss44JChZZY1x85VuXA2Mf3121O
fI2h/lliZkO9udXxyPEmyFh1D8eQZ/pdWwj5QWnH4IbTy2BDhKL5c3wKj7RwBJkJ
Yfx8rsofiXuhoce/GLQghmcpKj7n5UEakHGpE0FGIwBleYoLLvI/152/zAMrslpe
d7yvlWqrb3mvinLyMQvGxSppxsiEQZcYIS+2NsqyFCHTD4wDNy06iPX6hXQzXe+a
37C4OvXCKDFIuqQGKBe9WCtYvQ0Jd7w3z8cqYayrdvddF7xI4mXYAWBag4ejFnHZ
U1iYM7HOkpyjECqsjDFdpaYhRmR6/yP3VRilQiWwfJWHR1IMDGfbAb+c1eHzQvHz
YGUD9RoloKmvFKNPcnwCBV7hgWu6V/MWFQJyMrDO7/wXiSAehtBo84g17HfZPjLE
hrtpdrHCp0O1T8GLASrZ/4zsyt4pnU9ikJsT9q6pEYI1hqjmxnzvP9QrAUnrJ4T/
fFLpFhNliiWHRVVzPUBweIC7Y/2vIeyw8OnhBexy6gvrCkx3YGSZacSR0hQQd3kU
hFuoUJeESK5D1NLBhEL27RiYSabBADLz3Doe51WNi8lu7e0UhEqAyDFSwvnkCpwZ
mQKF+shGqMAc4NZtdJefaCrpauDTnRRpGZE5bz+q6LepkaRRqGSzRFVDDzsuZD+Y
ioGG+M/WKhZA+I9C/eykE5XdnrsRrzy3Fycldse2uXPr2qawUv7Jqg3VBeZsbMVY
39K4pYw6tDA/cDVitnfMf+CNPpoPcy/SddXR3UFl5y8qRvajJG7pRf8TPdEG7fyi
KnH+w91HVzrcmd9MRNcqqxSE2uda/H1UU4HcmLAB8eA1uOfaWlui3ut2qLSeYPT3
PUsQ2AjAApFvTc6NivanxcqhpKLh7hMlAk4HzjsSHbh/fAEWFqRz5vFqaPLEWAVL
SG9yPkrmWo2C+rkVtaR7aid04GNE9CxznUwheGu8pxGTsZ/C8TSUQmLM1s4SoPJO
tfsiIlbypK+xvaTIY8/rRg0sU/no6EiruFs+44zN7CSdQDdDXX8bY6DWJ8SNTxlL
Mw2HjQcnhEx4Io5T0v1WOrN82gfJ2CECT3KhYH/5uJZGWlxkkDzJi60c9Rh7eWvD
p8xiKFtHlIWqllwyew8CUYx/1HpUrZhkH8TIATP2MhO+UTW05+wY7wNP9KhbVorZ
8G8WYZWXdKIdp0g18TpIYKg00r/CPR2kMUFS4WG2xL98cL3E9/YOYlxQ7ghahmir
5VPKrZRn9TIKVMKNEyZo/I6uZdTtvgMlv3a7dl0kjWSBndDsn4a/TmVeauIwgEqs
cQEisAdWpBOZpT1Ei+Fw3ZdjzTeAiauGUKfNCTb/Kr4ir5xE9r7QjwHXv9MB3b0K
pPTYawyq/8J+gAyzQnEdryWaHD3Nx+cTg1o0kYu5zLp5KeNPkhItYSEM9F2gmT5N
H/TqwYUc42pazDmO6iLhME4oZPG0MhCUyJI//i0dD33Ac62QOmNyJg8b6bdg4gEw
YPKlyitjnH9MOz3Qqf01LRA/wPvfBQEVreTkNH3ksNy/sZmj/h1yoaCCmbsKlbTk
rcB90e6vxM5DjQon86yC1STXGybY6v4nbQJQLGg/0ds0w4OR4FqPqdAdrqlWk6Fz
EQPnxiYs8gMBxhkw27xjOFVNhgG0oh5WA4a+p91hCK8gRCY/LIbq4sghj5JMO6Xv
ujt8ElZD6cGb5oJJFShp8NCpRhem29dPBDaJcfAhSDZyZcLhGCOXVIGNtOZ44t30
NnauCEebZgqyPtQPxsQZXZT9QX01HoGDFAPNwgdzBWOvY3Y6qdCWnm3KPbdvu7oE
mXoFxJwledOIWnkgG4COU+PaiUqyliuiOSFcqN2daRp5dJxWRdR2qbRWzEUPXUua
knIpXvGJPQqVyCLeI37qwKdlUH37plXEB1647cUVHf0996Ln5PdlyF+59D5H9gs9
N1L3C9Ta2rDB+JSVqwuLN8Oe/0WPeDojfzis0GImy3j+NXzXh8UeIUsDdMgMjTbm
6ivKwVHXqDH//5HCTwG/OFBF+L6qT5evicXw12+5DiaEYvNdavhx0C5qgVegoq9N
mUzmWYm0CvcX08SrExTtr60WrVImwkNa1LNuDBzS5HRH4l1AR1wEoxVP0nfj3HQn
w/5Gq/XSD+0w/1Ymj+1anYMqMAu4A3xV7JwhSg2FlIoQ1t5cma6khDl22OdgnonK
hUUVLWTqOcr7i8MFzNn0dp5MSeulzca3qSvkRLzSRgggzokBcFM3U3XpoLUfc+4A
IzAIWhMBvoc+/Ir7Nda4H3NJGnb9xPwVIRuUrihDQlZLum2aM4qF5k5fKYBVdJbH
j4Opr9N/Fx/qRUOq2k+VqrbQUHEjUWa4nMK6KiZ0eVVxMbhY2me1hj/mTbOegbn2
lZc+4+fxOOxjYUnTwVqxtQgWyqoVHMtQ25w/6yTP5i5duClULNWvgveC55rZMJtA
qk7k8MBzkwG2/J0lFPrYM7+yM8TZ//TeIkBQQnHhHDZ0XI68UnIyiZeWSvrIGAC7
p+8V0CqXqSj4c5RGQ7rubztngTXsTxU0k7ZsYtI2YPl4OSFiRgoNAGqWgvlqQIjw
w9Hm2Ykd15nEE4AC5HvLQrLSxdDa8DxoGqIkR5irli4+mQEfTwvIkPrIXS/nUv2k
gtwIf+m1QItiXhd0+47lJu2Kb/zz9gZkvW0oUGhbNoz6xWfpNcZ3jnCNYfVary45
aRnh+K31f6JmHp5n6P7Ps1t3Lwqg25RLwEWWHQ4i9W1/hddTC40Bbna+Ql7vCOvA
nkoJ3FxSo6WsybXScXke8LbrSwGkonuh8kR3ffbgEENRVNoykKzRpWE6/9HRCfpe
UHqMtJpYeR6xqLZcNOWAvZFBtHMJYFX1OX1evBZMYfdjopBOkCuSqbTSY0tIog3T
UPpS1r13ZXxQ1QarQE9gVZdFXZweVvhOmaKw2fWQ0xd6WJFlkvqJnuGyd4KC1w22
yAHEcajqUCYYQYl7F5j/DutET4tVcKQfHVSTTUJbrBsExehcCFcnJQMvvGatnuZ/
MXwIerONx6cUHL4Y4yFYM8BS9oK5YtyyXv3kMFWs6sO3FwMwgCA43RnpbtAl8Awc
S3LRUlGmCWI8JGzCVG0RgdgCYmD4vWp4wnl0B1J838Ge9V94wIIzPa3OhWfqvVho
AgTjiURV4JHii3DxSVSbczsR0fDELGm0VM9N4K8LOUsoZnrOliOlPQY7/GZo7xuM
Q7N/d8lPtDPwJrr9d+uQfin6SQpWKUDFw0M/5XKVD17RdofMBiu6dXBRP9nS2z7I
0Sye0nnG3DD/1VmCK0oS+g9ceuwlmVxfp1kOEPuk8EJf24kM9smi3BFLonmlRnqo
oTwrxdm/lyRDz2swSEjm87eoQM6jrCIBLTdqXfZ1G4AtIW/oJLPb0F0L5LYie2l4
euzeE37uIUqCx5cWafKA1vx0KCTopH1IHM+0ImJ3X1WTK+wpMZowTTXaSn5hAQBA
NsfCW1nTbEVAxnFmcanwlKCo+I9UbTnMNapNvD+YcC63wl6T6IPfzZE1dI9ndRXx
9uxoLNKeSyBysm+vz8e8VYNhFhmJMRlcRG2p5dkGCxK/6Ya93NHHO5FKUjM671En
obK0jqpj1pTUPOyXje/RPL2oEWRwbyst0kNBMRtESwFNPLUv1k9PkwEaPBnylfQP
BwQ7J1uesZMyUtCWJiLuactOyn+m3OEF/EHjw3fG0OAygMRUcM4TLiaq60kfGg82
rrF4sVsYfZB+Jn9Xqxov7o1Swh834eNmza40aJShhk15aB3jhtroi2FPdvb1LHJY
Zmh8k7QLm9Zxs8VXXxeeFxl2IUyLKsR4ElVhkoVQm8hOahUGBgEB6g11/ohsYO5b
tZe7TqPcKOUty6Ks7NSLJub3wDTKp8EJU1B86v0vXyZ4sBuJu7VO4kO/lcUQ6aOw
YDHpq6CDe2h5CGJKtWtVhSH2zURjkhdLpFpoPObk3Yf6SX+cwMJcXAZ2hGTUlgww
GiQEMcIjx4CYiVDakf/r6tfHsfjV9tSKNZIwa9qcM2EnFRnL5WYa3HpIINGehYWG
oIWPGaN7VIXYXMIP4OEQv/7jv+BrHgnX1Fg0mUdqCRlilqONUJiNSp229lIBrz64
xWLRDsdv4C13S9t4BpcsoAS/oTzdx+4m02CI1WY3axIdyfJrq8JH1qTcn0OkyCuU
fx00jcObW9NKnLHq/EO4I/Fdtid4e79PhKnWbJvj9RmWEZwIJFohf/Wqsyf5+ATM
nLPjFZVR8lOresNpVeak83s99jtn4F+vy+tZN51F24sBpJfsQ/1eOtLWcl4NY8Rq
O2Unf70Q8Xux4Rhih9an/N0eFi9RNB1WFw//0uSehmcor9+YRgVsvXxI9PxG3Jji
aEWFUrrqZY/HL5RyLk58wH3jrwW7lVc5M2AHHLern1/exca4fJ5sQEYBwP17nhJb
ovOWihnGuqIdOX/MGpBmZPQKSAbM3d2P/Wp59xoLyLjPcclMGfkfcV+ozhPBX1HQ
zUkhFCcTIZ43l6IFGn60I3hXMFWfLsiP5OrN/j/tY97NZvWO9lXyZp0CmshEM+j9
zhGxmuZ7+vdRZrglkRutsNiDnL9VrxU+hd+C9hYEmwsplTHgsXNXhIqlIdThgUhf
Yc8AuqMpndbivmQQIkkzJ3VcxMZYRATQL2rKFVAmE+rM6izeK7NnLmHutGFX4392
lX6tFmEzAJl7MPNx3dHdC/PLBxdBE++tbN9g8A/YVAXWQ89tpHK3l4x/rCi9+/fF
PL3rfVt6H26S+IX2hq/SsG0C7rNRtVzkffn7JADVsEH0lAJVLPn5sgt6XFPu4L7m
6c6L/w0c3y+kq+sp3O5MHwTz+rNzq4rxmErGc18gnZwbyNfBOwbSmFcIbJdpmabq
bjfpqP6EBa34zquFGRTBH7WWsgSwpTBYD+MxDNuE+CLY+Su6DnrSumNYgw6nFGmR
rsZv7cz5fvVeudVSU3XjpGi1nVTLAHPnX2FrXuEba2usOMxMGrIzzWh599vewiWy
2GOnicbLrgp01DXxdFjsBlKu9MZN0peaf43+rTNxYHe8QtYolSoiDGdRvgHJF9Aa
q4n+21uSIKZrNonm7nSX6R4MyWMYSx6lKtp3301mE/1wUR1sM+W4PttFbkLMDg3x
2VxvEchHXQZd5XDB2j24DbHfWalR1JXYN9fA1R+7qOC66ny+pf2Wm3plD4hAE4yw
AqA2T872eeZCTxKTv9QTeNGv4sUMUWqxe/aX3r7bP/LABTK4RVmyo0OXxKHpgUzV
3yBL2tpe0OLdDc5oGELHGFABduntrHFufZa2Mm5qgm5kPU6cxQ6YIO82ezYHqRvO
QXCLaP7ovAOtplLxJmW8yZR9R54vEEohgZtfe9J0eGb1TsFj0ZzbTXFefn1fzaRZ
tlTxoJXKjyqPG1SGejd1LgwFhXrGyh5L7h8E20G2624lHieH5+qXCGzysWCDdnoH
erdod2eujXekEpxO5O1r0YF9Gyo3NlrR1xYZspwf0ObD2EKHwtqRzOPxExfk+nHN
4O77FdavwHcs20MbGuFSZJJ/f9J/R/puVxoHe8YXmIHbhDCzcLBPp8B3yVBcn0h9
8ff/dTDcxRUBEkAY94IE3rD02eWp3Wwz4BJ02xg4biNAf+SKmcuRtZAHFWw+eimI
8WoKklRH2BQBVEZ7i3xs5RsseoQK+JOwURi3vBLNRASjSBziakdSIXh5d74pfOnq
uwfKal1b4yvoA0/ngJHN7ty/dvvDCHktm4vG7GiPLK20ZymFq2CZGl88+jFdzIQ/
wvnSYFQQ7tTQasmiouwqFioWoW7Mw5ddznBxh5Q5luvUDXIcLTdh24QJT1F0tg8c
j43qpmBTGrWGYLi6+LVs/FNPD8eohp5vRZ3moM/jZXQm+Bw+Acx5h6thQNxjKaMH
Z3Y4qjGiTJhxX7QtZKnOPIK824BJsWVqL0qilgQjcgYX/Z8ts7m1MRd2MNtKoGkE
FdSgkC28G1HDIyrRFgSuhMDc/krAEmygB/gbTv7jMcpQCwUTY0nmt4q6FJbBzIeR
MCTsMJNFHtuWDSbL8ZYcKvFWxLBXsclm45r+dLBn/4Hyg/ZRDbfhVW3iL8pFP4qt
1ortoytoG7ggyI1A+YvMeLRy4NzRjBprEBOiyJG0GyryeQbvslqbQGLN1SIt4akY
faqkq3xT82eTHBXrVYMc+aaAY8dBtW9jKk8xYxRgY5OJtwVonLqxXg1zgRdO/YZT
BYuV773Z/6dB0COiF56LsuCUeMMXwsrH3qMFmJU6DjsKJDqXTbULgSQ+4e76oSqN
GhxuWyZ73DGRr3Gt8pT6R8IVXE7eUdb9dOzExGACiZOufmu+ZPeVlbJR/O+nRa07
2LGmzVRHCXBklnlVoeyfuGZR1/7dq8tVWHLtGdQ69JkHFGYqDFwGDbJp7Hwq/Qbg
ptPzrpVuRmhBF1gGYtkwfWwQH+zUPf9NS6g8d705lK+Sbv49PLBVM2kv8pcNy0Tq
UH71R/WvqkBxrzhXxlC34DQraeOXuk69hSU/gx3NUXF1WxZ1pO0a6zW0vBcAEads
sRAjaGYUL7KAn/GkRPd+jjOUXOVkdSt6NQV0xeUptDlcEduQDX7gJ48YnzcOSV4d
plI5ImOFa5Aj1pJadnceIptfEtYnnZMNko11vbU4lNAWAXPSPGDO6dxXrI9HxDUC
DQ+8l0fkPz/L15lXYe7TfDgkwZoxSKHHTQN1ukebvJiDERQi9F/V3yUv4bymW9hL
pRkF7LEjFn+AzTkj5luxHrjAf23co40gSn/0vnbgtuT9Fu3qwTM4XsE3tez3nnWm
/UJbn23F+3BcwFHCDHpugsMqts5XW0KJXHbtBXxm56bOYgsRxtpyjzAx/4vhrpi4
DaPZCRYCs+JEauAIIhBOPg89OOFPFP389DZh97Dw9s//WptUflN9VoX8PO/SX59s
zgXumGRziElQxk+nDtkkmcpi4QapPI/eN8XEHPbunClsssz2GVulorItvlSXIAYp
o8Is1128+BG9RJy0QXCOcM9CR1kPq3fhXvwaQA4KdS+OvUdw9ah5VDL7UwrjYNFP
Ncqlrr2zJR0O8CCn9LBICxppZ9TMCPvkPt8mXQYPPIRJuUN8kzQyq9gNTCO4bk3Y
O0hZo7joOkLiFqmCz9uGAc4kDV6npnrvJ8+7pTyTokRVY9W59sPikF8DTC9dfhEF
Ww/r4N/1zZs1hEZzu3jVtyIcS6GgKk51y+oQjk7C+ENNzZqAVphoSnDJUWw36RUx
sZ14ZWkByMNfnnidSzc1yxDmMt68WUDtR6OJtfSxOs2lZMO4tVfiMVpNgJv1U8it
/mbyfj5LeR+pEphVU2+UsHDen0CFxa24LYnP5ZDckRzMGDV4Npl9w9QnFd8lW81A
V1b6FqLx5ZevLR039vg2Fk1UrZvT2rmLsFlEKouZjesxg7+t5FJiRBPRuBhrf16/
CkPBa1gJhXKaHMcreQT3SYAxW3aN6fjZDTmT3V+YrSNxpchYa0N/TdEsngIiYSwy
Kd4/TGnAXgCd5hqewetHrSJ2d63AOqV1oQzbYYtx4LWwZOwToZHY0g2e7cSZg7hd
oiGIkYkaBgM7Kzu0BM2Pj3apiRBKn5LphFhpsjP8y1dlzebsJvhXIlDgZQoZA1Oj
BOV/suIewv1Ffx7ptnr/udKJ0K/cQuk1FpMr5ZEl3LJerP6LMZoltNa0whCfIwwv
8CKx3rr3kbq6Q6olsSr1Gx+nNCDnhP9xJZpNZJgnYUDuSB/XR61LOjcFZRoe8v37
95v7e8yYEDgMt09dJRAXQtfrx/10UkRLnjSyfgMS3wXIYkVbfPZ2DlMhZYIJAfuN
1cxFam1n0ipPpVfPJgkhsuk8RrbdwgJTJuuosluUBj4ecWJDiH3aZMfjRjqxd31V
6ybJCvAczxcxp9ZVEsJjstM27XjwjmhULrtv7FLZ1usPZ94XYtvBsXW0EOW74CFI
FriST6BcoF2QINXT4QsQxpofGOAxlGaAlKOqFbrnu7qzNMmhoU0xCWTN25DUq81H
YxERFs/Y66/kQLyuv0ot2Z2FA4hBp1iQBWKCGejTE3qJQcTD/WkiYaO7O6VtjubP
JDAw7Lr01mKsRkSY6w1U6BBfqVleW8fZ0GSu3uyt5x2bawNy4QLZXh6gHrgSIYEC
BqHvOuRrozsdNngC7kKP8CgU6Qa2Kuj33jFpj/vposTMSKAfyzju+Z7704NZSgy/
edO+XFMA6XYtV4WfjXkcvOiVNPVOxNmGsFzEctGwUCvTKon50Qbnbo7KVPfEaWST
034HOzjW0ggBfkIxUFlOwMG31aE+jQxeFJEdYKxPymqrpkQRLjLSbam9ZgL0ivZL
lRSbbdv4ighBc7xAJkT50hQYDr0ss5tMihz+51ifrrMc0Hg/vqwMsALrDDipuzS1
pOrWw2H/4u+qJ0mtUB5jWuAzcw4ZPloXYbuEZxKYpnYhm+x4kIjApNddvzXW/Y6u
ANRc1a03SCprcj6sAbRcL2ELbreFcBx/f041759/zElXTtlZue1nKFZO1oYgOHZt
M39aFiIYCejhHy6dTKT/FaXVACFcTdCbnyC1rHesnLvHwoCHxnCQLIZqPE17Z88c
xM+2ACAiGJRcbqjvXvSP16bLwsizDuKZBNlZx8mo8Y6mv4jKhIrgFxtA2ph/7ASI
X8nEaLcDVbt39DE87luXFXXxbeu2S9ySCHFdr2aB687f61ggsxK9EgoelPPHQvdE
RLXX7FZbEQWiyECYXnuLo5XZLwgie4SP+fTykVWN10ESK5zsGaJ8Fcs1jpQAu2Jh
FJUXwjLwqPdT3fg46OYFMoe1ZICbyjq8YV0cZ7GxjDH9fkYOElEBy2LI+fkfOQ3v
efA8z+IKXeFSYwwrYZuldfGVNyNcuRcvzWmQaytxtd3rqu8sHbiE4MgHM5UbRpyM
xJ1jKpkO5oVOnZfHlLG9zIXxktIb67LcSxai0ClXNQpqFFpeqaGNngGO4WVqKTow
0lcxS+gbtsI4aa2WJWcThXhl/PCrsXE3yaN5tZlR32IFff/FwEdS+wmMWyLLPosr
H1lX7bpLyns4JtjMhYEC7yA/D/PLAWnYaEELIlBS+cMXEINdBg668yg/PPQrVkOH
f43jMZStaewUDecUOaenGBU8c/1OIjkFhTfbjSd7qHOVfnnTq/S8S3DRyqYmhK+y
eWwPne0p2xlLXSW/vTOh4vvHSvoVX34eK10oYBIfX0saoFvWT207NpxoZ/1jYnn8
kUypAE/UeCG8FuEhpeNJ+iWxvhzS7W2HBDFcFld8HRM6HMUtxs5e4memCMoj1KOc
GKkZ/ezzLqzOylqJYZG+cARwWJsyJAkgxPw+AxbggNMRRyB5ZTS7rajEvXJbJuGV
KPqZ/ONeUx2M8YAWZfKCy9sO2QTj/I0fCb+PPcEXMOldnRH6pZQDWtAD0QPfVLVT
rjsGzpGEtnpfXmiNyY0j72Ynx42zUN1bLyUyiV4+vNprVKrEjjeJw5wESpu5QR9H
GAMAuS1jBIHLwoi1SRlkO5fJHBddYDqJj2z5EEkeZMdzgmuUm464YT9Jq6ACSXRf
YMkmEfVJBcUnsHO6WENQDC+Zgij/j17EIyAUZTfrsPh+yBhbdRkG3+HYgKuThsNk
KwoT75dNoKpWUWIiuiZMutE23wRrrdsJQIL5eeiiWJYSMRXKKLYujl7cuwjbdfR9
M6kIPR847u8zQq4cGZfA8GTm7wZlN+0/icqU5g5bJGnlQ0Jd0Jg7fshPJ2LL2wCk
A7df5wUTjQG4DwOhMLUkUhuUtgwhFlsEH4VR67+8fCRtDj+lZVO6rWx8C8G8jqaa
47YtmP/wyDYIGS6ozIykkTpoQ68yDrc6reWHkceWPxxYRHVooPbqBdfvgtONmBRY
WOmxz3fcOl04M40pw4xFhAnk6/UJSl+xcfnXFv6s7DWSTgbv4jYTZC8sMVSkfYaG
3XoDY4FJCHWTrPIqMg1JkKS15vLsKAX9NcdqcnND/rbcfs1RgP2V5VwTydXahrpw
m6QVS5mbKolGTs171hDmLdyx5haCXRxBmXYsOJSkgsAWkgyLFV3G7OvI3OZQ56Lx
M1GyRUDPZQhHFMsXrfpofprKKWFKa16OgoepYhhdSqWcB2oUE7G9NmkmcjXDu9qu
csXInN/OhXqtfVtVxRZ36BJ79A4uo/nlhH7p2T6nbkDWGwRPTy9wju2/mjvkYbG0
pF21DhvjVy/YEdGfjYIIpaml83acPbyTBtQtSU8UD4L3IpDBu7KRYXDfFN5+47+C
5wWzUuT5b314l7JGxNAQtVqF53oGoPYg5qL2ykby4zwfVMLebMMMb9xEVxaDSkfn
Kbr1hsTOACX5gPBCOKDxsJlO/EY+c9Z7Db2hn2ioiGDoyrJqDL0CKYlNFSD2xNUC
74g7kZiPktOHInQ8XP74bqgwgXim+putOYAuY2vDGY3wWhd6Xq1m8tUZbJlP+xMK
LMLwG8yPQ33avffLtorTcmujrW4XZEgtfs4+nZCLSYF6kJEipesgSi05xqXhXIEe
f/OLfOclGky6tFIRuqpZVo22uxBGWE9YIxld6IhUOBKtJQdJK6yLVxdTAPfcFz4u
/xObu4wZwwYVnirYqf3+YjKDiWEi6kOqjUSZ16joHJxcHfms0cTgtNyntEZD+Bup
oJg3dX3DR7Tf5Uv/tZt662lCed1tan36875STkb2Bs1dS77LKizB3ieFAnpPd/vv
Aduiw9wLz1TMEINbHE3Z5tPy4FE2iizGV5vOqcrFs6Qlahq5mNdpN3LjCZMNMf9i
qLNU9/CJ5yvo5U222RnGMcRjNSQ0lXYswuMajcPbxT7oXZOn3KU+/0FAk09cb2jk
hqf4BTpwdRnh5Bau+AkateQzilaqMuJjXJZVRysFx378R4TSyY+GGGBoAEPJdK8A
6avKrqeCkdzQN/SNQua3mFUmccyx9KuUL3pMcY1fezSmTSSiO5YaEF0iGqFnqv1E
4MFxrLm5vGOkmGijQnCuwzhAYHIqsmTnwSh9tlJeMdz1Apy21A9YB11nfz9Xc79o
XAHWf0FMsBkfDVWNQiAzfW97EpK4+AW6+HgnCzuTrYasi0LCbI43XH7roB4CIyj2
zgAr6CetpWKXFPbhXZ3JGNYGGN1gBgTLdSQOj8p2Tryb7cYPJvSkJJIyPZkwUxZo
SOrTcZmTFidazpCFHfDA5gLhdNZkqemAQiLq74yXN7qkKkLy+Q4yjEX6qEOAbAnc
WUb/6vgCmNPD8oCrAqu+qjEoMH1xXht/hLj/CY970QQA2o4qZl5j8unPKrxze6da
q2pcrV1GdsCI+/AKh/5LJGL3HxBFIJ6HTmR/yy/8H97vBRFXlkrC8pA9Of2SDPmw
F2LXuj8OcQoyreX6oyGaKhp1t0aHWOJQlH+DH+gDOjCaxR1jJ59sw+fJTqipeJ9F
1XsV9p+EoOeEswIr7gixd60RpFnIePoicGqZpLwzEc2kqd/R2mzFi/z0cfHcGrro
gIQdk+vIRkP/fXugTKKRQbNqFS3HKELWubf7zbLhQFYzDnZCGLOhNqi8pvoE8WmY
cZOCuC6BdjjVr9viyj2nExr69+mfWnbmb09rx5DyVRQlY9VljdZm0J3dz9TpRVDf
TWjDofkQYtwYAPGYFHuDR+0xv5vNX8onwP5+o6vWt5t4XolWPGRcBE/oeZob+qp/
Hs4FzBadvVIbeJYEEhBYId7LdC/VxRiSa9sMtiLH60Zs551YUl7Rgcvf4M6u+jb+
UkR5JVvkNvfhwa42QuZYzJ8EFYbXhfJ3Qba5nmJhYUCD8vBLxk0k7waUowz4Xtu5
n5tcbfAkiu1+4RmmvvSjUlfC0dfekZDjMnP+8NNMjvLvzaHevt3iZbWv6qT4uKsl
UGjls+tEhB9pPqqvlvJqslrFa9hnHJzQnReqVDFuJeal2QTirPD2Cw4faNiO21Ie
oswhymbr+C2ZTQbUP5lhjEdqaqMYVgm5JXDOQdwUwzsQiNGeq5tAykf6cw61udnb
jPW318gTLpo2OzObq1pRxL6Ta2GJwAzPvcF+wCldPYHrr6P73apjSF1fq1a39CeM
JOsHyn4LWI3wGmlXrXzHbG+IWJIA3GmkH9SScKIV/eNaDIV7VpLQOeGh36pP5jpi
+uD8SX0TT8W5vvnKoG0hsHowuaxPR+96J0s4Vb35+K/rqBqCPfxHDU637942Q2kj
6JwfHNjbr8kPQ1JaVExTDhanGnNluFjqeu3nzPzh/YMaR/l8L9TpMMTNR3K68LcD
w+StHIBS4sCCc3dLqWepf+Kx8FcaN4sJL9D/v4Gg1xytmnGgmZJK/2zyeGKq396B
PMajMlM17JjjZFe3LTA6KgC6WjXrZux49dcsTkBS3k3LSO6nB/6SBOifrUObwtN7
8yd5JW4moqx8RcOwg6rE87NQkhKAMCt2YiQv69Oj3TXvOU+Cab/CrrzF8q4dKjfS
yNrYuA5+F8QBmwDawaIanXbaQOUSO9rR+VUecIRzWObQkgwAJritWSm5Dn65JAb3
J/hF608Vk/Vp3r3KsWRFE40znrbbcJIRiMSYV1X7jtDxju1LMFks0lTIG9PcU7eI
n413MiWyk9bUJegp/t4q/lbnaMxwDbPcjtKB853nTEHSnCgVAb6jwt7bnVQSVAWC
oyL7+Xg6RvVSPOmVVhbVJP4JVkCTBLS2CKk24zkI4bK0MImkh5+nIs6ircFoYQS/
XGv7no7gJ+hRuAietxNATU7H0IYHqXL4Bfb5xoA1LVGdrlp7zVYdze5f72duZ6Ep
cO7HuQlTOBBz4fP/V86Tey4vkAKXFzJNMuAcnGIdwRBBn/SElTtAbkK8dXHmfPVM
6MA4kHlGs7AMo+uliAscQuvrrh1Uw/kY/QtRFPLu6ICi3UYoPFzZElVCE50sQVaG
pmkCiKfiqfVTJzvnBrfCJo57sUky/i4ktpG5uQptvcgzgkYwqAkDWmiZsqqVctrf
FQ3hm0p6CrZmvH8rxULBdFhnWZS4mULOLWBNXbNyWPug49yRWltXBG4KQTsU5G5M
Jac5eT+oT1fG2jtU1ezadYzhFWX5N0rWF3cjKjwqp+HcDch7YCWYIYuiVZFjcQPA
VqyIFQGsI9nLRvevujwCbpH22WhFc46KhcwyFzdB2pkOd4t2/api5xgN8Vl3rZP0
uBEuo+X0kova8lPKuZMOSNBfVtS0vZRXMPWr6yKThNIcVMwSr7YziOk0ultjkaGO
wBoo+FN80u+f7MvxqqbHDZdWooPSZ2x/Sk3nwkuc4wIpaqz+e+HSS9zkbT8SEdAY
z8UNYwPeL5LLrca99JCL11W0FwsI2qzadgmp6cZsCeFEJQ332N/LKULG4sztUyvY
TxHVQ5DcCyDCAcOvWhZg1gQHs9aucDiWRbbBiEQMoi36hAlapmCoiKyO1klv+GO1
qDTcEEyBluGj31pPCaIqdUzCgmI1Ht9pPBq+/6FHY9eWo5N6e84AK3N8gdqZO+NF
/WjIErjka5Tigb/usJkFMscMN0gAmvqOFs1H/btRvJ/nUsMW2xuSjEYOCe8EbuyB
fbrfA+XG3VYOj0fjiHgoiDQiOYmKp0MTlefJDALOzjrYP4YJGWEgjCsPawK+Gklo
fIqSrR2tuO+zPIjosIzJkgm/4xYYy8TD7uB9GkL9BEqxgPPyIOBv3ZoVZMHlH0v8
tRwOSgQz+/MJim1hlDEikvjeVjMIMM8cZX/yquP8dW4DLvKTgN+pbHVld6hmjmNH
T53dTHRAdn4eUqn+QXmdFgC5GU1G9U32mBYqPTpCT6/X1PcWeGRddekUmQx9/pEo
Pj3cSa0ACJR010Acmmt8nD2ngBdw84IxENfDjr/qlWPAymwPmbRQ6McLyTRbJGDr
Ws0cIubZVoEk0vjsTnvnW76hM2HVgncMObvhD6QfgAJNQbr25feY2kyJYEDVI+Ym
GFAtXLXw5BC4WeA1mYqWpCwd2MvJTQizosRCkxyZkE8h2amchDTRkVBsSKJBRk0V
efGxrK2T7ytwZVHmI2EB+L4mxM96yJTnNW8ofqTC5Ltirgh2aX6RoTKk4IMIu/Cb
4fnRf2cKbJoM361h6if5RPwJXsr9+2Gq6bkfxE1YhjUJ62qQmNJfZ8/lEAKHy6GY
b+m7UuVDZSSyikL3uGa/U32auaTvZE3CLTsbBx9InKnai4tpfQYPv/ktavwN5JKb
Qz/fyTjLsjZqHwuUkG7gJZjnoOjK5KHLCK6BTedQsyS//GtMdkg4ItbhM+mRGttY
Rafh/nHfiC4Kv8OppBkWboEX5X6MJdzCjz7uxkIZyV6jdvwD9kuJNMZpzxdkp9/O
Ng8R26g1h3X/SWBaDd1hJgQJWqNkt+2b8Kj/feNv3+kIDtShJyJ8M4fO2DG3if2M
hoaSAiwDrG+yEBiNxsdaiJmY/IAX8kOFeQyuFzb2KpLUdIO3kKuNYLXmzttBTdPK
Z4nuxNcBlXO21YvFyQndcZDcqExntuYvkgP3LS6anIvfEgDTdHlxkQcdiPmRi1oK
UKpvJlj1baWz7nyt1GjD++ypMDyX6Tm0bLQGuk9OF+2y+Lf0/BNikcYMFKib5NZx
l2ged/PtHJ7g8WbjBau9enrOC+10dFAWwqxtKUfPaU5yOXoozJdTqdu17Lh79o03
Ov0EIEDf5AMTwLft5pA6FAc0hkWejEQXsWBMkfr439o5ADvfDqTEw9VZcxHrCq3J
sC+c4MvdMaxI6eA1VgqhfliXdjfks/Q3TnwaC6TU5AHn12JS8zl8OoHsnqztNOej
L3nmV6iE7ispE2GmGeCG4R8H1ptF16WcRNgujOn+nVua3Ov1b6gC5yCRRRgm81GB
3qAh+H55H3sUCJV1P43wiFSJaZ/B9l34zrJQWaE++W2IKVkfLqUKFEd/wqTEAp+2
a+YZCP4EDSD6edJutZ3Te+eP/cb3r0DsnYG/7H+vcAOwrcwiuYwUAHiOsmETC16c
NmqqKS820hMK7QkP5JoPKS5zkajLb9VUF/F88+628mhI6RG2lD1Xz6rE0tGDP7I0
7t51tlzA/t/2P7UW7U4s5Rmatoo7zILEoL188/WvGWa0e+pfvkPuParxjcHgEIgc
5UuPnWAKcVHVKXP6mzgNSf/v0Ts0hWNOrIT6wKCeQBoTjHV48VttE5tEXq3ENUzA
ZeTej4BcF7iMWjDXQknlykGE0gKgDH7XVO2L457tLQC1ZynIt4oeS9AyJA+MBB+n
txX6Ho9G7Mdv5DYe0NiVE/ILRqmD7LDN/MH6gmCWrM3NNU1H/fD8jacgqcwNysmU
eUdWhxUwcF5gQQhhs4b0bF4WPXTxMxzDTrSpe2qAAeQA9hRDwA6KRgQmZ6JLY5X5
4PJvHe9WPyyL+KMoGkg3cE0YJvqaq2V92waebCCpLDyukfiKBZGA3LCZdo/SN8tx
b+pIUOMQ35497QfFFHVvB6Qv8fzonGw1+gdZdRe2XMH/Ie1vwlpIlq3c/bmWXg7V
8+0O1Q17M32IIRp/11JQZ1/6TkujvOIZonrxz6pMrpqFF1UbfIjJe/u7nO6tO+E+
QnwYRDNAFj+cb2UloWUjngGgR9N+enRoxkJ6cmNtxalom9cZdtr70K0ujxPTF09M
lN9zsD7RjnPW/4itMBT5nCzLdaZqqi3lQymjNoL0WxObLYV6ePQogBKutsWfDWNO
ago0V9PPqljRpj7DBi/7Q53WIgqVDy4QRWEDr9wGAG5tWbzK0BovwEebWqovxVmW
EON3PSII8bxikG38zxTcRn7j/k5ijELOrUEDfCIU+ZPklQxzaUeMDZ9IRVm/rolx
SxAl3TF7BHRApGUPnceeVK1d+l8YR6KGsdpvhMJ1t3G/Asj6wpmzbZSn6LB362xE
sdXAU+pRgAa/Ixk5EsaUyZaQBVPgVzF875EQg6NgM7KcwXzmQe3g/YTVhJVYQKWT
AD2b8sQ47iTaVl7vubAColkLl6dltv/bUwbcOsSVtKg+Du24nk8ELvAyArHJNkHg
m3NRzETTgE+Z+3Bb+LOIrMqs34rqPIYB4Uw2MjK215VH4vSiO/F2AqUco6bn0y7j
CIQQXiXyF7MoYBXM+YJimKdmH9Ojlr6IeW5SxMUMvKtLBh7y3YfSWqaB4mlT8Xs5
JMez3mG1QHOl6subp2xO9moysPu7OHRElGk+5yO5TwPw6UvzDmN0aXX5ZfKoPWRr
3mKuh1kKB8eNtbIKZZGLpVH2OeCUU/0kROVSWicL05bq3jH29McLOF2tqvMIuNa4
Fhcdutq8CGqpCmj+WUai9WPerdKrUwmNgnm8OlQzSpl7E1QCR9oCUtS9S8zuZ1tP
71FfEYXRDS+yi7EjlkNAWe4yT4U9fjjSv61qsmit+uE1OuYXwAkV9v6Ioxp2RW2/
sOIbsh37gx160QjOlat0hbbYln4TvOcEsL8UQF87JnTUf9PBnjmdOFsTODdlTCGO
j0K718Y+lfm8yTi0bphBEbgIQo2cDLujfNPtBGTYBJIHRGxZg8BVOyFdpObW73CF
UFWMvg4PIKAHbJrkUzUKzVSELUpjV2jxoZzzZd5YVY5KnmFO/kw4LBmAChP1bUf4
NXHuRb6v27WImgLp5+7agdg5daCv6boR5O2PlGlGb9xxNZSit7CmVjaTBqcLb3W8
jjdfr5vsS76aZtqQn/lTHWF4SDh+C/CqbcZiMwwYdsqq5h2+sW+4JRt0yIcULZOT
xmKWAC/l6u7wxfbZRZlzGchjVsRM931tnZEX5qi4i+P6JzvwhOAtYo4S/uZV6meu
+lqvdySbWPmYbJu/Ve1S9Lsqim9xygtQWW4iZ4H4bssQcEM7kOllsopZD16aCkGa
F0/FIHrhtwaOwJdrdthNF2NNuVNdN7BbXh7FZNfjiOwhezAjZvYICal1tdmNAoh5
62642JtdDNIDxmnsXy2yl+m+j/fIuLhNMe4e1xwBG5HXoqNskRdb3pBF6Eqmhhom
ke9XK3oizb8SdHsEp+Qiev4umZfkydDJgXIB8gCeaScuVi6r4jtkU5Qlo1LkDmFG
0gQwy7IyUH5Giznqn3q3iJ527Yo+zFZ6vUGTzI5ACxfA7+paBYdq0YrR4M5p+8SC
aJv8hz7X/ZoU1RyOoQC/98ZtdTs6LfZ/tbDp85miFg3wGQoNCfgCPGmnRxaNuU36
c0zONgJKiwF1C77CBQWgqLP1KzZpr77neA/U+ne1o6G0KJMCobHMFFcHsGag2TNq
ITUz6UnxHVYYizMvHnj6Wv2JSDKnYbjc873mAYBVe0SBndNSzjzikuevm98qjD8T
mGvBqbuPNaNfWkgqlrDz3X7iSgLRq/dAcavRHvFPL1vVgOl2hzOA5rohUUKEF9uT
Db0o5WH1IwH3FK6SmXHuPhgBt+AqhOfry+nBeLOCON9Gz+kJqZH9xDLunsEVH+c0
wFtxFMijUv/tyWoTUpZsq+iCFxaLB32/WBQZXuo+lvnL62WgI0vmXCWmL3A6C/Tx
fnOvJrTC0l4IdPmC0wXuPsl6nomIRuBf7DFLI6ZIhzBXquS7ELfTcnEm6LYFZrPU
1zgk9NuTz5qXlE3mmWB5kAMReTympgXf1BnPLv73ZAbxWih+iv1xsGsYQdtnWF0C
frGaoymvtILQFS9IuL4LnVeawVSiS4zFgBqtyRLox8d5jvopONgI7L13Cx4IfX5O
QeLXixA6+qxW9crSQMtF6ejXY1ocgKnEYH477GeJg9wUsWY86Qd1k3LAjesKnTYr
2VJ4MAQwE1hok9BvwhQ3MJd7ufGywr4lxhOLCY74S3wm/vW9+hmlVNSjGzRi3db/
oJxfDMcAQTwdFE9W17WhZEzkfMxpwcacVbQqRuqHFESJpvs6fQuvdV9LPqOK7YLp
yD7XCiAwkd8CRpB8IRpMuVM/ulJtD43q4Vqi7r7/qxcN8OuyTpvpxEtJPULgONxN
ZOrYXb/Qz4Dds7wtJOauxW36Tg9KL9z1O1bYWl4SS3iH/88jNqbcRDhTMfRSUvI8
BBzjJl1Fo/UBvLcjIG78YXeIaoQ4fN+qIDrRyDGqRW5+vDqshVRNtQXD4lm0PLDy
iubH36MyCNY9hmcvTxnOIWuimc2bCR7Wqjd19meoDfa3+MCsTzrvuWwskZegEwX5
PiY11YIvlWVwfP7O3VUfAD7aUgumOyY78H1IT3g4/lyC7NROxWcHjm3oeuOErc30
ipzqsdzbUoaaE31yVIpyVYUpD5hYWS1otvDuhrJzewa8+Jj8gusXotB+L2fz84ED
U1yz9qQxrB2+JaFmekSdFMLt7ULZDMPmvXGzHI2kM+wk/2Ar/ud/zyRTib6fqTfi
Ee8cbjoxJwwCL549Do9BKvRkxAT1gAkRI/W5uBEusVvHDrUWdVe+PrTfDcLxrxV6
UcLFLkVqeJXKI+FBySAoJIe69/frUht57xaS1cnK+1H/ZY+55paEXOkutUJ670Vj
jW0HOcHNsTRZuZq2cYqrXvOePyN0AHH9qUVVB5eOCLo+MjOIEZhSpgrAKXL3IuWk
iwgWB+5OBvqWGUkR0CFEGa8/R3crxe3cIPnbagYA8eJGyd5RyMDUGisCgC3OnBNn
pRzpN0WQfQ6MD9vPnJG89CFCoMqOBhtBnUgiKKvDoCsqCjONZG5kvwfiHjZnXJUX
o3uiW6UycnqdfhYRYQNDd68FqUjfGY0TIfB1Ok0nN26YbUHYcVz3n3X+S5UWV5wi
UkUSCzqdD1zVZ1j9cMmO9rL0k69BhOfA2/iN2vCpAQGo1cbg7sAGSD0BaegIhXab
tuOF/r/5jMzYT+Tqx8NxdFbPN/BpXqVgcCmh3o5e86krinot6hBA/pOWPxCdNSH1
ItVmtWCx24vM5h3zSR1dCTtyHPHG/ja5wzWvv8zIpb61RmYE9hjsMX8XL5df6OZ5
IIoMAc7GzhzgYMhEsHs4SROnIhumGGYWuVOLBD2jZK2+KFwdA38qYA5+U4aKi9Nk
yu/h6AopWdVjOXCK+WNcE+0T9Im+thPBAtgtydKrK2leFRUEStXN2DGP+PP761fX
9J7qCROv3F7YvTbzqH7feR1nBWTPrOfwMeP4MwxZA8n1SGqZ77dUyrf27fke7RDP
ZfKsRpO8Z4liQc2A2dGR35AAZF/vOxSNXH4GwztcAATbn0JmiUDe26kMPQc/CbM+
kkJcC1tcH36Od830/zGPMEr6/nX/qOPQmQrbTGaITKRUQXIoqdbTuFlYPVIKlA4g
svxNUanrAHVnBTsqHFY5u3WJfhSMoO88KUhDZiFRTa4BmIsSeE1A3bHwnYIz5ZoL
9bAi+hqs60TrCnOPQnnzs/mW97cxNwRoC62Gi/b+iYCycf2E4iu4JkjuvvbS+wBt
C2KeEqR80xtOLBQeESZYTDsLeScHHKylIwcnnlHs34C/OQL36IIpcKpy0RmOiCU7
SCH3wm8YvOD2IX6yJsL/S36U56/dxn3LeiuFEGuImgUIL4QWdOUlyPaltFBxetbo
JfRFrJRrz2suPcFUlvIgc88tFF8ksmprdRY6bobtOX9VH3c2/heSpGYPzU0X72Qg
dNkfXwwDs4qMxxILjgGxRLJvjyNt7ZFTye8zNsBwHicfeDXBIDPKKxSsgpsWhFSC
XJfi/WbNIjLGqNu6D46FA/Xd0JmjcvcZpI0eKtQTfu2V02+LLcjQClz6quLSIkv/
l57on+mVduzyz86Eyzeqhftd5JelB0HyzbmehMLkXw3uaoV/uYOCOjHEIxrzScwX
emaJxon4+Jno5v3hYZg6MH/bYwqQw5lHIGmIrORlD/4ta5esbZHBoYlWw5Uks+L1
xq9agWcAkOZH0TKKHV7UXgk7fW5BZIsnJ+OinI53uMVwnCQNfzGHQrJN4YS7LhaD
q55pib+1aQudjO9//zo4z9BTf5VhDpoadN8lOHvSygijx1KyBwFm+ewN5HGVcp3r
DnXioYco71LX6ruXfU9ydBi4DVfD73T/u4QusYYJJtjrUexg2NF6s5Xv9WE1nEOZ
elnIF+drBNGkeqm+EOquIVHV1pwy5rzgvXP+g//95a2E81h52Uhwqll/zMwDCRF3
TBZ++toIDLtjXr9yFLXpXFvf8AcvzhoXUZBZtzf5EytguX1iIWsQscnfC8L308qE
n1vR+DT0oWh/03xtTcXTXlr1ERdscabK6w06c/8f1OlKxTQNi6NP5weLVUwZUtU5
8yUtWZ0IOHu60nJiVBTruWXnJI0D96pqpxauWL8r2tqSQ1XWZxGzS6hpXS+dNxVS
VMqeTNcL8qtmO780mL4TgfsK5H67GPMdzg0TDe+RcC07eX/x+kuGClSkSFUMOINJ
a2GujofDETqOJhvJmw4Lwycct1dMsOA0f2NPp5ntMKmNYBkei6rlrTmuUFgoP4y3
4Mir86iMlRYfTUROXfq5qFGIawQ6wnPgAzQbtKzt5J2/E4GlQOUBaS4tti64l8oa
6BaJtDMjJVy051AfAZQIiV4srAlf2IH4DkU9J9nnL037u4oleOiWJYxJ4WncHzyb
qfVrDzOqWSNe5x2mdspeDy/FZwRjQJl/k29uAmXMAqwEEQUN9ZOrw54Q4FE2G4ui
v00vZ/+92n67zQyD4H0eehZEZJeTdOr/5wAmZkdhHaArmSzZzv2bcdBGCgIUBwPW
KDRDfBI8S6QNMLK/jeffkrQ82rANh9ZcSHHQ4DOnCg2jWbh8m30WsN1vNi3cXLwa
ceRLe4aCTEqobQjLCn7eECuI0lbszPaalrw8zTMId6Ln5YOGU8DwMRun8VeHEvFm
F4SvLSDMj2D7qoOtRYhyOrCHNd3iRWmvBH+kGoauHZeJDxesLYTf3VVAjG+bZA1z
/8Bk3xM0REMf6HaL7fCfHWzZc97GCqvo0GA5Pv6ww6073/BCS6ergBLDr/A7HEBX
r+IvGljRKn2KqZp1gRqF11LfiVxxKgw6QAaiXldSkWs6izuz3T5IN/63AmAaMiwc
6VdSf7v3QDNqOFdDvIbnWCLHvelnI2ie91zV6vk6YF9WHmB1j8zABaT2c88A7U3r
tPUrnA+od+DgyMUFL2zeQUT9ZHZIodfL3eSWiKrNB70VX35Dt1VNG4ovbK144sEf
EYt9oZoKrGg+TataSw5Ps4AwpxE8pPdABrJD1H9PNIephMGrFHFaUVChGbizePmV
5w08x9pzds1zRBPJh1U5VmkNxzAkvWRfHZrVK3QFjHiwGXpmZO2pK+soBDAuW6AH
zuxhsgeaV+iKZqjYIWBRqGDo0dkJsmmpRDbgl2N9yxRgpV9/vox9NfaBxPuGme0F
UXfy1nGaT/RPaZH6VTlipKtACoySlpebv8MAYt/NKHF2BQstPkzv90CtOzk7EzD9
0iYfjaIs/5SNhCTL9xZaaON/98NQNQmTKgqKm391flYrWGFLoTOcfqWnIPj0w2V4
ltXvm2IXDlXcZ9MAsSjDGAGIisGZb7fYO733bs4Zfxu0dMWzOV37vO0BhIqcs219
VvCp14rg28LRE4qaQf7trGUTt6wDgWHO++2l6dfwpkt0e+5v5M/6meQeWiUH1Y1o
zAnDgDxoga6KYLfcqPkKqlObkILX4Q+nEec/fFUYRVdcR89bXn15a8wNB+LLT9Id
pSaMZixl+ffU582oUGD6LsA+UxlFiftqsKI5rFK0pcIhgLlk3zRQntRSErz+0xpT
c7HJBjeFDGFyRchS/+bpBXnzDrc4PIte3m2ibd4WL9wy95ownTO9/pdpKl5jo/c/
q1oSe/955pBxr3bsr1nSPMKwGNc6YqijC/u/OotT/v4iWZWsdbnLgWXo18WOPakz
JtEAuaa6FndYFEufPimlx+GuyEdOKlIgl0Q15aWIMQbfyWQxQDS6LCmHDC/DD19b
9Gku5i8Lq2tcREt+rXRdXGbfzrgoqNsWB4TGqYgNiiSrZynmmR4RhWcGYJn9oFfl
BGLbiZVzVyQIoXJ+5ei7ny00AAuW/5LNzgj4DP5LiN2aQgQwEEHjEk+2flWBxxFN
DSHFT/9dBtbEq2rEjGc52d2X+FPD2iyTa9uvrC5GNifZrZMEPJ1eCO+PZIFBvpd4
TjyKQ43qOlRDpowmhy0sP0FwL2N1b+4PtfXtuCpBpzjsERR6tG7wZO9/kgy5NeH8
by85RAk0jtjhdHnC6tMd2Fl0lTGHq3oJArIJnXp/JOLDZ/dGsW+11Xaw+ROD3/au
yQ3dsFUxtlhWyfiUUqINbFeK0hp7Sg1m/6kqYf4kosA0wYMFK45DJoz0AF29Dx4G
TRrRPCKn2/zruU8Hox8JOBvne9ldQoVXxnECtgz2/pupViTP3kRIUR4gm/nwR+1D
WTucb61HA1ITC3k41UKYYKN4OnOIempzdrWk4RBrkPJFh0XcUxmCLq0+TkNXVNex
FcJbTvd/O5CdoY6ewEF2GeVIfVoEkUcjlxlWCevX5PJYyzfXRd6vZLhhOBrHj0bH
ZIraY6EYBz06NkpS9KIhMEBtgi+Zsejm6B/cAwB032hg0yPOhONt96IlsaR6dTE1
pRzI3tDmr3xtqnIH4W1TmxdoluO4KpCFgutt2XCpMWrzlS/+50kXlbSCwZJut65S
Ro9vhaj5qDr2PRIt7LjtmlsFOwrUbrug0uwq1Ise+4m3XmWBbKLcSe2w/0VGajJk
A3cShcc2gkO8rKVgjSbycvNxUDKXRngYcnRh24jN+2XeM+JapO6xmsRBdZQGKrYK
0/XlI4243BiFG4mQAVvwcYCfgimvguAIHCmnJ6o71cx7CGJSRt/G0OniY2ehW7k1
hRWnevX8hq1H83t+c+atHbcBeyFTMY7MBx0YcRkYdaY3CsJnUW0KL3iiIkCv2Xy+
xmG0KArtfzVqezUUIqf3YUicxOhUvOi8uvwvXSeA1VKt10YtzKOU2tZFX52uxaTp
07wjBZh2+h0uH3TgO2Y5iWO5KAqXYScJWpHlmEPymIVbzVqO7X33z6Q2VFBS5J/J
S3lJT4vo3HdoG6xP6sLJ3QyDg2ijxwqpEJRJmaKbOUXoPKqUtyVAKydfniO9aJ1D
Ny4fUrpUg8xuSHmHEForNz/EpWCBoN8hNFvmzcGTEfspXsEqY1EIh9eKnjVmGac8
83G88MU8apdCI7cpKIyBpyayyOBVSMhZn5yZV6tPVuMebO3AJ4i7nYAmDAnM8WMs
rMqcD0MhD/de+Gd3zbRbIKtpv/Xr7RXWHm1qnkHXvqTeirImwaFs13kh9/G3wpi3
7IxRpBLObuKGIhZl/BPCvN3MYmfreTLSxCW4as80NTdEOfGUYOI9/Rd/yvobxakr
nvjSHINnesFfViOKIOit88blY056L6cCAS4f7hvXMUDudqZZJ1lvtm/h2zY2Sn1A
jca2ZRj5jDlh0OMRL/NYFiyfn57AG+ahAeGIdh5E6ozWE0Wpc+68g4Tujv+Ap7WL
Q/DPZpCYBPKtz/s9nOC6H7fQ28CKxVGUEj64lxo6uZLsLynO1cNZYqxxBFh6uejL
nJOt5B3YQIMKvzOqFaSRit8QMSVvRrsLCoLH214RJpYPCjZsrtxZuc6YlxB7UKpU
yK2SeXoWNi8/yPnTKGMa0+lgMnDdIE6yP+6sTlk91yfDwhJ5VBVqxYSpcDA2eeOD
jpyModq7gMPisAIPnaWZaf1r7D/fOabA+uAJG7McuGt0z8Qme1y7w10WYMdvNFjV
8JAjweFLWbn6F5iEdDZwEOGIgdzfW4Oc4G+eM3vPcqOlnqFwCJOA1dU4FbF8HQSI
bvErVRE1UT2rOwlm4tjVP0tN/uZ1tMlsc11VnoNxwJZ8/SqqIxrcU1ZIkWCJ/ScW
+gaTmnVe3ZdFLfeoUtmoJeYd1nQsRW/X6S52+LeIHDMnIIXQy6zrb4Olb3jnU+P8
6/eZNFH6hTtpLhBi67Cn6eFZ0VpWtOxavkP/Dkk/RRVB+Nwvd9o/WOHhzjKfDhu2
cARN+ZKpW1aYcfjJ4KSejSwtYIE9qSx4OalH8otTRwMUpzsewwXXgsww1y7rQF8j
4swGz3ttz/ldfRODGh6KEnHH+KEnvfBUX+etG9npPC+8n4beuwyHOORQRkkTO/c8
ru8IutVNh5Iw3TN/G/R+lwZwM6ScALQpK5Kgryc3gWrh1JlZ8MrO4cftGzhbIh/f
vVwJ7In1n9LJDwjSvKCyBk9TZbFEINSbvQVwHAnvX1WUK3lF/VeMxjh6crNZwWrE
5s7AHhNhgq7dSiHM72bbF+YN4kdi64GyOp/c+1xPuSvhjc0iJZvebOqfEbTjBPSU
TRc5p67xrrM6bgd6e2ccQB7R/D95GjaodIJxvz5XjkHEsrLtAw6vHLyy63bJHman
bb5CZHHsRXzhd9FlZjN1ny0HzBH1N07ruul7grCsTYUg7H8phVazNIeqhppZfYSR
WunZqrnvVIS9iMa+k/Zo5reZXzMV7S33khKDILoExgqwmo5kzvXy/0fCj/8YFzyx
weAFP6HhOAVvBrYyZei0TCfghZM4gdzza1YVF77JEiak6x/j+rWXKCTH+6bscYfM
4SkgZVOoTgaYGVHqPC1PMP/pcX+tcwP8K5BUPT1r/VRf6LDc4cZhrQhiBYkG5TPz
RniZ4fsVi8wBElM82PXllF8v1bJcmJS0Gkqwti5l4IxubyMHNwtcl3ubZC+d65Zl
w9l3V1pVwMqauAlcNi1oREj0M7pY4Q9X7uSvy5CChZhkGpPz/lC53HjOT0vfvrXu
xXdjnFJtzXoErM/f7D0iAFB/ZhSCt14+fjlJE5gVDrP0ztTYUNGTWa97XQS5u3Wo
vVUx/Gty++MH2EPxfAjzBNnbZZ2fFDbeoZDMmAalkIvHuq03Tt9jJDFvcb0w9c8D
REtkQ7+cIkHxDbw9EHmIe14zKDNXuZ4JWTeY8QlfXF78aeQV47Uj8h4KwTptttV8
L/gEl2IFmNtb32idx/6QLK0aPHdh8pyj5SWXWcRRcGTzM+g8UdwM55HnESwsr9yF
eA8grgwa3GZZYJYtchOYdHVxOTt+vK/x3K2UQG3GbBSZ5EHX1o7eflh0ftm/SzCf
FS3XDTkOOJtmhBhQAx6CfgSd3huGxA2buwk02fJCFDE1bx4+qqNz4OS5idG5niEy
t2H9avhp8hv77/Yrw0IchfOYySxoEfG5pdw7Nc7ETdveFjkIonrrMwvx4TuURQIn
yf5ywhRtY2u8kqiwftSrQaDv2Qomx5HSjror8r9tabIyg+4bip9C9I1/L0YHaAoF
RPJqsn95/PvPzw2E71xe70Typ2Dmn3vq5n0NKCoTVE3Tkhdw4DHCmsXS7sKAyckN
szgnlzBCWMyX1mSzMFXqcHBbhSZ2/SWzsNdHnqYhkVPNRIWytTuEWI2t28XbwlYM
QO3HmPuVGK5eRzSQpbb1DtP/wLoKZuIBNg+QUzlf6XxPoIu6Wt+BaKV9W0JfG8il
IO1ksM1N3J6vGONuP7wN+aWLDYxYqnQWHdANrswWeKP1i1IeGz5HmIj3paCySfSI
4JZ43AEm+VdjPacfrWSULEDIwS9kMTNE4ro37VGDiku9R/YJBoqQcmp7MIwnCxgB
csJwMqaVwPPNhgwXLuZe3BMk6568Ww5L8rVS7rrZ2gBN5MSgAWWuANYIjLUqVs3k
p9XbZ0fjWboBooudK6lEnE9Ay8SSH8YFxspUxOjYzWFs3rRejY+FHi76hAfN1Wtj
fqlVhCIETq/X4lIovHFSeuJDF/VAqOJMo4JaOR1dHlaqGfk9M24286QKOX3bs3D6
QMTzynkR1FDJWL0dDStAI5ICmOyRxRyZ04qRTYW/HE55yk+sOI9GXC3bbtObSlXB
ruajMnWelrLf+JWtfJB1StyWWfEwfqVL+Xi+KKo9QemJp3IvQlvHaHPXcotNHP1B
wWH5m5xOPrp9rsrfaoVdRk9ONp/Q1CjIfPQUVmX6kOV5R5T9vDPdID2nvCwDij9x
tIarfojbT6WlNy5r+9xNv26alRqPPaqm+PxF8PbdN9/3VJZhyKKGHYVQIT0l72a3
MjiReqiQPMWB3EKLjAO3rQxXjoCvIOVmaiNOojFQSxoHFK7CIjO4RBrPTLmZcaxu
kIOGGYt4fjZwH/i5S+KUV+62XMZQVSnEYcKJypUx4KH8sVo/SS7RpjOeIruQlHrr
zNutJEsSgEhptd92Vwj2fSuHkZgZcVJqFtm6rcTicLPfH7Urr3XOg38aIOBaulJL
IdgM63Gba9PsR4Kohvgktkj3Ri0fKq98eRMWwFV7wtk0WKdnCwOeKbs7jzPM/eIz
sPMrdgoNeMV7VYYYnqR4D6XXqFKF3iPGeG9ZC4n9/OpzGIFaBOLpZdXrkyQvjDfu
5MpBKFtcdhehMf0+NPjI0kWOkqBvGhOsJsOlPoyK0/stYLnQfpfRH7Xb6wo4VtTV
HIVjAYIe1A1Ka4wcE4MbY7qEX7XXPxYg+YIqRI+wb4aKq7yjxuqRqEL2jCU0zcOY
k11Z5VB1l8Uq9uxUohPxSSKNm0hZ94bJPggUHSwiHbX95bFInN41nfsellq9Xmwj
6y+TJPeT9bVn8Jlj1WueKyHC3qx0ddI8/9sZwILtR5f7iCx3l+Iw+k4unRtwVj/b
MLfbHtbt+65IU97cZqnG+lMo6DVZtsxXJW0oD/FrA0lGINROkvZDXwQg8Ig/9v8B
CRJwRDh66oCzKgk//qJngjGw4aBoB56a4sZetTKm2F8nvUhS+muvDi6iC4d7ec1I
kMW3vMJjzc/cwA5ndIgKZ2Wkg+MryCIme3fey42xbizx14sfH2IYYW6JC96CZbs8
NXo6v+vDJwfHj1q/Tpy3NQrBtAC7P/m3eSfrFfU9ibDy/8aG0eMIJ3thRqN4Lzg7
TwwgE2Wqxab0WaKkf8Rz3JqSaCEOqYqdtHpisOsnjscL8U10kksQIYsoyv97mFne
8ZzSKDzzc3poC/xcVszaytxKmHe6Cw6x96TOmlI1T9SXw9M6ejA8xjYhVpWztnDI
Y9ZKQ7G5AHMYV0ft3/YkrLEHQyIH1tD9mvzl2ZIJY7WL2TRJ5/MLZZZaItqc5BUx
m8faxzehdjP9TzwHgF/3FwAYSVZ4YKTiCvJ6gX5yUIJTI1IZRbEI4fiiu3FP+H+i
K4lvUR1awN1fBqT2V0D61uCbfyA1JXY3zAH/uvDA3Xis9e8Z2Mo/tGFXwXyHy/be
ueVZ5wDELFXTJKEKCGqWVptbO5ECjHrPDVKi3QWJTozNp9mGcAKlMRpWzekE6Z+d
iPBgRr9hu8fu9GTTgVGsgXTFYPnLAgi3jjPaxL5WHVZyxHVvi2tdB0LRJemJ31w0
Lt+qkU95Fk94IRfG8qmjSuISom/4/CI8+w74a28sQDPchsY1FPBEx9kw22Jf+qUm
v17weQwxeh3n++JVO3bvwtP91ZxoRaTsU+egaSYxcedf9qCUUVEgz4nEK0DPsSKf
5EuGIym+63byGF260zn33DxvUxFGS/tLbH+XDaU5sfB9gzex1BRCaNiyvg4xvDmX
cOvBYXGgwN/FrBVMrxYQWcGE/b166YTADDJV5K8z+AJofbiew/ev73frXH46wqJr
YvJSCjLuNu1CJG0Ij5Mvb+iFCMYJIJRup1yecDbagGwTkypPeQdPvMKvppeiX5Av
wDKhc1s913Bd1I+St4tidwWa3sZYgITERSzgvAb6rnzefnAEzqDJ7ObWPdaUal8a
51SN+livemN5WFwTJc7d86tHHakpqPPk1f0t2LB5/pzsmTH1wnmpgV5JSsQPRqMJ
y6No1Iff/f3ygj1/3PCV5OEKm3l7g3swGNDFsa/Sdi5TxLdi6DdYP6RIaV8ypxj8
WwNw9Qh46YXuEZrqIo6Qn8n1hSRzWszQw5x3MUTsxbQnIGM6wI1rpd3VFdugXEIx
1F6YSibd3diXqpXI7816HEdyGZdFg+HI0VQXpICA+52oX0e7O78oQbl44z231b01
UYZ2V07Gv1brQWu2Y5gAv5/yVXIjHXqcWaVaQ+PGBnXR+uY0X8svUSI67uHpkb0i
19wZRCPuJAlrv5AHwMEKbkDjMhc30C2iRHC8+DioA0I6PCbpidO3FBr3P6h+fFMr
CQI8NetGHK41ZPGV3CkHLlkuOBZgo37FbKL8y7BoP5Ox23IvekSuYsHxvU84V21t
o7b0HroaTvyipTf3he6X/NCbFQu3uWMMQTG4Mo1rzK8u7tYNAkP/ACpBNw0himjV
YnewDqGbf5BHcWT+m0bpPDO6koOUrgqid+lPxMIajZFkYZxgFNwsc/kSjpw8sVQa
jHcJYomloTjfd8rplKp7cADx8WpOJ+V6gkklalfo7v68HsVCYl3gVJzw+UHiYG0e
+IyLusPIBLppfSTzG9VEoqltYHz1/4YY4m/c2mN7cD1NvzXN58DOhnCXlkMPEW9P
Zajs0wzINBk9M4IjORDgqUknzEgHMbBZLkDoBMBEojCbhV6T70EB0pBPp9/2kmHE
ybRnN0eDjdXNLuo9L+m/ZBHUv2iwUCLjmT0XhimpvziDrKGGBxTxqCpDqlYa+FDH
Tu14bDnYGNMQSCgdG7XDm2ahkQRLwTbTsYpNaEuQj9s4n/L/mLs8/mC+6RtOijBd
+DhHjAbjGV4f5Dh2w8xLnBeCZ4mw1WFuvhh3rOtUHcLYiF33sIVJM17q+IneF5k2
88Fh7W6Qg89j8y81e29hLMfs+yBIiHYchSeXDS6sdko0HTlEZCWN1BWt4S59Q6Ae
693eu+Lxguf7/Oc0XHKxWN/CHgeUYdlpFrgXeoCkCkmF9KBjtlkGNZOjhPgrgZhK
f0zizTxn+4YypWDImhO3TohK4JyIt0q1MaNKd6Rgc3xW6FnwX7YCvcCMAtdNRgmS
KzMyOZF8wEYXN84f4ego6hWmAptkRxlR9vrXNYYfWiaSwpdL/7R2TbqWKygh4/Zr
fGNSE68UA2hTYdRjzn9cCNxHUMCEo+OuDfXKRqx9uXnQxGAUr3TT1P7QgFLv4MiG
m/b1jC9cEAarGTsewHu1iM5atd71SCrY4Ogr2YlS+gRDBXpTcN1p+QrVnum9z7qo
OQkoWAlSsCS5xSMQIZVm9PyPsts9qszTmh7m474I0urjpcjPd1kGM7/nMtLRm8oM
AK7MuobULw4+469JsDSBu2/6mBhdJiyvcpJooT1rcAHMcrAt4F+6EYtOfy6sMakn
HBexEis7gY1YkjmgsUyqPayoqtxavwztZOtVIfeobKrlCMJr6Nyu9J8wuyt3ee0x
OtZ6cki2UxjllgOg7alJZOlXLQ/k6JMLpdMFIxfzjWffdc08Te4S3UFp9NNJ91P/
dBjkKnGGLfWn8pE3/tg32jRFu3zC/mMMJvfXE/F1CLy+x9ejQakYXDa8iMUO098x
5sF3md151AMqfZVyPaSBurrPKeeIG5n38k+8lp5FsJ7R8L6bUmYnPXnpH9qt89Bi
yVe6h2jPTD1mk4I5cNRH3HLYxdpmyEcbGnUNtTnXf/UbuIns6ceZY8dllF5IA7sg
PBGQGHvrlO8HGLp1Wj2pErUfh7KBrV+gHM306E+YKo6pLDGtzi+iyntb+wWomZWw
ZmTDt0VdLJ/siGBoX3K2UuwwxNGQYeChwRANcP9CVRXx4zGhT7tNC7+EIcxA/bEO
ix52lZ+p5LXaHa5xgVZnO6CDM1wRbJWPeOjf5CFPBhY/AR5q3dfkm4Nl0BRY91lr
HJlVW8Sy/KQ/nC2HEPaWbQn0EvIyExG3Ii2DVb+K2oQ4AsO1H12fRiLIqojDgKEa
On3I7Ghb2SO5cNrdO33uxgc7o6lQjVOhe26soEnf0KYEvnpNwYgk2z6Ci9IUuDxG
EJTxrr3dQj6FbmQpSm0LrMpmHFx0bdoa4QrGAfPQpNInoE+E6IdrivFYmLyDxsZ8
4EqIV0xNaNz45McD+GUxN1ivMDAJpesGpa0gk3qwcIpl7GVlvX5H1UBkNMyxGRry
DIuyrlxXVpcRoeEduLS/A2oFA09mljFDI3V7eFPgRlXUv+A4dSKXrg2kO14g2VEe
ON5F9nOsH2ZEES9srqqa6wpuqVI9NsZEnrIwJLW71Zinha/GUeyybDoeNeoA2q7T
TTXiVIp6ez57HrMtFEe13EFMcZoE3qZ9nIHjn6kEmyyDUxiIuL0/0wwef7GurSQk
mF0UyNm2vmF7IXApd2PNMrdQ1ofivZldbq2oz5PTCBZIgaVRyOoNopz4nIcEJvQl
F9NuXR8eupa5ACKBIysXezcS6y8qSOAaaMBQ7KesjhI4tr7RmyxPXkxTA7BJv5Np
nNAALI002xxyAEnMUEZd4XIi9kAX51YVPeBtQdhskJ1ZDZIp+f6jKbLx/KCAvtD/
S/3XkrBzLbu8MocBNqgONjjo2Z07g83mm4SKMP3sgv9PQ+pJfV3dGwEVNrS5CvE4
wnAYIHP4XdIi+sztDdojrjAp+uoLey5Id+lOIVG5bjRC0c206yfIsD5F+MEtsVH1
NSS3I+9Hh0kwxXCZ7XWxBywj5GZ/rJLbqpM2TsobAaQE8L8YmNzAziaoFQ7zbj1k
xcF5vWigTlc7wrLx/M0Cc/LfvsV8TPGqlh7MCWX5kRPM4anoZUBdjr44qtVVxWvA
RoOdBbUoamG4EGtHKjoW24BCmrZ39Ytd2tk5pM44kAU8DzQcIeV6YA40y9adcafY
WanI5yek2snoOu+t7pTmcdr+x7RNJFXQ4lpZMq0IUsNyeQ0S8D0KEw6G9l76MPZD
9K0V4VGZitN/anCaL+fwxBX7rzPFgqP+9rrh7uMm3S5XQX6b/arQ0uh7rwz2juxU
sAE4IF5VqY6ue5eB0orw4AD1Ld8rGXGZ32KeW3vV8Bzhgf7037laV99WfbqrTyuO
1VaPUW34elIzmnpjO36aLPGHc9ntOAGbIjxwydoxTQWPp9Tu0AXx0oBBl/BlJg4O
BzQgEzvxPvWdUmYz0Rsd/Hw2J5OJ94yn4ZNnXSDLQyw7dQ60rmMxsHphiYNlMc8N
J8RB+92+epOVXYpBkGPQaOgEAv3T049n9z81+COWISurlpLNQsuBM+VydIGRflGy
Ihxq2tXoH+E88FZo0gal7juyJfdPXA/os2eJpMDzXYLrv3Bet913IK209jZyg7+8
hyd1WJOS8mr2B3YFcwDpgJ+7DiDjNhMEb7weaRjM1aNb7VMQwuf9x67Al21E2Frq
nrqDtVsPy04A6PXL7+gXbDOgcaShVUCInh4cEF1AH8XFBB8y2zSqq84cYKPHYTyt
K09JgYLyA0zyK4wXI3uR1lYpofClpz2eqf4iyDoRTX6bhkcz/twHdBqzAf3nNLNZ
2qIhW85yIykm026WaNs/0knD7iRSLg8Z7At7rvrVmxE3+PQTYBA0s2QrpWjinOT4
VCsJ9rf+uW6/8HVFetRQBqm70Y1exDhEbA76DTdXMSyyIjwnyoarq3B1VuRSEWNz
wjctzNzG2f+Z82KaxZ1Zq44S5DMib/rv4Fmx/gdTmje/xU1N6kKhbPV/vr01Ri7h
FYk9cuYsV20g2XJNfAB5ktfGjIODA76UvCd9L1uED4zki+4aCPtUFU5TyCJbRayQ
3xUv0yZJ0FV+zTcguZi2WOFlQxo21ipi/H5gSk0BNaAlnZJIo/UaQ99rdyd/fj7M
jQJcL0sCp742qj3Cxnl9FCgU0Z2tLHuIvbjdElrJazoxCEUN1GThjOFRsIcwtVqZ
kslKbLWALL1/UAHrVJlRRz+RVD09/mbhmPFGa+J1bdeTWuQ6wozcBZsEHCEcCs2H
zq/ee5056seAjorn6h8fv/HPr0tMVnKfqjYJAg7zMwyiX3S2n6jSLf6NvslOjBMR
+ixHmybiirF/X2Om82k7zVymW2o23z5KmMdXcUj5xgWqx7rfgLtuImdeiT3NDcbp
xC6xbjgA1aT8gxAEoDT7WkWAVWCJUygprVtbRm93WKM6FonkR7l/8SklWAsmTFxn
lU4iFTVczd7XMyqziwsAkVNJnt8oF4QzGLRLhAuJH6klwfuT0ew2G0f3hEa6zhHr
Pgl+FMPjaPtLMGn/xrTpOMkpQhCVneSUfb/w9clLeo5tz4OVx3EjxBYYj84F/EOx
rfZvef3maLADjOR37UZnOggt/S6rjoYMQuM8HGW+YLqSwKXpjOkswzBry2JyLudC
NR3Rs9IgdtSPvdknhh1QqXME3O6k3fVL7xq4V0FwfZlxENXsn8gBPlpqL6hxQt3Q
TOIJyM0/oj2k7JBcSDRAerDa0a5n6hasNLaFamY4eRqdf/zRpu3MfHnnoVV+hsli
FUrv+Gq13I37OGKIbLyHj2U7OkNCWoKD0PnptkLPW1cCHKdXUIu+C2/1sAYFWKbs
2Rrr5gCFxcqV4Yk9XzchaYIEQ9Vew4922SaJ2iWhp3pti4akq3dPZXdQBClc1T7z
fxFatEN8A0l/L8ipVrQM1dvWR//Sawiy+zTM8XIhZEeW7J/abFy44Gn06K5+WI6L
CuvtzIjMcTnVpKsUXNviypwyvnrASp+ZdCoLoW9DfKnP6D/VUvmz+11dojqNjdGW
Rdi8oo1hmtuNWDzE5MUpPLltjx62hyKUMjlGdlyRmD45dIAlGynluVaVJ7SCaq31
i40jDGdLvp4eXCaW5QnixjgkKO1UPosoKOOtbMKrqYISYzdSykc5b+gELO1CgrKp
719OH0wIOJ/6Oqeb+AjB6clSc81hMpxtDt4IBTqDt5tKhFEPL6o4eZoFrtHkX5q1
eGm7KxN4SVFZr3YkWUgxumf2gALtLUku37cFZn8XxUeRAu9GHw5CjuZqLPb3+T1h
5fbWctkrxgg94+c4AVZHn1U4hYv/RDmHrPRFR04sy05FR9s9OXYmzO0Xp0wD9QTZ
n9avP34T3JrJoEVqu8x6wwrxaOot6QVQLrpvi6OdlK1rLv/1DWKj8loR2DRpp5Kl
XDFPP7FSexIIzn6KCavu+e8M134C+pgZftbloyzxbtIQlsl7prpKbA1NjQkrhyMv
zpQVi57E6ZLH+cuZZQpKm78Z/Z7A0DwdWVCLnvktJGso70udDkYsZXrSlMnPB/aN
BYW0ylDE10IF+UASLW7LtAjO1+9cOm1C8tOXLM4yybAoZ0t6USQxnohzYWYIzxXf
usanl+8IQKfH0vUuQTc5fly6LPzc2wgHXZUJfVKm+bhDvPNkenERmI+bQ9rraR/G
sVUo0/CBWVZNgg4FbL+vEwpntkR71fEAR194qt2DIz9pxSs3Cjaj7ZiM7UBXzwBF
Ybu2CQr4WegW+p2k0H02lDV1/dfMpqAl8S5Scpd8VwHFC/ivxyQlhIHrdVqEDHCs
oaJ4ZQ/hCMK+xTLY+fTBSS6ndErlHoG+hBDMr9rPkbr7Y7vEu2ViFKs2CwY1sq6A
qIN8j3k3U3xgeDiYza7W6csiKYjH1I3D9+Me+Wq5LACQNnwM4C5nI94LqFmBqLmg
RunKaDE9fkT7/z9RpBF9XaR3/cpC55hcLalw0Fa+8cZIYnmF7M0X8ootddSNW99c
XI+Tuqeq1AqeCJQRtpIFkHSabRJ9xFVRLRCAVfbbpCZ2ETXPjdPOsYv7L8+AfXv8
Lox+LhISx/+ve26F0mJC+9GCayt2cxECQqTTvsUkcIxXKxH4V39G4gJR8hz2or5L
tGi5XtGQkOTEv6+wQN10pL+yVNOXkO718XDwTKWR4hKIPMNuhUNuH/qHWXOt3WxM
ex52BhKOyMdejQeZZSWhHyZySK1F06HcdF02ZU6RX09lISuxChEmzyZhh458h2gv
VZiVex0b6RjBo4Tw6pQsAyLPkhF2iOWPVbQJNCnorEhfGuMCyCdFtiEjPojqNSiZ
wIbVyivEmCMt1lmwa9NUVycYTLWbZFIWbuQSBR41Gysy79itHDCo0lH8KY/omL5f
ynpm4Cd1LDpUL97U9Gv3QdCIYwkaNDcUaTVceC/9Y/xnTozK9DGZpBH3CuWUZjKn
/Ctikyhdr97dw2+W/DTWLDG/vjRIKYuxP/1rtdTR344Dv9p/QNpwgz5I/4oRPI98
6uEEYfrEYcMe7M197nPIKtepHJNkF/v6OiwE7KeyCE3PcpQsGMhAne+2rHm6UheD
7OI25wuBifsVFTs2YSzb7c354g4aANmVv8cFneeFlB5Z/BbVEc9aVR7eKOv9oy0Z
X0sxw5VvdilAIpzXfd51potlWcr3T7aeyFkYv5xntEav0OgOf37y1qorracpdreO
ZZQXhIBmNs1LzmDIpekjNZ9QoRJ2I4yULQh10/FuZOB5q96DmdZcLpyPj07GjzTJ
tWubgHVVllPFvnM3eCmCBn9DCp1Yj5r5EWaSM9JtrLTXKl4sPFU5EFRq8XObNeL3
GbHgJVKEyIpL/R9A+kjbEJ1ooQ8qVMiqETOBY8v74L8VKbsaQCe4spAmPJDPfFN4
Y0RuYRpc0ZoaOGTapuWJlMo4Q6Z9j87DXoeR7aSGlYcVYGuN6Cr50OWiHa7lWI/I
iKwMCEtyl4iqE3DdHpwPMZZ4ZRKf6wy+kGw4XWTQ4LoParW00+CX5UIQkDyc9mKQ
JS9VD37gVkM/EE/4X4gQw1PnEoqtx6sZcFyxV6w887TFqgRBVv4m0mP9tkfGQNNZ
FN7RBh7PbnU1OggeMJaq5TBRrHLMjO8mpueFe0cT0yLZx2OwdPwhFZoi+c7V9myN
uG/MY3c5Rer1otp0/Or5B7UPwq10PEO9dsx4d5PIqUIS0ispdT8oe68b2SGKTsOv
BCumfzrepiEwJGv/ZiRT7kSIaS3bKMJ/riKauF5axgBbssEf2mvd93LOtQ1ELGkW
ZrC00G/nAVosSpnsyXk5tcjGIbgPvQOKp/Xv6Wh3VKzkoT5g/1rJFNMqlIeHYHrn
F6PUOGeLIZrOAGscUarkRkGawU07pyBiUHk+IbyGj0ywF/ovA99q0u/3IMNyUmsb
0wC6LrxPBLse7garFTNHJFgxFP987VM/lp1bJKrRRFsZHnAzqA0GSdFvMLv9S1Qx
aokYdKuSHMDtFmUYq9jCX8uMOx2UHWClqNaUAKycmUD4yD4wE6J5ACQ30Gq5dGX0
It6v6f132km3tAb+FOEgDkpGlooNEiknsXOY7LWKC8lZouq6uDh8vY0HvRJ2xA5r
VBh7Ak4ZC7IDa04hZtAocHqLOaheUKYpp70jw5qJLoo7JWTpBbEEMzE5X6ED9TAZ
smT0VLeWAeifAE4/85pgDLEkZAkRxySNNsZUoB9KC3rVw2XGybmQr855s3JMzkAE
hQNu4oe1slaNHxLeK1+Na4OFJhcRFhL2TlXhn86M4iFGtkNTzyFpzH2S61ziT9Wg
kh+jTPAGkgsaPbG7lU8+k66VOfK2N+WpHt0jY3W63gSkf42Moix0gQ4ElUpF/Ws+
ALSHUCFG4obmK5pvMK1ggYbH491l0ZSdMWzGL4bOOWByzM4vDRmSxmHvnGEDcSXf
Xs4XqfFUTfx1tyzCiXokd+VCg9ckacCBvh5Ojm4kJF9fmhnMgph0Eo9zOZ6MO0nf
Y2hL4Eo+jNyHe5mEY2UkD1Z1sbtBvSXgvozw/SldXLfVpls0hntF6L0RxzChcPrH
RjGxUTkrDSmaZEG1pTJl7FaBj8ZrtGhvflXji09+EV762SDO2SNGlT5BjwFed3V0
IjBE4nHut4aDwx0e+YiSd7tUGo5v1l8Z3yC7XGllucNpiPX2aD3eUi3pETRSze9d
N8wsMpeU/20j0E0QIyZ2DnNYXF+8AhU/uIISR6/zkIVxMbtcaeBU+TALl0UBdGG+
HSeB6TjhxtRehTwYNLxinECoV6pqI58U6lHKn2DHREA28cnBX1JlJlcZ4ZZA5spw
ShAY0o7jZsBG4e/e6Y/xzNmN28Eo0mGNlG68xCiBbXnc1XUD5tTrnakQmHCoFNjy
acayBSMoU51wpdVj0+s1u//rrsoo7UtdFghQJ79HnPZ6he+Rz9Ph9uNAR/IZaBXU
TylHCeaAG0/RVUxr0lDQhPY3t7DLsvx58qayYpT2+YgTY5JPK0hq7oX/JhGqaxe6
ApoWcgG1QjqRwqFpXaoCbYJ4KoR9vQOe07bYyDmBsMfDK+CtUct8SaZn1s8xqLat
LKfQ51AAqLDkOPPl/TBFqJQzunfZMixBW20n0aXr7zTiv4OVbwo92e08u4vqZWMH
2o/8kBHkFBQnFDlggjTTrYaoJ4iLerClwh9hrQrITG/q6quUyZfmSjmkzrOBROU+
aFct/0pV7e/BSwmIse3uFTxMXvkl3ogshLSlS5cV/4shfWZvSTCbnkUDQG2zD56u
rQhP8nPUGKSc+Gw91SjcrkGVzn9h64HmChIXnYI/OStZ6SEAN9O1WZQoZYN1UWw6
PUlFhyKmfYPR/K/P990Rnh+vonbfg73R6BQrXI8AeQtVWZ4Bd9vgp9njWCkv1r6Q
MdGY5YLnQCT03pEphHkRKUuhdCrX+TAztxgqU++QnhFQ1oecJjqqWfKfiYjCYkO2
05FM9+VNNnvZXjMfFjoAtev4DQIH8Kb1dSORNtbMypvirI/1NWOBXHDmhO5qdhUd
lHftUvZXUIQ96OgEPGZOdcuCEaFA+m9Av9gAYuBfmxRuqAQFC4tluKjy33CtXAxR
sUnvSdmnk4P8mzoOMqh2W+BxzmZQvWbxlmPlVBwBoiEpRCsbWYi9TXLlYObRdqMj
zgLrzH0Nlbjc2pqg2jG29wLeIonsbtp/vpxWR6WfcjViSJnlNdlwC/4r1Vp3jB4D
Wkfu8Ij3MEMo/54tF8YDHGRHYnmr6p7b703BeYw3ndAhMxrTdZbBmmBQyJSk248S
TzUvEcWkYSDGDa+McCF71RQfceReXdMEZc7+m6MiReLiU2+vdZRl0sWVP6vzCb7p
PlQwYSVS3cj3EGwK5BJr0HrD+Y7DUjH76kocv2s6M27CAXCnvHG+O/j5SWg063EK
oOZRixr99G5fvjElW4nZ0PdV6/A8mb8c2kZ9wdl3JjvQlTFrTLTqHtnYnppTmphf
xAR235iySVL3Gz+mwbfrPxpwU+CB5ivOcwvpif5u8HTuA675URHdtg4pMhQTVJoJ
ITXy17/EcjLWIZa+3lwvfAXRVmmf9PqAYEQSgC62m4/E130Mt4U3Vc1Gse2yajPg
y1o2ePUehJ/zLXsdzeln6OwAsMyFmIqqwoN14R8gGmyC26+vCbUOfhxuVdJYBu7D
CnSrswalL9cNU0vOMCAtT3Smv6NxfN1jwiUmEtud8X4wmMdacI/XxWAW3U7uh1yr
rXB2D5XZ/THx0SNys8CI8PsGbxMnIFAIYzqS2kicqg6ICRquJZX5KxONi8a+seU6
LQtuwNo0nAsFf4NDtLCfRcG/gYNnTwEnW/hEjdirBLrJmkEYiRYSK8G3j+Bm7L/q
HthXHa7VCx7w2x/6ZUdKoXCOZVUOiZDYlChUa6lObqYdLtTNZUmrglSN2gNvYt05
48evSCE7R8ZzuwAshu/mkewvsxbR9o0EsctVBIsUqtE4bogzq3IYeYU1zCcOZQwG
I/BiVmiZCKMbz75dSWi3aussIbRO4e68qvTIjSWsNPpZcoJwkAtJemxr9oqaS65z
S7k2GfBExp/dZEcOFlawMvs2WcS6GbkgHZp4+wrhjDgcbNCz6747gcDJ0pfXEs+0
dL1aKL5aTSgGx1RCuK2ohTmdjUOhAW01aKW3VT3sv3BSYdQoi7ihEpk6bYGDkiFp
Qf8Lbr/rmChYEI1KhWnx9QbuRYIZAWJ3hG5uBv9sjlnfN/j5fDg4D8ooEfxz69lh
Y+KZuEeIFPcV2eohEufreXwwbVlhdUVtGJ18bgUDNr5X49N251Ok63tvOQXarI8T
I5q7S++Myhv+1edDUkVpTGaaBli7ti9W6CX6HHDwmMkpDD1h9VnfNU8Za043IOGi
3Ls45MYmcJa6QkOYSsbVHiUEfi1ppSx4gDqN1cfLJcf4+7znlNGOc23hb5CkhZdh
EFtJ8dYxDDjR3Nx9DdIGQifqcXbnGcg183dNP2N9qTXHZBj9iV2lzA5NVAeJ+kpx
8SQ4iSu3jayztYa3r3KCliqxO2VWG1DDlR/WQh0XEFuj51QOSNXiBoQn5CxMxSXV
jxtuP3IKkuDeZgVeII8Wt9KLfuDcWNGyyV1ju9c6xO9+LRU9tkXtoTylhooUFbWW
Ij1fPvkkhNKtlUFMkC7p+B/e65wfIEbvcS1We8Gqwy+2nqoNQM9THa5Hqnd1m2pB
7ZdNBP/56/FI7Xbflqa1NOg+EDrRvgJ3ej7ZW7xQkbjnGDWnUlBx1VkzeQb2H2eZ
+FyFkGMQPFHuGF4rf1SKdhufeQLpUYt6HTPjd8A6KoEGQQCeYWxULA0/shny2g75
jii9DSCYHtXrI63t4MrjMhoknawHR9Cuwi7vfI6K57JUyaIQzioXScvOut5JGz12
Rk44wAGoyTyMfyhweaYj7NOpFvTCa0w6S/wmPnFWbTI44pUNrC+IHgXibqm133TC
fV7Hhir8TojwgiSf6f3bg/2lo+gq7KOofmqABOUzaAbxWiNHXrlu0JnJscCy7O1c
TLyzcJ0n8T904t9nsRDZMeqSaMI+IvukhX8OEeb9ZfypS6c1mKFbgHF375WYAgD9
+2cAopg5AWMu87J/r+/uyGbFpDDq2RTuNMrBGW+51agUxki46KtGbrH28cehXkIo
gwM6KQJqsPzTfwQ+lGzqsaiQBWqG90nepXNXqnOP+7QjZds8/HaieYMVby0dck0S
b1Q+td0YxhBGc28VzwWOQuHGwIk8aZR0i/ygtvQtH8wC51LmWqNfOp10+uY8Ss9U
3PVWDTkixLkfHp3LBfctaP1Lf7dc9iH2VFWZt39x2PV3tGI5+MLAycFkky4BWWwO
k8apoucLg34SM+Zr45f6ghLPP99LmokUXo1c+KiY/SkqdYN73IDdgPpkKdC5x6ZR
PCGpKARIpRXLVyFrwA7yyRvD2JRC9Hfz886uAMSM9bmZYbQQJb7f+QH7NdkH5NXa
T1fbzJceWcwkcWh8tVeHQAZHaPAiAL0+F4KI39kfXjmy9DLBcLkXKC7F/hMHNY7k
EOm86vWCULHfkkeQjJ8+XTQ95uCKF78G/5XtEHLEliKlY1dezZ331zgOEFqb++K3
urFyxL7ti3JPCq+e57e+kzaPJeyTY7GeJY0fSTRfnGcyAVmqYcarThGjUDR/xfQ1
AmNcKFiGVQWZmkF43h96nnf0t18im7B7OTAgE1Xudsi0iIPdvoyBcGiUYOw5hbws
1mSIhDEln693DMENk32Vp5Nrmu/rIteDDrZ8bwE7Q+2zpYDmWvdFbAHeVFpXEzcA
81XOIEYEeeRltJqI1rvP2pi8DJEP0eGgbWrtafIdAa86neel/baMOkCo0C5qlgx2
jnojcIIubLbRwak/tH7VdDxx+MLf6fdCei8qGwkHTYq36aY7ZZ6qdQBeCmty0G8x
h2Lq7eEmdgnC7Tg3rvZrH7HmmgqLTQxghtwzZk28JiRuRgBJb72gxC8xOAB/xt7k
dk6/mBzLBTXeLdV1WF6AmmfoKT0kMo2f5pvv0bauVPrx9VokWlgKjYTmphIJfgwk
iv8pdfaCPl/JuSgDJ+n1Gc2+aDJ0vuY7VGbOfofQUTXSfsMWM7hnVHs2ru1nello
XoE7Z87wsMX16ElT5j+zoh82wVQmDTHtgcHMkp6wh0x2YHXC6qPM/0Ql7wIuD3u4
Ij5ioRvw2PU521UO070vQQ6gCwvD7/kqN2UXbeomEPLQoWwQSTkQSEtXr+RutosA
g2OHVs960cqTJ5ENTZeE9VEbMDLEhBn6k+eZW1hBv9pqUi7d88jH/2g/iB+sKs11
So+ZbWZHX35Req6WK3Wd1u571iCXPJocMJV/qhYzl/ZIe/nqwqMNkyGu3eBbWKNN
uhq1jE5Zg5SV7ndISYhv/aH1DTkF4NWFr+FarBnkYjXyM2Kd2d2RjQZUXj+NrKKT
7BMy/5ubiNPQVN4/ZzFGLW9yjEX5LsSFcILvqAPTIUTUknpuw3oKk1N/DH9CH2e3
PnktORrLQD70LhBz5G2FX4ZrwqUxPCi08aSG+4tq0OqwDz6nTJ4QMvUsSPEMpoBx
eBITQTad2Nb/fCGza0dks86p5jp/g3LK8BY4gEG6AIC+QU7arPBQ48MyDnXFPoJE
ZNInSaauaEDrhzmvfK0ny6zHKP7bDm6CdhW/oX1pTUYBcQhfA95zlG62x69jOirH
6qzQdWV+uVke0kdvLO3vDRS1yHGjFpM0YDsRiZRB30kejleB2VeKWhEFGWIm31i1
Sie3y6RTvx8o4z4JRQ1tjk0wA2tXpMZUJloXcUTokmYK50PSBBGbspyYnGaFiiWK
nTauxCuHO/E/sKGJDKiKMf7cRd/yCLajj3LerkpN3HH02UxerHC/y4MXU2foDkzi
1GMid33jfm9oRHPdNOAISIL3VY+1HdxeZCXseTWAJfJueOmW+QgMMSvBkjepuKUL
rsMzDYaAwrJBYWQLL2n7d2O5KGa4QioACATW4fkS2lf3IGPSHtEfr0brjnk2eYCL
L9dHELG+MTyiTCTRo4YW3wMzBaia2zia+AKrH2lRcgRjbyyazBEV1VK9jFeTO7g5
2Mh1YuwADfJK2znlmBGnKV3a071Q5IoqDya8C94QOmJdA7kR0sSW51tB6/VPgyrl
342L1GZWlVl+qUpEplmp4sAVKqlMmuCfzsw8rLcJ3mGAZxN/r2YdByrPhQaj/HxR
qB+GFvb6c6wF8ADetGkI3l8zCXF+5ouVZc8goV2sehDklRH+q9/onJ+PRpEedUmW
bDpn3LaylegAXiG7aK6fyVN1fmGxJo73/PgzLQ8V6irroM/LZk8lRhp9Ou7ri9/B
wELa2IdLCBsnC9rMK//SEDPD3oZjrdS59I39L1kfhrp6VULIPoYvvBB8zqX7P7gQ
LOj9AsYK80ICrIp+HTx/hDy/2SNOd/Jtw8szlowjbiNdQjI4cMBBA5LGdS2ybGNc
qZLRyPZvAy6C5tpJiDuGsfQj74M+qussq2duFcqYgDqz9RnmUWds2Bg8KcdTRajo
5kWEyUP9XuSzThN+fLdSmIHJLFRSwaIJankwTfDJ9Gn26aa2JhoMA0qMoRMR9jvs
zyKUOn9KM8xn89mXny4qGbsWU1Lb1KksQRWgD7xzaLucabbAMbI9M2baZg55ebDe
u9R/bphGjS8lCrqfBLbDU+unDWF1LSlDXSfXD/0uSdUuOkpuwOKxHetzQkODwgT5
PEtT9vYiEORL6l0351uaik2f4i1yWGL7EwuyIqRXbvdNuBREAvIsd1sxej7SYQSz
XchrgvPZNqcCcgivSKdn2Qk7azqenBoWt2FX+I3OP2O6EvJuigo/cv3HCYUKWPM5
RWO9ZSsZQrQtGeSgetuuJbcUOiJyqJj421zc/+qiyeG7FJMhjz+bLQG8X07oGKK2
lRcgTukhu/h3Rxx56IaxDBj+7ex21YxuDXbepPaueuW+nn/yW6Vq9kAqrEFxbrVy
R+Ys9IBPkJEtMQYq4zK5DNyr8fGQZcQBTh/n6EmhBXuWAJFS3DmvCghJPfLfzRou
4R1NX7IOXHepASsg6FQRxR43JTfYROulJY7fsRMQc4l+t1aDnjU4AyHP6MJ/cm1X
NJEZg1f0VSTi+nyOoLGEhz6+9vnPTm1dUcMYaj28q3UcVEhVbtnZ7aKWXYfTwasl
9hy7zY7aNMIwy+AR2rrD6vViouQK2w24uJml9iumGdrBsOYa+yPh5gcrf9iP9NPZ
u9mLZsQvlDj5cX2arPyuVE/O+I/1FBolBa3UZKN4wR6qsYLPLLankvvOUHIjFxly
/ZS2Qatr9pg6VBiEiQzPjP3PVDIbEZ7d/35oga3CbaDegaMF2AdJTBbBbM8BGcty
BegKBZNZekofgnFkI3uiuhkjKZrMa8gsJi7B7F9SPP5wq4z77cxOCGraj/XQP5ZS
khPMWFcK03gZxVS3Hv0leztF+dhC7AialcunZlfEIn+O6MAXs9Rhe9N5O5f6SW83
ZMCUCkKTHVSHW5bDlDkqgwT3juoX556vnnRaDaLwPFvYMa7zSLC64BBrFUYEFwtT
rH+LxFvWXG7VtF3Ip6pgv+vmW1nu/dwTitQsxjaXqEiaZyX0uh7FcbMUPszoiyOx
OeFLzaJCtyMgRsVIPwajnvwJndkxuFilnhImOPw0e10E91u/TZpjNjOV8Bqo8Jgt
90LA4qAXiw/hb5Fb06LaNs6bCt2hZaI7bLLSfDDpoke8tdUkgM/5xB7ALFoEfXW0
WmoYixaFR/ITcp5zg875+DLDRDwwPFxh9zBYZ4vL6MEGl+VvpxvEujQ2ZfSUzaCB
mr8pTqK2aVc/pV7fdeLG8KBR8d6XJZJvoctWvTEhS+LGuq7J1jPnJCmgeUdItFZx
8g0TI5eZDJ7Oj+BLnOWe7Qe1pcv3hhubqNwbJ9EBnW3jdvxhnQteq5q3i7FDBf2p
YXHqYywe4nuCpx6TBjlWJxVwY1hiXUoG6JNPxMs0Q5rMdVl/mWIW7nIYqXRTGcKA
SDvqlgP1BsiqTgj2jYVWNticIBu2noLTUVge3IjKPtMli4FXA/VDn/FwBtgV0of/
x03dIoM7a1yWDjOemglid4UK+IHrpul6CcW3oFMbAQNx1clo0OZ/+YyW3gbQa3yk
utqc/SkNPyraoWwC0r4iq15XgHFrM0L537iGBtdZqxQO1CdEiOPRzU0wacbeLs1U
d/PV/E8TnoQtRz07o/yI2MJrUZ5f1xViXzKzcM86DP0sjJKCmJHBhL55Iel2Duqr
axAFDFlVbuOZmV+AsP9pyA6t2snP2KMBR0sO+VAqxYUcRgj50wb7hDnMAIdxmSbX
aLQP8CRCZU9dZvl2g8XI8dV6Evtph7D/OF4RDOHqbPIz/kvuysCp3M7SYoU7cbTz
uNWzGIQG70/6JERoWmepoWiFlMpBDRTmnIyY2rB+Ol/Cp4QwP9VEbkzzDFaAPZgG
FzP5LX+Es+tZQMeJ2MmnLoOqo7UDc5qS/pNiKU9Y6/Q2YTqvp8hihVZEGhF0U2B1
WarRbLUZBMLcDhYAnCGCMLF1QAur5O1OvGg3JhhOkEqrLGI2KPzMGwD9HaHuTbb9
7VxiPpOl3FHsMGwDAt6h5BioVQ1eoqmCkHu5y/9peeQhtqI/h5f3o1jdrXf8l5ZT
hCPfRs7GleoNB/k1ykF3dFh8lr7K37N3kCzH386h1RgU6qrTqMn6DdE0tjyozr6C
DYYM7DKOfb0Bq4NdJWnUz0UYjsUam08W+gtCW+s77CTbxtyCnTPmFSxNkg1keiuT
5E2hDP+Hh6DZhu+tRxobXwfLcMKJbDZ29/Df8W3nZwInK1UlR7nucfkiWkHu+dHC
JpWahHqNfAzhOfX+pyg2I0fd/EHavGx/cBg+eteNSRvgKWz4jxyUmpQw7LQhJdDk
n8BedAaXExNAusDzTmecedYqxgKzIK4tLIgwUvUIsD5+/jByZA6+UW2/r7kGj0kk
jmpa03AufWyKRlpFs+IN6zYssoOg91m+WNjXi0xB7e5Ap0Ex4eRNnEBPzROmlzQE
u017+dAG0o/i2YWUGNrfBzO2EvY+HrE/N0QqAIkrLBdHEr7Y72nlQ+MqT47c9eo6
HR24fuBSxO7aul8qvCsDZN8Y0jnd2lZ9s7z6c9HB19Fq1L7LJFYwJ80sEzwNS65g
imC/AIGslBJwvX11AK0Zz/52H7RFZEs3Usa/LuKtBdMH5dAW8Su5u1dNtoqQw7mv
rmjiEN7yzSXQIh2kSl4zPuoKoExVAAcLhrhSl2JkOWDfWxodAB9Xh/H20tgvg1Tl
ptYy5IdDbsXuqaFJW5cmVAC34OdDv2jwBOFfxxXlNDiS9I6qMXBE9D5XQwRYXuof
hbeVGHcOqI4FYLuvNHmLkrXvArw2zYqPkLH6BCI1bxiMWxMkuYceZeMII8+ayA+p
lGIZ22k8HPmGYGJeYEBiTsay5CUzfK9LTy7JL3MmMsrwnasbLDlZzBstJJax4jKd
apnIVfFzQHp79FTYlGIOxU7Iq051MLp9Vvq4VCLsrCZKqzB1XXKHvFynEbGxHSGV
ANivKTR/M/PldEq5rxuHvfHgPZwo3KiJ4dJenQb2j0ltKMcO7ZOHaQ8U5NR/cmtN
oWGl8pvbsH/aPWuZq3O1K9WS+sw/VUacwPMqAFnBpJBipM5rDaNlgvyu0HylXSlr
r/3dYMZJb3qpkvgOo6StpbWdeM7rbLktYJjdoyJJ1gmHc5k48FiicMcdgkHwDa9v
MeCC80dXl7YBdv8nXocVvswui59qe2zQhJZ9hKAixsUcbgMb1Wo1kRemR7OmclC/
o9jb6iRErB8HRjpELcIatxCOER4dXbQzIVG8iIE8dSD2brq49xfa1z0F8usXXzsx
UI3K4A6yxfwerqESsESgTvs2tKuPAceWmvUna3h1WlxgOCd3kN+q6reWlCYgdXGj
+2KIOidlzp7kMaF8jFDfSCskhAZhl+GgtaT+Ub+2oSOI2fV0LTfyy+Hefj/lWDz5
wknwdob8/Qmjn7yPB9JT0JI+1cedWM0UmLaqZSzJdbmMbwdL8mSUzYu/DQFPie04
Y8thdc+TYomkIf/QXMPzV6RWb/Y6RkVG0KcMSvX4GYFsWVa0GoJnNk08paPLkHLz
K+d98ueM6DSTs3l4RgtXdBk5SBYYtfWvo/qUa0HdxeKgXDVZT5Hzl1odDSg/TngL
OwSzsNBZCsqzaIi3IAt9ZBPKJvFGv79QdNP74rjBVNE2kqJt4q9aWPMSOh2a0OTJ
R7yAdHewJdoh3W350qnSeynDhYlc/jiNtA9MJfNdUgfWtkrjUUTGs16cj8URpFx5
SQICOcA0XHrphRBkpdJ5T+iRZVrdSTFnfeOmDTPSUDqqPyVmce0eYas6nmCHtseI
HMbRj+fieQQQqDACSp18KJH4xHcIH4gXtaYy3Hinaa6/L4J3Y9uGEcsoNiSJe+Cb
NgoRNt+AYbjE55ZaZ4MfNnRFegM9BZ7Q5kUoc2VECgBdSjCOd4lqcCJnZcSkD1j8
lZIjREaPaJ7N5RS0bHTtTWMIlOSneW4y901renKWEaGax/FYJ9cihRGe9INOPBvX
golDyL9fOA+O5cw6z3HIQJOuA8837MIlECVTDc0ezc9s++rC4F66MiALk6XzGBan
eDd8+2t1BsJF+VR/r2isDrMs3k2yA3KBA8xbGf7hHoNGECZnhyBNj1YpcIkXDbA1
FuZtz0yVine5pVcxbxoyLAyeXXc+WBj033BvtYr46fnUDB3k995F8tKkzklaaXiS
rN1jF4TvJSs2JvA203gOgsC/0fWmX97emZwmnu8uWkOTMsUUJmUY3q4AI5inU9OI
c3ziPTQuL4SKuaNxzUV9hIa4NmjYTMyon8SkJHpqod3qU7TxFXuJ0SPBmDWF3rbk
FDaHdxeg1KQY/nlAqJi0RvwPJU/O7ODdhWszYXyX6orJCJmE3JIS8EFxRRJAwUKe
2dBQhh4CyC+jBZ8TQQEo+LZjRzus9vYsl1RmiuAQVD50ntf4AwIFlrZIDq3HbpfK
7fBqRfhon6bgFtNJmDyE2Nw97h+UdQy9QSKfv2MBZb54cBFzae21WO1BxdV8qrnO
+6tlhDfClCp5pL8XV0s+gRyaGdGaTBaF/XNC8morltihxNWIiNaHzP4Df52lyWMO
i93JGgzMvslXD4TVsin06es0IOspJI+ubB6R5EzG7XH5oM8W8r9vj1PRXWB3unlo
i5kMpTyUOD1xkjqCPuU/FT8XqJF3O5TE1uJXDy/K1h6S+cjnGYIA3Fw502EYAAq+
38QoqIQsGSh1EVuC9GKpo6nI1f99BhehOVNm4Y6qApQ48IHZucZriAonYKgrz0Sp
xQzJo6yUIXo5fyInblk8TyMuDHDUK1WcIYyzqu0zggOI0IRFDRyjXUmeblMOM9YV
p3Dw+Pqy/8hbuIUCdgVxK7ul2seGge3tPTHVlax6l3kuXeFBVX6GmoOlOKNMEtqH
cyAZW0aIRCbtxQE565MCJRCGyd2TQ+KAVPoklzNpcyGCy5+wEU679n+2ZPUCTGoL
UZIWqZu2Bm0KqiiqVDVfBKo5bVl9G89Gxeb1niSd7+OUGFqwyU4mdv1xv4JNfE7J
giiv6jk1sRVS7AiCv1wAJhCq4iCODh6SYyONKJnB2wvcXM1beiPHDatl3SDtsnn7
FjG5VdsLuPfrpFsP1IUGiBHhxep5MszJji6ZxB1XSpJykGxQFMU8Qzgs7O/8Sy5t
8rA0OXKWVuYPhrrFAtHnu81YyoxsoNzAgLnYz90E1fbviGnG/2t+ZqjuHKk1+Lag
qpmUAMCwxBEw8yg9+tNRtkQbaWjZ69QvFpRQUf8yztSei/o6/0mRJi1nEU6N4oNt
LxNTJ+EfSGndPdf8o1l0mLC4r4bVuJ6mzX4fW2kYqUEb8m8X+V+7DVR/kSQBzZA7
nzrhxuXkyEeE6WMKm0CiApisnnOLyoXLoimfX2z5rdzh+d+SIoT+lPruUVXHAWHI
2/GmLxc8dZfHcbBOc5UNnU/0wKX6z6rMf2fGqxeT8yY87cyPKJqHUtvpV8S8+x1C
HbXGOnh/xjj3e+PKdQQJsLi3eB5AjFUOOlgg0PM+mN2OVPetbmcOZaLR/SX94EZH
KnnjYtT2u0TROjpYhAhSl5Gh9F+1hhMfqFv7DpfPStnAy0aCMb9YWgT3PsOztpQX
/6bGuV3tnngkNlg3YyZZAeTHmxtj5w8/8MsS8Ohib8ddzeybEVKRJEJGF2E2UKwd
s7+V15Z19VAldKr6p7BLbRmPAdwKF7EbLXdzOdzSskqU37PMWPApVkIyPmB5JysD
OdfX2Hh7sKrCZ7cGqZFcF5nNJNIJgNcWnjpMokrBALITI5yNCeOTJ9ZnJTooehVN
tn5TozFmq2SkmYirQECo3gndut+5LywodM9JL+xkRa/2Ifwfme2d+TRxzK7ATU31
QOMm7FZz0GRGRyaaqfKKsDJqTbJArxz67ZVUhVmBrfc7y7i7snNYoJFH0G+KWHP1
/lBRTmSXpuVI8teio3SkKNSo4zxL2cfi7ISOHKmgTK1ebsHWzYdCANnsd3Rzz3A2
ooYocIw2jwSywErn71IsJGKT0BOb9sNYYY6rZszxfczx340lGWPuwpDEO537QM3U
ye93d0ltCkr5W8CSl8Irzn7y167z0JPbfVG3Vv1A7uiVoiQH4n0ysH1ywZiEXFBq
J3RLcG8Qgp4Yze6olYMBKpZF2xj43EY1qRTPp/C9WcSLIt6ztxxnH/0uctvGWo6l
lNPF+RVwUlbe6HodggzCC+7zCcVXRkPhJmtI1csZW1V9wsW/LufZQwfqTzdtQ74/
CzsknIfZcwPIl8sAygArfU6zkNbyTVCpmOi+HWWcUU8wH1cO312YBeeM+r24Qj5q
D4VcBck9O6nN/w6VAMDlAmlmj6CQY0HnKOQGW7Upho+TZe9Gqe+Ktn+GZa69KOMQ
nC+wwfrE7+n6oI9dtsG+LoE9lDTNpTDuH9XvaEBCOB292i2w/RdbXtxnkcDyhsjD
bgeJFYEjNNPesaumyHXwMtJ7IU4p6gFUZjfeSl9rZty6O+1KLVgxTfRQ2Nlrbakm
ae89YdKLHngLdjsQ1uHNI3GF188m3b3MkdSB/E3OrOpy907FmM2J92kvVm/+Tqob
MYbFOqplHR57jJ3gLVWJLNvpCPvH9TP4TeGvYhnQ9L+LE8TcEm/fVnV+ICu9spb6
65KG5UW6hVsP4tUsGa4sQV7aqqvIL7XiOLehO5x8Iz8YvrYJnR8k96A2rNehXLv5
hgy+gRNk0ibJVAXzVV6+Ov30kmLkBjGYQZYnTxKfMc655C8mfuMMLY5DOaGVbrB5
B/4piebWy3TmZ3C/NW5I8w6SRGx+85xWq0cuNUuLuPBhREfkn71hp2W/z6cHaG37
LqtG/polqb4vqGcpJ74Fq+s6bvt0kNRAbi/hl9SB6+WNIf9y3GvSUCNSkf9aKVP7
g+bhEITVW/iIE+j5/4269DKgp7zHM8jkS1i917XwcJCeviQrMi9ZDm8DKwmIIqiY
Qdv5ckGzPX0oyK9CgGYF837uRLMyLgwPx1bBX3o6pkJBcTRZmObOu+h3GqzBF8Je
ZvJMoE2+a9q09u9qqfdoGlYC6ThJoyf4+DvOiQMJlQOGF5uNZHBy83Naoqqnq8hW
jou36g11TBB36g7fSc3+y/ipsSKVf9nHu/2PQwvXk4ojU3yLIAXJZSk/IXYLNtX3
1SIx+f9Y6zyff4sHkvnOcu0f3GKVohjuaeOygQuJxzwyH8bWAJnNCLZfnGctgpnG
JL9PoA4uNsPKxrDEAQo57t0zX22L4MxAnruvjmH4VJMfVa6mEQ7eGeCLHrcA65QK
VV7loDCeX+rMPdscPdEQ1aZ2yo+R/pTeTfi+xdsY+RSVdgOeWSQZLnDFtltqoBnY
nQa+bQjlIh8bX8lRzeT6E8y2lPsBhYDkDw4Xet2Lvug0VSaujdR6MoW9lri7yZ68
BRuxS4EEjIpHsB5sjSpQHAHrS8L8ziou2z4d34NF42AfMlWCl3HcS8YGG1GGLM5L
oKtB6VVTwdXV1IqD7P6BCZgMG7Nfyqi487SVUosgylel7OClRN1h+XdXGAbyn8Jl
phmDeIjSXcG4UBKkZyn8X6yyXCRljmzGPioOFZzH9ylSBnGijFOJ2C3bWPofECU9
qy3h/ZeVse/ew9iiJUVl1hydcMxs//hNQDpW6wYSrjASiqEnjYFxjkZlBV4W7Dkr
rDkM8EEsrq5HVWlVD/RPz++4IhzKoYQbhKp3bAa0XXNAKpS7S+uKTDj6hh5nR2DG
ph55Q6dxOhMndgrINjkdwC5hTCYU55F4hoFHQPLyp9SBUPQ4XAbLl8PnsRuHHZLu
pX0IaMIwakvbdgTTIAP5c00FuA3LUwYW8X+BQa9/WcNxVINljIA4BF63WynKbIe4
9BFwJX7oMrn6UYHu8xceopKizSG2A6yu98kyO7q2hrkXX9GyzjgcDvSjwbo2jH6/
D924nKFeT4Uo9/2U0zOIvzFgmP63QRMX4A+IHMFrJnPfi/N/Rx+xjXakyzTD8RCk
VrskOG+Pfco9CTou1QhL0hxz6FMC3Ei/hls4Gy078PXWJGoBGHmFmti0rDcEZ/SL
wPFcb8AUN/PZs1ryh3e/eM5B3eppjka+GC+ErjjPDaMLaruuv58VF+rcCusu0aId
clSAqNUNBBaizS+9f4s/Mns1nMnGHjE3yETyKAEJvBqOO+It4dHbj4jM/qKvzH7i
AUx9N7De9rfZmKLgMnzG7LQEWObktaSj7JUnAB7SZZOUcrQ3OQpgBzikOtonC2K7
MKMEaOMbWmXXayfZrLZhfIiph+XIytfb6oYlSduuCUh6Tu85Aa3O7DI6S0WOC+Cp
BtieZhxo4S1v34DBi5RPPbEqQfDIhXSYiqncjji6lUCncNwlTE859JQFQvjusPTe
AxKfy14Zyn8GHv5yTYZHesb0Vn4ty/aRphpuNggm5t6AGVgNDBCmpUE3KMUCsORo
jfYbYA/+pnvQiBvlKbMicm2ENd+EjqLmCBAQD18BFuxGmd1V7N4yg3wbiZPQwsMJ
+85eEJ9LlCMEe+e9wEXvqCvvTNas0Z+tOcZ01thvWUGw+a5fTsOTd6hvWRg1QgtA
0F2vEa4YFgQWOTSJ3ij7GUo5XBtukD9PTHDoaLSz8gumdQCfBNzdUAJNQveuZF4u
W/cVm7o/7MCnDTlrEveXR4n3iMHIsczlu7HL1OYOXpzcgc08k8cYyC0DFTUneU8Y
RVZA5RswhE7zWEWSgQnt1WF8ekDwPfpJs05IsOBJAelou7yWsqhZEKLM9YgvyIiq
GbJKJVFPWT8gkWNsFehyWlrhFTw+QFoSweEgNvaL0mekTVhW0/nWWFUktpZ7uEUE
oy4vlsB5X9DdN4cYQgd7mKsnglhZsw6vD8GTks3i8izYdyavQrfku3fMk/I4T1e6
W9FPA0Y6gSA/Sab/VhaU+3mYcBCcfhb6AlJGfqnxreubELVRnPS5DUhCYViE4OPk
hc89wKsHVV6xFzjrZHbwF9mrQKph8KXXpBy5c5/4cSmGZutc40zJQbhFu7irPgFD
VbXP0BIxmuDgBUyT//JEJL8G7dPmEqP+06UGwttZ3S3jzQGkrkOM6Fx/+rQGKCXN
fISS8L7zpbZ44TbsdyqHdG+42Bw92PLFgJ1VuVEG+QTnY05Q7B558XY8mg1s9DJR
jRfUYap5VZfaZrIL7eO5dHgdXHpZb6JtnRFOtKMs4QIhSAsWQZN1aBpY50LAFN+x
7pX+VOMStcP1pQNnjRS3nqMIn8v5NSSj0VKFuEdnuZ0snwaN1jFUiJy6EtnuMji3
ftUoNQr3cKFfyYctsySK8Dd47dbyXfS7Szgxi22njfMCyxKzfZ35OT8LnEmoGVGv
kRRyqwARF9bOEndyez9KgSJETKwy5l4HLBeL7F12GM0unlDvUMSI/hSySzfAK/r6
MzG58lBJC9RZuSdNEHoA10hcUDJ8gfYOd4IpUQzYfiRDmwzJHVX9CtmFvFbcVmwk
lmDKrkQa9xkqowuUTFBiLqdLH/x3SE8Q8K1/a6YzkQpwxvT7WtUTU17DpG3B370o
6AODpQHb6PT3eYuQqB4kmZEjgW3qRHICEBu3zfBM4tVuW1zA8Kg2Xi/7939Q5b+W
vWco8qdTP571H5ZijZq992U6IXZejbpT83Dx1HLuWa73Pufrvg49e5DR/pC4Yp3J
+dqvbGLgVTLkTb4cjnP1kYwNIgQF3PmOPJ6CprzEdlw8bJn4KPG+9whiEvqzC6mD
S1IoLL2URfCJUPaf+dY+xfGAg81nwocU4oIhCInxq4RCx8aCHJWEMS/jCfQeWdu8
8N+wnz42PDSp9XmR1rD1vT7A/mhSOV/USfmgfa8KjXcYYTDDqQ3I9vuS9I5qC83j
CK+ZsvilGx1Em4qiifokvzanzozRiwx/6gJ4G+7J1J8YzrZN7ASCGLOoEOgR7tyK
WokxP03Yj8nRrjYs1MubRw0wIakrwxUXt2xPoJq1N4H7UMFjcUnpVGnxHiioPevn
w4ukgJnYomrVpmXGcNh/pSUYjNNHt+bKfTSTfrBOtCaEFc9kCE4yjIeEv2ohVcSj
jPvUPLCIBMm2y4CRn1MXUZiq3K+6LdNNwr1Zj1W/Eo0G1AcUCzCg8+lVMLC652aK
KGdkqLlmMUMbUDoWgfgnP+KKId10VOEXGlsCAg82QkU6iqWCwwW8wuYx6ls/eC3t
BAT8aTTW4MXsivkZMTJfBXnGKEH6XFmfS0x3jlzNxxhase4Tlp/c3d3Iiks5OWJx
86ppSPKtbxezK1cR95EBfwM12djVHLrgNYHlURhmJQYELVjLDTSth305Y/srsF7U
BVIoE/4NzgU9M/kdoENxaE8luoyHCh3qxC63Yrc4BkywD2/ROvqAbkteJ1epyRom
aWiF3u1Ecc349fxIQd0MXbEtNstMJgZr0jN4bDSLl4lYlNrzURpyl17DvXjymz5i
7VfTr2SUi12Crl8TVMperz5c0BFFqW2dbxFxX6kzxqBJEGLQYlL8o+9t+GSwo2Cn
Xpd2rYqiAR/E5GLJ8Rk75IsY8ffB8udESx4N5kBe1TLnvfa2Wn0v0y/MwI8gjHr4
c9dMouwEn7piqWLcjO8Q18Jnb0GXBTuHfMzmHpRpvxk8eeoLTWBwp1WVwzUoE9Ch
753fI1Sxokes8F7oYIG4teKzMVQ4uetHoQuMy48dn3D2eHHD91C5O1dTdNSsarqh
16oPM4LaWhnKzkEdxQ2IEYBo6spWhO26+xklfwGQDLgH3qwsN2rPaCr0iddy17Vi
AyuXtmb+GcMD2QeBRnel/tkbJSb/9MZn/GhsnGT+9/Skn0krmk0ZVdEiQ1pNBhqG
EuwScX1tzT7Vh5A+gHUnpH2RLMdxFT2NpUm+TydWS1uK2mYt00B1UC6qwlHfxnnu
iY4b91TsqWr0AHfaoWpzw0XyzyfA3cqGp+LFF5QQvJw8mJS6p8lUTzh4C9BZsRPX
3eZq5slXH68jZsXS+heXv3Yfn9wbwRvJq0kEAcNyfrf0Q3DXNpJ2XT3N98g61OJ2
NEavAKCIiGy8jGB4zoq33H9N3ba8hJqq5AIfZZkrbXycf3gotqS1welpWfHweLTw
XvbDQuUOP8ZKgCsc/poLOejYMTh6c8iNokEtkOOkeRiNgBseSxWmO1rdX8uFBV+D
jo6IazaE6EAEtqxNWmbZNSqjrvcmvA8mIaSv/sYoEBchQKRa7sYT20JnuGyZ1shZ
5SYsOUFJOiRf3ZWMqb5g02Dzem4ad0Zpayd9hI6OKmXSD4qjjzmzxVxVUmWkaLzR
x5E9hwZcbuqdDwgUYMMWd6DiNg58J+U1DdxcvBytyM4/jbeVe/9qR794A53gdryi
j5DiPIp1sJeAIaczjKBe1r3H6c+t1Ctk6NoiCS7LqdEp5bvMBnUPfo5WTyu4ZrKf
EkEEiS2AO5GPOkOAwE+JNKiYEqUErK9HR5q4KT3LiExTK46I7gAdZiqB/CpplGfM
8zKNskx5epQmzg0WqjDOTMqZABNs7+LvdG1gt5QkTJFpS2L8vgW8i3xqVd782Iyp
p4t/tGctbmlEEKyl0u56SVkK0rQbqLoLdWqYltpie9Muyxm9kYB2b4rUvqhVFC0c
ONi2qMbkh82LKGLsPzxCGoaCQV65RNsskq8OJtCLxz0RNTAgNnRpixhISdZk0nLI
R6jijBY6GgkHWZEC2FKdbgEW7HzVgDmgXbxzaqy1KU2OYwXvRrka4J4dYGgBSVYx
6V55AfG4kbhul0e5glBI4GChB5DNSdVVGBedJDRnuzVTq3CdevT/ZTwoOzPEGxdw
FNfIDI1FErRTm2TX7VVu+wf/3irSDqBHTr3llwBMkjKIJVLm4PNDrtETSX1RUzSp
kYmkTluF/qKXSuRu4d6WuwzmIhH/UHt+VXMNYcMSXDhFpbdejy1DQUqBDZFGOHsW
QYP0otEqwbjIzscz6ScfUjF1jWLYYZDANQGJJ+aEY/nXHQ3fWSydrQ7nkITyUd9k
zTVPbvy+CGMGa4WQv7hsk9EGvAWdcv9Dk4hRDOe/G08syLE21RJpCAybqcVdbeXR
qj0GbMzPgQe4H57kGw7/wZVcXDgDdfNmISIJ3HuU0xkgoXyqvOtuaazgX0CuFIeM
US3j2pp5N2IY+F+j0SZndAximpPjvD2sTU711dUyEcacd31l5UqEEvVWRIEAZdJb
2mfIHtNrJ6poC6Yp4c7Ng7xJBcMH8HPomU/8gwTNBMoLO08Sw9xzMcZNJj164rKT
Xp+fwT6icjG+RqSy/BCneLDs7sYjGrE4oNT/BjxkPyaSStnPAh+ZgMzGfL0GsWLI
CgkrCHl29oYZ2VhklGZF0tmgJhUJIiL1uNbS6SrTRMXNYkPVKYaojscyW2l6epdT
pNdvI5p4XM3PWhwNGRfymi62SfrFVMP5BhfdPFKg1wEUfFcW9MFHOaoLlNBw5DOb
WH0RKs87Rrd8GaEdkqClO0+UplFWmo248HUs4TKsfJd3Pu7MTxjB0+x7j89J9bBK
yjz7BDcOpne/+XsAeYZPAX/bSVqZ6NntBCeXmJaPufTonhEt0x5U5RMcHy9qfo43
AdA1mlXvWGYKTE/lr1tE8sqVfpa4Q13XGxXov86gxmsizGGGKW0zAN4vaFW1nH1h
gddeozbdqVbTgwbXvpJx6PwNCRIJ5MvgReKgk1hlnwPliQNEnrSXDcLJdWrB8Xph
q+NAl95SkdRxdeGQUATAhrsbkMWfW3mLcgZuZTk+0QYqi70oHelWWlIRLvTuQoMS
D61FDMgz6ROTDiKH7Za9DdZX4YjDTT7RGKHstpkIILecbEM/eXOGYECsNPLBRknC
5JrZwYjYM7/9VLfeGIKVF5/Q9k2kweqEPOMehJuBXt2UOWmjsoHKYhU8fumnD++9
lU1opU6OEGJTM/ojywxTkmMT2JwAzpdZRoR2gcW7/spJdrkysS1BgNixCYo4Ji4W
JHmICAzy+z/aNwStgUFkYNJlC6YmCPFFTpYW09C8HE8n610830OHSxmdgXorqqcQ
92e/5GU4tdJZxFus6CnglkQ5OgOM8FhM7/viN53XDtde75yNvpifvXG3yCNL5JAx
9DxlHq4GAIjGcdpAzLuZXc8uxy4lRlzbIEoj+pPaKqXq8H4lgbGvdPT/FDvRNtrR
SMpBeVqA2dboAW0aK0uY+vcaThXdBy16h95nIETmAjEfwp8j+vmGzyS8zV8wMDtE
Dp2ls+ZJzlEJuq7r68ecPFSt+hfm+fuVEYW59leb8+GxGdMA7Zsn03fjdBgfVQot
2DhGNWzjCyGloQbd/LFWYiB/4FQ7qvoW89ATaUjef6/KgSWleNQeb+ZcwfQTw2iM
vOg5IVO592ockrvHJqNP98Bilf38mZWFQBw3D9XM54qFSmUwGRJLW03OP5DkKhBv
QNJv6wvSb+cSctelARvElPhctXCRBlwUACsveCYUkMGDR08ivesr47hlTFOQDkGs
YRAJwOnB/XRmCcEJ/O5RXGxnEdUeJPc7vTiZkprqul0K8qBK/EoBxXcbf0vCy6g5
3pbypLjgmq7L9FNGfKoklF0ckzQqJOSnbeN0mYjNpRjRuRd8TmX5ou+GUHhujGFu
S1+2NqIJlZqCUQCaNtUKT1a/cdmnehahjosi97xqf30Db/mJFb1QtGJK7f6w5LRm
mK/TbFtBePACD/AnkX0HnknDBvTrTDai8TBFrtC0raSREc77xB1udPQ6g9psdxz6
V7Erqzdc5gzMbKeBore2cuzjGvP8cfXXouNFfVQ7kzBG43uXRwtNWqaZjy4sfUXF
WqluT4TD8cwk2uc+vHMbmbsBN3cnPeZ2PT0UmMRJ9DnuVrZMXQZLBQNmUhiAsQE+
OwItXAVxM9IuZqHb6bXpc99gAP8u4gaIrHidiRZq+Q6rCzh/8fn0OvUjvx+I02vC
iJLa19DusDno3D7gQEP4PQop2m4O7HgsUIYRgUY3X+jkXw2c/5FGxOmsD6UYCdxH
xmFdeIs3gR25aEDBbjszPWuAfWlNHUgKw7tWU6uPWYHUdqAxYSsNdtPfQ4uxHGPG
dTFphJTD3Bqr51FkrYnNA2sz7yYsVsxtOV9GOmRAIQojDBw9mXellyzdhejoHolj
O8RGfXAz4Q8FQ2ktCPwRjqnrcgC6kGA/HhMnDQNj+I0cotyInAyC++DXaRTuTS6H
a5+ZQ5Ry6ExGk5AqBtk9UE5t0eT0XbU632DGK3JRYSolTEZEUi26/EZ1q5GrWN7j
pPLMYmo2cNf+hybFe3zpcKFnhKraSxRNRAfMR6CP9VkVzefT9HkVX2N/i5tO22nH
MjLQg+pmXlctp0fQs6v7yTFPRdpzRk+wlCJxiw4naTQvwJUCkzZLo5/wtGf88uH8
+C03KndI2ReWVqvinwn7jidwqzr2f7VF8JzjBiwVZlJupNJ2dOR7Te8FWD3r+rAt
fzlfJZ+maztbOmoPieWzsRW6+yGOvAUB//Hs3ujMWHChQqt/spxJGX5tJSRAL0WX
nXu0CuwB7ajHBE4z+NqpcoiklA3KTUISm9CDU40qw44zyRcSxmgA7m7QksCsSX41
WJG3eLoAgDH8KQUilOSIUsZ6vGob1e2ZQTPEBKIsa2sIPmuGwaSDNch1ivE8hdQE
ka66+PKozIinMVqb52uw6JYLlrNmw2KZqO9pm3DK7Z5ujpEPwfUDa1/k3cqtZh54
2LMsatIRN+M5V7JwLrocPmJqfbpY/I0fs2MpUKYE0JjYZyGArbMk8l+P60lsflAV
gO6yCyfCXlkTbycnkMqjiGdlgNiqNemklxrZeQCN9un6xqHShrDBm/x4WrgHtBk4
CJjcX/3zXnohqDSp+RZpPVfg3AvxBXOE9B1OqwPRpW8TejzSnWIGTgIgJXbVzZ/Y
CsdH5GF1wCDF+GTReIphPhc2fsDNUcD6lVcVBpmcpjWfMqFVJmhKEcTFVAKA6V4J
rVHsT746llhW89Is9M8dZ+cjFWaBwp8rqbCPG2MaNighvYOYHKLQ79SonxkXO/ok
rJ+Qo8YJW7ezQJQyAY+NzhkUeGN0t3ajTyzds6MOKxVCgZHC5UyGI7nl7GLEy4C/
Z593IHhQinLE3Hu/fInnsOzI8KTGJLdj0cuEWbjE8095epMKFCsyIPVCBAxqsXrJ
m3TavOTLqNCm5PuoZIeVQUPPIPgA9+nEksHAwJbZhH09PlxS/vGNYlcSF/wQ15M1
FJUcTJmcj1Z/2RpgutpETl6lqs8BpEFz7/8jZoJeOp5nkBCpMe2tDss3g2bKbm3b
FmUukKwBKtSpXpwLVAetxyF0NSlOj5+QY+tsZ6vKU3aGPMiVT6i8T8c2/wtMUm2t
hXEkEQUsaObLqqsJpA90mdbIxUQfdokwD5h4OiLkxLIZCa7ZIIPsI6i3XdaeIVCA
fXIEwqqOvLctxU7UReq3GQBxqnmJdxs4EY8QpoGMSW/hrRlAHkdJ3+Zc3qUsgYYz
mEjhHpawg2vsnznbLk6P2PN/1Uy7ymZgq74sC/oAXDqCWWYd+Ktt7IJiDFRPpN9L
YwNQofeg1et3j5O2DjTcqPC9mC7plYKSvNLjJOr9KM8GilBYTb1wybp2drOw7qot
fe/B70Pat1DvKuWvmZD4yD52Tr6gQEivxVJd0kJMj5/A9jFEX3jPoKUKTgUT6K1z
hDv39Av5xlHY8NQuv83SxJhTmw6BChj75YdyD71mQg/ZkfH0SimNuuto/dZfDYli
I4HR3ZePfE2wKHFKXvIGPE3Mih8a9OTPbm/n3L1hhp835Qp7euju4/e/iOKizKDa
3atZocYLZ8mxZNhl8zj4c6r51hjwxxaOfLmAfqeXCeQ9DW6jOomvY3OrxLSYShBn
qLw7vkgDXvjQOxBzFAZQjvVBHctOrhmMN38wImuhckiKjZLteajRi6l/7MljTWZw
6qlr7Eh4EigtMaYPbh/TX/wUkpiIYxj0UVAQlucT/6L9LT0uuSI4zLHP0zeCU8eF
ASPhgRMC4t0Pvejoobhs45BjbCdTXvUMQreT54Fkv2zQp9LDGUetLM5J0PzL+myT
WyfW4zy1s68pRMQtww5dW1+VGG/+RykBkXvNB8abI1SMvet0kH4qOgtuMr9SX0T/
QTRoL3k1f8gdJSYuIxC9AJQVhXXyJhYKbvwRhCzvYBCabQax80oV1Ra4RhqA+ZFv
sCbr6bHJyIGwQcAjYZjxHu3JQnfMR37uFtpVyQeYteAwWA7z7i1b6wvZUmcs0mA1
cVyq++oEDFN52apXDkMV5xduLvmhmhXiyo6pWeYp7fBNUZXQOQqXOJhGDMm3egHR
MO4Vt6R/cRtFnDHbkSXZH96tkzemp0jMTzzPLtthMbnwQdohHJwIyxHk+LiPOuFm
rqSVwJQiwEmZm5I9pWo8YC6VUBzl12LawVVR2xUqpXQ/HN+2XXyNcinUoBtq8SEP
O/Ibs3hbuLWEvVt4vc9/+vAB6dNZ+Z3g5CWG5VItiGcqINSKPlqRFl9m+73wWl8z
EZU/nbC8aY7aihnzun+4QWazD0YTtgXiTlwzbwaK6aOd8rRCC9270lKOnKrQ2HDq
CKQfqIAhUcVu79L48bXTvCOlGxEFZkT3bcTnYtd8YexzaxVblCZR9425gILq6baY
56D0weewf/6B7DonGaJe7JcxV/m+aMy/qJyWKXFMIkyYsHMTxGSbGRTMlQoyYjCa
KbNQ+VOyaNo4smQLueJ65DnDHW9+mTfI47b2elxbqcIdiB+RapHdMCaUQHhuWhN3
OYq9/voYrVn+65C39V2HSt0BKQ6fZDLe5Qzq2XizgV5LH2MUKPtBgFe+MJOhw4Sd
7c9YPbgjIHIda2CzHfbu+J8DJkQdLiM/OER9VyWj6OJuuHSeUwjn1AKwHHxBNlIj
//3Mnff30SLp9zk3IzIuPz49tZ8ou7SjgGng2Y/h25t1upLGDazQwBtw3qFTqox7
dLY8bKYZYcgoe/5ZTDBxNVVxk21wKsQy7+jJT7aBT6ewzzE0QkRrsTERLHehmWPp
TWoxOZ/9LhkyKK0pZRL6qlC0r17TC0eH+BMG1isMwoeijKafxF3dgGzLqBIIbLve
jODqx0R2ccnkhN67HnVu9EN3goMnTtiidERGMhCfV75PmCnXyul97esI52++sX9+
Psag3vFklOjihXPRrCx5Okyi7E2fubBu4k/RrjDrYEqsZkch5n7zhexrqmFxUpRr
2KXLAajCYl05p+y4j7YBs/6eu144tyIgJ+Z0i9TaBeRg8g5k5Msmoup2h/prUYuP
HUPV+g5Rl3RgqDs/UW0abA+iUHlgxUYFCfzPLBtNSJiTeI7BXLq08Itxhf/440dM
yepctFNSiIIXilqpFggiBuVx1B2yRYlbdBS7u63OiQ0eldpAN5oFOilhiDOQKYNu
O8HB1KkY7DBI+rJm5chzjRHjqKluvrj2ohYnpV5ItXVozydtOX98s6+m7Ong1jRg
ke+ORcbRY2gcFQa9h/zWFdqPDgofuks5ckoqCJFQmw7DIcqh1cgbnp22UaJt17Kt
h700ZzeZCvy4FS88vxZ9UCl54r7nBbSbc2E/1FiNhRaX7QopUXr47JYVGTWx0tlg
BHqh58Rf8KuRQJsN2E2nBM5trixV8tcCWFd2hfGCtShMqwLeI+DD+tiPs08yDZOp
+GBp4owwNgWrXbRFM8Qd2ie1SNajsc5dTFiYlDAhgyVZY2v//2dxFYYaMLdxekN8
tJ4jtkBymCh7G8xW2h2WEan9HLbDK+HMyfTHepp8GC6s1oUA1trxDFwr8iJoMNig
3XblnpTyqjj+0J8ODSo6MBjyhFlNmY2Lo+Jd7rekUSbpPy6tl/USox1QlApocIJq
mQeH3fTwDoCJjtIqzJ4D6vjRfkQ/2v4pqwNuKGwzJiux2+WEbAM4Y5zkHfqR+8Pn
xH4ZHDMyyH+q45H+an14JaqrdlDbbR5zTIYM90nfPI2dX8qIILKKCp4/8/HB1QkX
olY/5U97Lg6YUT54Z/HvBAIQriV/dAsRIyM6gulU52wsohO47n241a9eEzd5Uh37
dCTJgygLkrYC2FmHGWK1UGY/NqItgqeSdqrSZGM+jDW988Xh3pNn/wfL32OYk+Pw
kxaVgrksQln3yTUiBHIxmwnxc5ojZiooxnuoVnmbc39zx7kAozwu2VGbwb+5ZRqb
UC+yQszowEIvni0IQT5QVV0sFj3zFtwI4uEsrGTEK0yMhhvQKFQQ8TWx5dnaDYQK
9wbNzdIaGO+LIEaIQ2wiWxRfS+mmJGH78+UtRDAM7jQsueztValx+xmAIKsBXx5x
stUEZWlKRVVkaJ4aXBZG+MGRz7ekPQ2LBptfTSYSW1PzqlSWneAL01FfLlUkWJzp
1LyoEaqdlKLMr5L8uyRF5T5aBeUvFwhU3/+vfF2K1Vzm3EqyRrPkpAlVdZ7MI3qa
RSC5v+kewIe2oVzyCZxotorVDsVX3P2XmzazugtjJrROHr8WhDtsdfm2frd8Jjak
b3eHw+eKs4DWdbuu0uwbYlkEgwrdVfBJhfg255gClmR4URIbhLKnAxmXAZyfewnX
52nzLGJLaJLscEuad3+PBBYq/2oYLA65zOFtp74B9g1ZW4XEBEhCqDNrZBJlciL6
k2o3zfMu1bG6+1cdxv2sRaGV0iLNYlVhuDvXQ8tIPj1nrPjUlZXz4XL/RLbmkKcj
CwaMJELiPclKDLufEjP6bzSb7giQcGs1+w52PIFiQ4V1ca2DFdaZjBo3C+n9RH92
d753vzfxJC7p0MOv2T+9qJEvXeGB/fvoEE0Wp7hWLcTqVFIVd58Nf4t6LMNInRji
mDTheCoTZKBFE47N5Ml+blVXy0TVXQdANBgbLPUS5qGYmTsZlUDfvadPiZLFluoJ
USeItBlPaqf73A0oWbTeQl9I8mcLUhzb8HgdzXvLhbGIsY8zzHMt5Asa64qzILm+
lLlumXuYAenBJT3qyLLusSeLE7/zSEIR+SJiLhtYaPXNeg8JHc7GhjBbreIzYCXy
4HSzoJGpAxlOs1wCsoprWkCJUAEq/XEfGfNMKiJ6IPiFzaKdd03Lf0LpH9NUxFyU
kMD9SPnS7jgfFldVxT5pQvOR3dc5vJC0CJWZ9LW9gQ/lqPHWN9vns884R/uZ2fZU
Q00pFdgmG5q7YXYsRQR1p4tZixDFiC1Q3TpZPPAMOxBAMPcT6sSz/VH9B3VSmZEn
fLbCtVwOobBLsmwOuJiIYVQUp2QfsCcTm3Zf4t5m4kwBnuJmYmk+ERnZiDrR1oru
Xs29DhZ8rL843sxseYyheNb0FoW1sSX5W/eIpa5vZ2FCF/tA4BuEYqofbI9P+v6t
J9Rq/vUrGlc0BHyI9QX2UMZfwl7/8oTCDgg8Fb9xPGwJ4fwg4zfI3mllC1+GHFoZ
AK2PjcIiXLzI5KjTkQWmACcZsYoci1VAC1q4JLgmyJ4T6cBW27Xipj8bZYNsncrp
9jB8FFJYIGNlFoqcQ/K+MOVzGvtOFXntpEFnGEQKHkw2fAsxtOvkTNq6XvjoEL8J
LsbDHa/3ndmI642uo6aIfhZjAskGZPQpJmDDlQpbze98F1l2sfwofoEw8c/jDcXE
KXVUkj7Bs+knz7oJVLM/71oZ7fyAE2se/IoCSs8F3SdMnc1Ss+317UyfK90hTO55
Km+yObio12NHLBwUq8OQB+moIzf8Hx99ISIG5/aKN6jHNPGYUNcMo8Evfu+ezZCC
NK7XBo0x7Ts4VZwIEhwJMwkyDykF0jc46sIsolE7hwH4ABKsy1wNppXFTgKHFb1R
7rdeZWE6xOa2Oe6oxG7fS/qaGSLCdgSySToUG6fB8cH8G0lyiw+G8QP7GK6bJbrf
IXesMEqI9uH1rnJel3fS/zCI+qXKvjvEIshsdDEJsMAXOpvaoplvaKnwlxOVI4Ym
Yi3aJo9eGv/dLiKHIaoYQIUoBsNl5Egzd0amF/lq8MMxyfq1ejXdlCg57G5Zf04i
/btBnafLuBtqalZonsMj1P/EDKuAX5jOMMPJESJXZ24L0CIkcnBXxcW4XZZi8oJW
y4C9cNpLWsharyQcCJdCkPQUNu4HdmN0mxWUZVKTL4ePejsmRBYamWVSyB2ysBnk
l/AgCeS6wv9n2NJH2ISIytpGXfrsY5QXdwIsZHWR0DSXSgJJj793droPaXHwDglj
6eE5GbVKCP8XQUWpO78V5SyWwnhHtyrG4ACcLeMRo6zOCEl59gnmTn6NlMnbxbe3
AQT6TTgC9PmDFiQmXS9wiivjD7PflES0545FhkARLbpdVM//VBADYLfPMnalGtvk
DyXE3RSfc59trk8r+1nQwWCgJ+05RoZdeYVrEX5xhkNZ16CUH6EAaxq4oy9dl2BT
OOEzyAdS5hV4EAiQgYdljZxE2DkkSfMmsdVmaIJgHvlRKJud1o1VhNJFyhCpMqUo
v64kF85I63Ym+GYSaE+ScDPl2Gdhs2qOZmlqRKQL1GFIu8iit16+FCGA/X4b5JM5
dskSsFazycYScYArl+DpqZr8iUnAMKr+7l+ZFVSrYLiTz+xoy+4uvPwkaaoNHSRZ
4E3jf80r0UVocisERvn4h667T+OKoJkViI6QSphJD1fwOhLe2o7aTMEWHJJEzm7s
hcmVp/MtbflDHnSU+cHpRogAgP5szE0CfPx7zX5dqXqQcY2sYEXC/LoS9dTcGmI7
+nnfn7Hv8J3n0HAL5CgqcRS2jdj7RWWI9c2mVU7CSg2qfOdagFoGsoJzwocfYOU5
OR6vVLv80ZpSJ5LLnAj/eUIPkRH+PVVU3aJedhc6UCcT3eRC69HfaPNJS+pDu7w9
lLX3X8dTcVr2grrZ0U6GoVSAouvuhpKxuXvzM6uF4vLQrlovZ+FTFG9GUIDpwzhK
TLvD1A5/rpI9FX2vpLIJPgZ5Ioe+o+4GDtqiPz2K0ScOBYhpKkayAedq0mwWrtIP
ovxmOjpwJLtpcUHbU61AJDGfD1cEEXt41vRBOkd52G8vbaLMAGQZjsgzInAppmjL
GiojgDkuo+1eRmF+BS2Kn7iP4Brk29jwgH8jy08vm6bPNJUuPlG/KIfYV6xHQHLp
a/fgXnJeSVVGbkrd+gp7//7YU2gY2Vt0rMrr4PKBnqJzr0hWhw5EaTSQ/+XGOIfS
gvE/0CArsLmGbArVlMBXQeiTro9w6KxM1TEIu6FTk7oVjKUqjZSQUCIYnbOdFmmy
kWc0rVH4EYOIGbWLBIDZ8D2Q9vOKf2yU7iFaIDiExcB9FdFfS06sHx0jYN3r+siI
rXA2USj+fGLmG7SD06bDq6RN5ZwfWejf1dZujz3GgFDzzWPulUpm0RxYKvT3fom8
DZG+5Z57qxfEm76LpC+7yZV5mTuttWbv40pByHKxTkEW+9sgbm/B0mmmrd62wPb8
rp0QTgOeXtnpnPGSYvssnb9bD4/JoEC5Qdeqbr0n4wTKv5cV17n2gp2pw0/FKKVY
2bnnAUSVt5vjCcIcQ4gWspd3TynkmAqjWAzTtnf4Tl62TsGFJw5l716pyA0mF2Ew
oY4ARYw7xkxKpROPK2sWUeFvwfA1F8gQWDUWJKt/825E8EgquZvPPExTG5QlTP7K
C1tcYLPIYYB3GwGSwLtToQmh+WFuUD8Ek61mxeLawh8Y708A+GIjmysl5W0knB2G
P5wDunUe9bYMu1bfeL9W/dznN9e2Z3CxOds+l68zBcTbnLHtZWbbRpUNzEvdQ1G1
ZptwDa7L3du5li49ZVluVf3ID/UUOllOITNi6DRX4BSrQF+uDFdNtF5UKTNu9wto
ia5/xe3U7Op/kXoUG3chEQFpuG2zJgyjikuGeZ/LkIk5lMalIja325V5GD/MZIHl
hpd4nvmGLzBZiprBqAtI6OFKgyt0YWYacWgffJKMmhFnhTEazkS8Bz87pb5pnRsl
Vl2ufZ927uHVUG5GbpwTwKuOvAwXrgFLbXNQmRyrmXLFLIaxRtenW5a/E7dtV7HH
sS00xg3lX/xJ2BQPcAM/0eKjtmSSJ+wn/Ei8iCNGGcWdbZPeDXXYOW+nMKRLJaGc
Q//nRwBaS7BFCN/lHB16KM1CU1eFK2Bmkmx3as+JEVme4OgSxkAhEFNFA3aX740U
vMv8cCIgzVxwxnh8wkHwj8dUx3qrIneqQyGfttt1Rq48h2lh/1LLYFjVZDF2AGzK
MTptpvGJeIV9ak8q34XkvURtr3OfejudUIo8C2lqa1xNzRCFtDzzBBYwvM5OED4g
UY0DWKH1dwvxwQtJazfBZcAUwXqNQ+UhO1xSAVZtM/EIk4jfwSSdX2h8sLK7ydXx
0h90jjcQbosCl23SiNYqKaMJf72LqjmER8aEDYcazGveb1s7qFGxEvEvV3dLe3LW
tbyvLKq8PwbMg4fU7qZwMtOuoBRGkkp64jEfv3U+C1zzQJdeCFy9mkeWoAzKK0P/
ngz5zFiAty/f8qahydzpgtmpPuAC4NO7/IRAUV0DZwnccgeEXfWAB+DCU+eXSIc6
Vr2oIiYLurkQzcrVMsZBzXnTPEMRiv6ne+Y3VxjqtCeSt0IZwza0RkqJyA/Jjbi2
sPDLnce/9JBF3A+eo6anIhGFpkNzuwaa7cOsoUm6dAoqMcn2K7KE2dMtrCVaqClu
9XT9VSLP9YeVGztgDTv5eOfNUTsvdSTY9CQnJkCDkoFcht6O4hbiscgYjEf0xJsr
Z5s7OBUWuYiwLstoilMeYMCM8WGrGCOsQaloask0pYvudOxozSFn5TOwd5SkSpp6
XSxkJjJr2iBAOUdLkDwX5Gf39jm/uH9ti3Pu2G97qDvVEEgc1sQ+chkkq6QOJEny
nLp4K6wDRAm+wjToM/b461DUM5dWv9UTgEpQQdTLZAptU4mKZQo9Akb1DjaKuFWH
69pcygUd+OZPfCY4Xiwel9frV+fqPNl2AQUFofigVeqSh1O4Uhw1TvnBk3+iMNmR
90f2mw2fUIg/fHcysQ5HQvAGheRG5Dc7bOSn02QKua826MLy01/06UAkke4ew+OZ
AKXs9Qtb1HeetzNWaj/ubxHFWTxwfXf8QtQ9DeflDDcMVyrxS+OC17pi1ghb8Rok
8imrLgaiCehBgMSyRm54Hbh/Tsm/aO6lCbRvWZtdaMDHLYeBEaQnAadgIHKmJ8CV
8FT7LtQ9O8fBF/nvYdmJkTTCuQq22bBE5l88+F/tdn0MHR5NVs0dSbMv9FvgWRHq
6OQZXA1FHzEDte5psb02DJs0UAxDeybCd6Kjr3wIyCkCwWMGnwvNn6iYf2pZF29+
aHSOyTlYl46hMhF6StE4yxQv9kqVmuZ/YUevQ9ASbZoaAKNAj7UvVhG2MytHe61H
fbnjku+6wg4Y8ktemaYrywQgva5ARf4yilQEi7Cx02c+164PmHUrUAcTvMQTCRJG
gEye7pxfC4JVBnfi9EBCPQ6KNznn5Zn9AeiBAV5owYKD3uMZI3NQ6TLlf6du3H3w
sZOivdq+61dmqLGZwN/Nj2dmfhGDsAH1ATScL3+dfMgv2kHFQfQLYcnPCchLrUrx
Tnz4xfYgiqLZBspOYSUOFpVPzOc9OrrRbzOb01CfFGMkxLX4bgJVfMiFUOJ760iO
aUMSj1HHiy6Cu9YI+Xr2r9oH2dYoBmRtV0yMxvB4LUt1oYhg0630Akevj5jd4tmp
siKSVzI51Jl8e2ZGC3sGQYNua7j6wr5iL5cfkjKc1KObm8A5fD9nZU+dxph1myPJ
iBbtmcTnQeIOfZqX4rCmMU0jYQG5QglQfSyQBMV1nfxhTipN85gtfT2YtAQUJviH
fjZzaPlroyfYaKt9QZ/DdRl60AJnXvKqNBp4xdCfmMIL9PR+Et2Qf9xx8DOCSJEq
BenyhV4rVsU2oIpf1rb6BBEIsm3Sf0GFl9e3PKxju9M8yl8irnuW0sguTYZeMAg8
jM2Bps9OC74D9w2wXG3uMXBSIRsRTpsPl2vxxGcxIsPUJhDumlGmEY9jwql18eM7
bwGZWsUYW9KYJ92OImqMEErFWrON746sPVXohEckYPCRLAHyWFartQtZdS8b9eOW
0Mq1o0jmj0iIZ/a8kL4bc3BSbgyUtrertr0bXoD5ba4R/oMduigQ5oss/r6RIgRb
mDad9aR2rBE4XILrr0Lsl9+eL1z5X+AwHF4wWc+MyL+b/g37ZQJZ9KqtX5sz7B50
PVfDsUSheOxoTt5wpYnlCnyhFctOGCAoHxl3fx9vmP/1Il0v+2dt51+rU56en2vG
DNje6tnR5qRUipiOfzFnZHYv1Flp50zeDMT7oSE5D4LLEIsgps3SfoM9YWDK51c5
t+ea1PpKGobs+gKhWiaQFIp78lhoVAbhDg+1eLcB7nnfh9Si8XochBepBp1pbq8M
83cEl1dlZtP4Xn/W0+uMbN+fjdXF81Y19guTmxXZaljCyEl1+m58gMxWUm7w2qTS
3vAeZ104gBXRz4K7reDSFZmz93pVVxgeDAQt41PrTCfBqMWh/osGgKPa4pBucROj
1j95Up+dP3Rt9N/t36OxXz6X+6VTUTM0a84waV8AKw1lrRmUgj/6/7X7R9d4Q/zt
LpMa6vyfdcWx7S8ZCHrXv7Eeb0Bad9HPY+wC7xvgyTLrJYn3Es0sSHW+ehAEOZTt
1FXFpt/BwMZzAYFcu93tkKw5dJ0jxLkNPbbrA4umXsBIcdBYDGhPXXigxtdMFneB
rKfgdynCKcTRMEPretuIz76ITJjH7yq4+Ywxxf/Z6YH5WGdH5p89UMlBw/X/Fw6q
j3Iig2KWGtEInVN9ZScap2XzmECAcdCpSftBLt8YPtB5qB/XH5jHL12irTg3IJS6
0a9u+jieEZ/1gIufN6TQwpt1wGQp3HA9QMcwNpBi9ZgiRa/Fr/SBoDYTIvOLN5D+
COkjjWiFPtF97QAb/KAIdYzvb8XAfg9UNHsTopqg9Z/UP/puIkD7RMyAhnIfCXuJ
PDqkf5Mq+BwvUeLEbe90TI8ZusItMZqghR6lJFraSLRqEsZwy8QBjrHZP5bJzCGp
QX4ENLch54ikOQumT1ts204ICdRt4t4+Weqg0Sq+ziSeXYMkf6deXguVCwYK1LwQ
FtP3HL9IZoOpDnKoZajTOQIeHVzjSzjg/V+c3PsdJfM4xxE9Q9mNPR1DeXvIOYtw
AQF9XVUqu8trWdDGd/8bs+eURBb4vwfFGc+yMWIxp8RPOJmLhlsJnO9wZjciIJxP
xnepHBTT5MZT8WYhXMTcgese1BIM/iDJ1K8rDPd0VrYRVUO3LhOyL0K+opXLjazQ
dKvWXZQ4UbYcUjVB6QY4DgW/vasW7OA+LgYV499Ha1bDz8GwTgCua2n5A745kvd1
OpL0/o40PNbNiSgmS3fi4Hl5jg2tz1GpfnHkbJIDr7HfNI6oMtB0hQX0NrAb6fIb
xVQODEkhxi4Z2G+e8wgBN02fXce0qyal8GOVKVqfgC8eR2sAzoTzCbOTAfMJrhe5
3nQ5VRe1UY54QGxSJSexoRO2SjZO6mTyNIVNRBEJgjH9vOg3zek/n8ywk+y6bLuH
haXdmczmFyZLMQoHJU1BWNfXkTztw69KISZw+1puhNhooviCWjKub0w/wKyqfb+B
Z8ND/5p7i57jvPfP7TM0EK0l81HciseoUIVDz4W5L/1wwNtRor3tSTRBAZZU1Lea
metwx1HDcl5C9mxpqz6gLS2COhFbbUBnK+ceZ7zqNZvu698Od1nE7WZJpp2gHyOZ
GpcbcdaHUN2/Y7Y9v81fyayW5jLhEcy41FlODzWQ+vl3fRhB9tuLFb/JpGKv1Url
kYzD5YR07xPSwC6oyyjchnR+iKkmndIHVQGdlP0WimQOJG+WR3MQ9d20iEde86A6
OT8cuGhZSO+zcpr/gbZPiJoDm5AyVK/Nm/pKNwtrVihzIVNzy5nZ1LMFRadGLP5l
fvs1CzEYOMBhDgh6D8JqXFHmizyJvjn87fqA9P/2oazn0e3esxvmN+LJmhSAcOxE
mFp9RD3twBeJzuvjIlNXNGmO9//7+JjtEstCucB6mcjXs37Y44sNjMq43INyQRRM
XAt48+NkdDdNsU2SCFr8s6hmmOL7Qt5H0pZeit/gIg4q5k4vgnBXESlVm0BfCq/R
M3x7pf+xZtaBdjtKwixErI3zH2W72wSYbPVq6V9/eCPmtRjbUZP4TrlfQQX7LKLr
Daa8ge7OnsaPQcumI5ZOY43C2vEo4V9HilEP3MGsEdJNuofe5bKaHW83LeczlOCX
NYsSqo5UW9bKU25hkJ2+g12PBRCGrXhvvGM2Ph+uf8w16Mkyk9wbqECBx9bdLcfM
pHV5mngaRGgBWwXbrczNssl1CYLGZHca10Gj+3HY6lZcbfUbqgwSwxwnYLQjmJwm
52rP8rhPeuq0IUM5n5SoUQo/CAEMLOL29SPmgEol6vorOdge/oPEYnBdF2DHX3hC
49zDqHlW6P6XZwAYUm62WhPPr44fn2YY6+faQfpI2IHoWV3edbmPU/h5krtJRycU
XqdNOJ1KwBUAKXoiFPs1KgjUPYx0u/if1rN9+5BviAOaitlKjD3FbIuz6Av5h3CG
7BaTxtWrFjo/HWNkU64JxNyCQGFVp1552CAWb+Q+P2ywv0ddDQOQs3FgGOMcJq0B
iNCngYhgSsV0/Oersk5sTELYOCeUg3WAc1/wr2CCJfU2l9gmvizfeIxrGdEIYL++
nT4NRZ+ZWgX2OKl4+MVunIKl/kka6a/7J+OGiJrlwcF0FX5e3vmDnkXR7hZcMKxz
VeZWGQqjd1x3RHZsOAco/09P9CPBiTzRu8Q/F6zoNWzTKJR2sVw72W01wN6827bE
KdKZRF8OaW9LgBHDPWr+duRzqOAjm4F2NXhuARTpwfEH3vgeewaVX4QkuNZZnGMt
KrKtBgZi/CeVH8QUBPagiV4lAFceXuS9YO2qLBoEsOdQ554qk7rRmYlAefeJFCqf
+0v4sTm4bIooJG/BHjVGwSQtiFOiChskmcMjPU5mfTAskT0qJlQcM2eRs20W1c23
YVpw1tXig20KQiQWGCwiL+zW2kRws36SKvY1M0oLIf7Cy9ZGmuaFdYdHn5Y6Wgdx
LAfPnQunyE5N3XiEwQHtas5zEudmTPDAtQJQfBoVunnSeNl19X06Uj4LKDzB3R2d
ePAcvwqZauvoac85Q7zPFPxeEtFhPzjTltYiYNLcRbtGSDJLLRUzh1lav41eLXuv
F1OUrHjF0BZ4lZyBWwvQ3hPw2PhVhAng71aah2GXU1WnEZMkxsX1qdw7c4LIrjYY
qu3jxW1Hii4XDia2Ai2RcPR8jIy2YtYDJDtBAdYNW1umK75ZsdFkfbwBgKN5pkae
sFYfDCPbC9HGb0bpjfIRmytAjAoe9w/opBErWfnyUNZOHnnaDsPCLPDEkz1liiVE
cUGk36ae5ZFFPzTLCPokfgUFavOvKrPdyH+8XBFJXZaGftmBPYUYUxnf0waXM6Ox
Li3Nk/ph/0I3vnYhR/MnmRrpA4OikZVCMjAxHdgtgD1rJLfFRDErHP3M9z5X8Tm/
zCeI4+z6HXj+fuAQSTh+/yc9tDv7vwVHX1mW8DI4uHJpluIU8idUUg264aBzj8u9
zKCxZod22skGLBDauqcgOcukJKGwkR26i5gh4XjPCSxAs0CNgsszcd5PQqNC/j1l
NLxXtaTBGYVJGDHFdZ8cdXfr4uQ7zy43bqphTPAqRzsN5MCtd5gu3hhgwDQ+07j1
k2smCwN5YKZ+5+bX2Q+3olGCgJ1Qqbq6UU9Kems2Xv15jokag4gydCXA++kM6H7l
WcrNPuBgOtqiHoEq0ARx/6xUdUrPLiCVLbv5kRMC8m/rIP/WIXLh5oRpiJWbuN7A
gfDHsqo0vMEAlXVW+Y4HqylcAYH83Kib5pfYzKgRtc8/KQesi6cnPtp2JM2lJe4e
oxzRt5qztgL8YZFXQdvfhtqA8zU+1wjzjNJc3tsio0YYO6Le0NQ4pVKvHTaSH/7d
CsWEX/zo8ti6wRVXN7KYY2oEiCy1XdvQ5jhPUSn/fvYo6F99BUB+XsZjna5Ghqhn
VUNLN0gJTD6i1qLEEAJs4pDVLjC6lYgwWrEglMrdNBvu6MkgXDsWVsy6rQpznrdc
5+ifsZMHNUGLG0OgpuyH/drS0UPKSlgM+A6PNOdwTJR5o5uUIChTs7p/7pbsXo6D
XaZZFCu9iSBueR0Q7VYz2ZnKIocuY9NrtHXX+JYI2ttWglFmcLjNV8QzYX1ZA1tD
dSqiKZpr/oHYFd3g6Ktv3qArA0zBlLnHs9PXnus6VJBP8iNw6SqcLdIJWtllchf2
nXz0AS5YSwhmcqUOVJCrkmSyRHAykdSuvlR7GZbPOEzd8qoA+hl00yFX61sKnYTc
B+Imq9mT8r3ZKMi8b8ZMPOHujS0WxIq1Ck3YBS0x21HFb5quhU8MfZ+X1EWKKINi
17g10kh0b2RDlQB9XamNqKXl8EXb42+l70ytNsH/9FtQlId68OV52oRk3YAhCScX
xEB4+uHg/lib+L0JxOAfanDNEMfA9KQk/VpJRxxAFdrpqQh7MpcvIwPJS0pI32UZ
R4WYiiepRSv46k6OI1XcXyZNc6p43nIDrVFWOL+mDL9Z0DmkCHCHsNdp8sL8C9zr
sodQKxEJMRY2cqpWPdKIYroiaM1aAejhXC3r9qzjB9GhZyX72W/zAv38eGtuOWLP
JDIa3Y6jtqsVUEq5yGSkXBCdpj4fWWThtyu9ecwQaN1Ro5YFEItcpK9526R3Ehzr
acKpkzcKt3qica+ACiHkhzuX0jRLiNkPRBkIe6mIovQb62oHUz+364W5dugrr+fM
I3PGsKmHjWM+c1DumWmZoHNz3qEUs1vafepAouAa3ya0Kq579eQbnNwpLGpm1nEE
Mqm4KcVunSqutTvz0VOBgkVa5i8q3o3z47EQhva507MugB7F3EH2Wc8yXdL0ClrV
uHbuo6/8sDT3Hylbvy8SgGyIN1UgZud7DuWTvpQDD+5P9hWsTO/O9JdKGM1MJ2X3
t6sIwuafhGjQTVMKGLmJ1cx4FGmQ5k9wZ/sBiINEpFZOHKC6ihmQHf1nWOdAifV8
8JW4VoYEWxB+eyYYLVWyVqcVq4W7qx7rEsdWC49c2I3Is+SGRfqUFiH6ZgDx71Bt
qYbs3UfNM19yXyi75qv1kncD7ATmF5BaDfaholeTBDK2LgSuKMRUJBWGJeXX5JIZ
TmUOeifNqOua5e93F6jusfo31ZS9cfWO6HPtZaItgDK9bpV0GVRsYNTfKIOUhr2+
eS/OrETPm+CadWSieHK3mYRQ6kIPpELtONlSFrmeJHy7JUGQwsvY8KVr40U9n6HQ
MhPoyS54wNaeJkxIxvqmWGnL/G9lN5Fi4OrgMrsldc3qGqULtLS4440uUc92p6m/
ynMr8PkB1925P6oYfVCltsIkz7VNmZh8qIT6gBd1IaFDn/+plrUyARTsi3g+FncP
03P7lFmfonTyx1+DJAvBrYeO2cL2EUSXNwN9WcTaDbUl9n5Gj+7lLUHstvpofaQu
uC1yIa/xWcK8LhTn4qKOQAVVvkCaJUi/xNkLdseb/OuQcy2CWPHPypLJP9AqpGrF
+MxuxfTWxjCZUogCYq30IRS22YZQlP6Fb1x94dMcTbELk9q3tzu14rpjD3Wr1cXV
zgTiXA8/CiJkU3UkDAeCrH+b8tsvlVh9SFqQe41RVxJ2QdxYD79m4HQdAOTcZd+B
/PVkyDZC2AK7ZAGuI6SlDveYnlcRKbJe2IBsEtm9vrBil8Dm+jNb8+YAMRb+Uf6d
cLYdAQLHwpqU+ijuhTubUfAGfEcDWrLJ2Lg1IKWYdCQpNhNiihVbzbjozjwztTZh
K02sxnBbCPw/3uHY9Kiedp/U7fYqiwEvum/sfGmKov8KAhnsuR8NpSdVmDMuUl59
Q7QWcE9DcF8Ukrnk+Uh6EtZSrICebU4RQ2pWvZ8AkT7reomOp9x+6vaLRSI1j/lo
UrwrsP+uvDh6QGMjmtCJ7EIjbikwTaKCctfo0w/bt3lXzS9tVAKbgNIJYB0bYDAZ
WhP+3FOSxy++NImT10xk3woAPcP+1kqJ0+TOd0dr8V7NNVBDEZ3bBfm6kzlcc4fe
lxPoSRSKHrdzyFBRKJrLkluC8zdXeB9xTX76Kqa17KjNp1Eya9YTH7FJD2mkGIQz
sSNmz6M9BKIWFbN2Z8dEZEhhKEZ7omC8Ftj1uOT+MGB90mx2Def10hJAgYO/tWzi
v4qD2bMPtSxnYFNlpUZn/qjmjFdTmNnMJGaJYdU4pnT716Yh2X5oLq4rcGOyIwwL
cMY1XXGbQNaZaaTbq6yo5zvpLRgfjk7BQGtqHWANtE5U3lcDZ38MlZ5GmlXU7k4+
pQ/QhaVVOfBlze9bObFg9ezQF8lFaUxvvtIDM03PLExBtKfcEwUxdsaXnrBCmOfC
wZZfKDeAeUsRzxJOwuWimPG0dmWTuc7PyoWaAJOwftPh5ZxcZn3jt5CXJozb6qV0
TgSWN7pOV/feGASdhgFo5oVOaetoLcIyxtxbKo+NLQut0k8XbBGbKi2U9i4yWRBz
8qIPcJse2GmhxXz+Yv0pxEH+iZcvcjZxquCvHOr53UrvQJbTMLWNZ/vZ/FOLEj3J
i70qWsBx9tCxHIlvee7pq9/w/+IQRpPA2F5rifPcAA5+XyA6Zrz3KRs+gRQF33ej
1g04C7nY9+4+vZya2M2BaTIiNi20peeTNHn/HzTg1/EXg4gA3my9rOQt7grjvUNJ
8ZFRZClsLvmrm0i6Uk+kNY/jjHL3bG2mxzIDdYBJOqUXkZJxngpYT+m0H3f4ZXby
QLXy6iomO17gMffItECIj2+VgI85PxSQD4X1CmlGm1wZOFacJreFZtYxw0MWeXiT
ZER1Yjr+1/d0+5BS7TSJLM+SbWNPHPBJRjaglk6b3d6DBpFlFR7lRHYyuHrH0XyY
S2YsV7hC3ZtOBYeBP8P3AyHsAYMfuc3M86mUEQByDv3QuWP2PeBxAGfQdyeHPkxb
4xOvX0kt5/Ud5Uhe+Z8k/NZxwO/75xPpro3JnebKZ5keS7Otf2X5YZ1CoMdvoo0b
nDx2zH6qkVPw+IwMybuFHHrOSIiH2GDPJnDhSyHAm7EQE4c9CXcAw1GEoGhODkWJ
uWKA1wNZ7pU7kw/BUl/MBq89gERsmVtAyP05Y7AFOxaLk3maB+lIcytnxrR66BGd
fYkKugIUZluhDJGTsaSiFzz97ryAQQEJYR6ZA/UO2UVjeLoT4nvxeA/t831uw6y7
HkwW5e0ibNiVo6hL+DAu9YojpqNnvC/bsUNeuICETs5RlAeGLaxrUH+Wk3TNnxz8
JFMh+qKCB05OpQsdcmjNOSPDR7NJB4lYYHAPWJYy9EgFOTyqHvBUjBQeQTwJXfXo
8udRHTiq4yhBfinyHrwcLzo/Bccro/ONVaReUKEeBvhNRNnN96+7m22+rX9v2bka
sGeN94jwPzzIB8r2vrl8ljo8ezsEz8MMzaIdssXt/z+7B5l7qPPhXjAE6nlCr9kD
i1YNyXZu9qN7EUVPkE6HlAY9fIk+d9Tsm6u+NOn4kOvy4Kh3MQNiQBYM6gSSyR3t
H6i6u4BIHf3HV+f2PKO6yClzUWLjq68B4jf7PM9W9sHexU6kqKh7YZFEDUFeR3Rk
5bSW7XmLfb3k0VQQDWKyPWROTai72YU6FC+hQmMW4v5r7Yqb3TcXPRVoeQl0q9F9
2t2MYLzT9vjtclRwmT0s3qii/OUAhTeFhP3asi9LtukqitJAY2y9ZYzlrieBv8fR
ZYf3FVLkT+RT1h7hCk/9rkPzwvXXOO9ApO9vk80I3PFOhVgcV7B53Y6JzkgG3rWN
im+mrtRWyu06P+KhyRL6vHO/Fbu8GuFZTUGRgbWTKXgSlyPv+AQfebPnIo3k74VN
p7Kc0coJSBuHcMKi71JUxok6T8giKHfjV3HpRS1ByhM9tCN3ZjpTEHYbjnkkW3ai
nDk/yKYBv4i3d2ofv9rFo3yTCG4wdk9FsXFJF4m1ftM2xUz+L/dxrW7lvFwEPjP5
tDG5t73aC/2hUo+QWg5qJkYsmSKHInqN9wMeU3WqlKwV1zH8ib6f2Fr9iA1rHSp6
2qsRQCr5AetVQYkNf7e7hperW1MvseoQeG/oIrDByI3QmkmXNBWxK/A8Qz1K5BoW
BUiCGMC1raV8EpanhIrKPMPrdTOCJU9nn5xQD/JlSohMtev9JYwwTI8LP/Opk+er
Bc9WqMHgf8YvO1fr5XKbMQSxgBp+AQVx2fPGRzo5lXc2cY5I7TDouuW1zoMk7lSQ
6/W4unbiRoq9E9DnvKM9lLF7KaCXiKfyVJd/VCYN/iMsxFr0LjhppjyD0oopDWi5
BEwk3DI9ROZXGMuKAZ9uMNPs0weSYMfJncMZ/lECvRc+3MNuLaQBPxxFBDxy7nL9
9KGSzbIZ1xj1ggv82LYUSKHfql5YFhzWPhMB6V/SCJenTwt+kyLNXNpfEypV5OYH
zZ1mz11zIe1LZSrzf3bNbQeplsPS+CsYEziOTGTPyojt9SURAYbmG/7j6gPm5w4Y
QZh1So7hEASxZwoYmfzhMJs9BlXw5/1tyZWEPEmr+oXVfv1+t5BGQEZYovSgHGpS
XS5OoF7cayPv9IUZLdiBWVcf6/HTccA9LM013g3RqzYFWdUfoA75idWFe8jjGs7K
vE/70vTrOxw8qAcEUAdFCTTDoPR9ShHn8VvVoMBEJ+Amq4b+km0Ojs33olNZwWNK
QBn/tJ8gdphhHHWip1YsFZtyZtYRYualBVLHLSHyuDnlH7VG4RBOKaGrtrXiV6FJ
28X8b8C+ljpwwL+RH1qwE+C4VYEBOyXUtnQF4GabpH9xmEWcdVK8uDo/hV03maQm
RHLcnawGjRGBGj3HzrcGz4XmtCmtwu9dnGP5qHVV8BwkoHm2nHqbz39e+agq2A86
aQ/jbHJw7MHc3JPS6TXKtuk75S6NH0K3D6rhL2CQk+jZWyMQuccxwWegtSyrL7z6
S3Rf+0SGZeEnCvKOG2BsefeT8xJqeiu1j67L+dWVBP76ZKWV1+Pp7BJ+OMEKDLi5
SI6GfPgbwFgO8Wzzyla5H8L9W8klXUAS9pG78xbl4/6OqcoPk9pKDnaT7mWwfjUA
Xff8uphDwmE4DlbWXU0h//kmDagyg82ux6E1BH5u61Qit/ysVyeGx6CruMonLjeL
H411QKxVSzgkP8jbBZZoqm9wj5Z6YvZZQ1ylarGuRWG1Jj7fKkl/2U/lIRox1xNr
mALy6cKrSVG48lqlxn4WNLbcqu4xDJ9sIXG8AfT23baMsWWM9nHzKGdMhFQ802MB
6TOxh/0LBDsaOjJX6UeaZMG/p2D8x9gsPZFhedOtzEpU5UbOUA/6MTxJDXi1dm+O
CoeT86biFDova6sU61B5Sl1nYEi0aV3Uq7YRfDI5Koy8KwNB4EwzOhLi5+yG26kh
2zHw9ZZrQkg9DrBrWUCT+jTsKSEY5R4XaGjUpBrft7gAy2OGRpFR2QF41YtwuN/n
51gwpaQXVFdxDJVvi9ypAMLgqPvHi77ECpMzc0iqJcmBT2fyF1kXBV4iSBL+yvrR
CRXTnxNXiAg5BnkinFMmrUNk4gE7kfKMGzC0uAx18O7lpZNX1crxRHxIXdXLFS7E
s+fFHxUN8TETL/fouez0Bg86ItrpDaJKXVPRYb/9K3IB20rnCRMS0932TjkNw4uv
Bl5wl6SSeyDRV78gbsA+4mCDshb1KX1VFjEprDFAVeFrXQa15utQr2Y15nkvv/4Q
mTypWjg5mfh/Z2DMAwnSpiXPUJK7AIsjPdxOH2Nex53vwYoIIHh28MiHSBN3MhRd
jb8xu70OSYPMvv6Gn+WykzGhlptgmkaotHFiRUbuOsts0N9evG3mPkgjQYxGZ8EE
BAzYFyHTKye1UeI1LxAdUFW3WKOteof3IRDK3IGLAYWdqWKPVFTUJXxx03CvG+9T
HQTz/ANC5z8qfhx8Yjo6WFnqXAniglxx6oUvMrqmDWU43uwHHwLL979T91P0+0De
g64SuVlyTcR60Y5nwK4+TuC8oivaJAznlXqtYizH/o9VQIpxQD9P/rZHnLEUW2CO
Gpgsj9/RchzOlJvD2hQat0KGPgFBHwe//io9F08w9f3UvWgrdT7/+xSJirOsmG3U
CLKyq6oDgF6ZXZ3Tx/hncdJ2JatwvPQO2tcQ+c+HzVPfPQAXUC62ZVp9TTOGahrM
Krwljj/sM41iAtitFt57BCNcx1V/XS7XBdjYSKxXYm0mN0B7enqeTSvtR0scoDg/
tDyWjpIHfVBdOX/L4INvqPyjQu80i4as4UjJfrRrKvc6GHPZNLYTQz+zgdgWFUul
+1gXZ0wFNvhKzYLEr1q4/oHId3xT7vZvASwj1au8e4nYddxOqEJy6ZF+kzFonsLR
YVPUJvuZTPuMl6Eg7CH1+DJ+mK0aHgJQsqrE155gTV1DNeN25mvyYsjYBeBDuD9b
MDdWQgIyUVNaIV6KonOuc7EujKVuJLxZ983u3W/oWCNYv5hnqnV9+DGhSmEhxsGU
WIE4UysVfdxtfDbF1kyQ27Qfoqqwf4Q1bLbWIkTvz7+JkORv4S+EyGZts2/z692L
DclwZ0QaObOkxlRFuVF8dXBeKbgpOs++XNUc3pfExnF/JZEXbkJqa3R9nm4gZFzE
EmSZaDwpdnoryppEHe8MoI8gm+PeY7UPb8dgTBPCQ7MPHwSfkhxGap/0YYNRAXXS
YinXzH9gFczRwXDhNsWmT5A2kd6cmopqL7LpwWMZudvO4eGrqubwk8g6fF7WjQwQ
2F+bYnsde+MvTRCve9WBn8bwsO1kkyOBKqv2kP8vj6hsRcigkDk005oBI6CGS6ka
9EnQlJ/Gogi9BOD5yF2BZyxM5KS3RRjdJGD1oQu7MdBdJJEqrTb9BkMTacIyBlSB
Zijtb+hNSXa+FPCKZwZuzaOxYFW9Kf3qhuoom5bCpGty05zl4GUJwdSUXRKEPpKt
hO5BnIkJmc9oVxnt6W/sdX9SG7nCMEibesDWKrIJbiCCztbEspbDj48OJ9T/8NMA
Ma5buznf5XSe8lYn28c4H/LRZ7jBSdqIwcZzhLT5S1S6BJRsxJQRGqtbbEJN/iZa
qdepdTkIyl/RepcWrdaQ7D8z5NoNFhlPSH4zzCYYhjKjQgTF5dveV85O/Vwx91WI
6NP9ZfuSsSb3qec06efagngj1EAEsilnvExa+XyLSEGMVkvjGDwnpjS9EjC/ejeT
d4megE4k4OqGh1ibtbcEWVeXZTuNrLLd7DXIlqm7lBz1cVek0/TzgSjYeegGxTYW
SrNiBdVCTtVGrpssTaNH/Ooz0JidXSkd+QFqAN8roifUFA0AoqD9kTTlrqBh7ayv
3Wf/ZIILQ1OcfA3T+YX4gaTgmiUKCvv/JW5O2RFQcWCmBuDHB9UuRzMnuqxgv95k
Hqie5C4xjAA/xfpw+cMmqOejMF4ZU6j9ENOvk3gkyraH8i0Ei+50wG82pKmnPCWl
DKfwpopJI2uF1p4HK/6eW5prumga8R3LkqdxtceF+yBhmvdDtSByFaVBKCNTT9QH
bu2c9O2Zexik6UBFO8EBf/5sypQQyZijc3IWS9H64tC+mO7F3gBLeS/RGkZ5yDtM
Oy3uAEFFr2+tjAtsi+CiK7oqIo56ZMnxCg6YVD+LB9l/k5uGIE5KbQjpiirbXq4a
GGCorRBq4I6J63wv/+O7eD5FEeOEkhUgDvIJd3O8WjDOk68LWZgY0zFR0T+Cj/9T
ubpGhWWJMvirnmep/FG7ouq1FWpi1sNI8wWHHz6aiUS8QaG3XgYXo4xnXmZtyTF7
4OyUWc8vsEyPklncw6FkAnnWybBPJvyIKmAXIBwTLibyFQQ+yJwfCqYk3F/BmolI
Nhu57ydY182OLyMvppBzyV79WUOeUJNozhzihP5rsNaNWwlLgTALm1uq6b2GqxTO
ag3BA9nkjNILr+fKIHyl6ZP14cfeZYgbhmrdxDhAVqf7UZ2I19o17dex1RuaHin2
uX4agmx3JQ4CjZORL2tzxdu0iVP9CJBBxXdfZw/ArSMoRUCt6jXbLRpy/40urROO
mIbUtbR7TbH+odfAzoA75P3j4mW8+5iBlXNJ57eyfuU9HxZfxpvbd2852wOATXe0
XAGNb6EvBu6uoRurAfzjDyOvyBvHubGtmoIp6GZPcnKLRhE5mN1+PZQu0F3bDIRG
l4HSD66c9weisHBXXx6OSQ0iwy6OHxSjda9J3eq4vtvqCruJGQ6vXiwtBz+U2lyf
IfqFzjm6PHhXWS5riCf2YwxtYHxx+/arefQ/IItuEiWuGefryqjIWuYpL134qz3B
xwN9NXVjaBmFGupIbapFAiYMWrE3ZRy79I4tSvMI4vVCGqN7B+XwM59+99e68O9K
bN1pV7T3lgJGBab09ryHulE1IqlOP4Qb6iliI7iB2SuHy3h8ILm0Fe4BWCu56OYX
dGaCjjmi7Z3Qy3y2S8oLlEbZ6dNrEdzvZIm6U9620xb1V9OHDWGT2ZaiD6YEItfh
V7J0H38YWlaZ7G0J6XxtdTM4PKdDKMiW6QgtFasJVpqC9fBHGBdjZIZjcvOiTFjs
ixSgpYoaljaROAd4QGRgdiyRCqHQXG9qwH7yct63VPe3LKft4Giq28XTHL1tdot1
TCVqTMsG+31aJosWu+rCFTSRPUN1TGG89K5dCgGpBc6UQAbHF3HSjkQ0Et+BXXh5
T9Kjpuy0En3oY0Y0tj7PtFza/M1T2GrIU5lH9uX4xD0H30883pEwOWGaD9mHE0jv
Q/p1OWm7zxrEel7rwtA4yAYC2sR/48+veSAIPVNGuIStObQVEqPx9TAaYhd7O5Of
N+er42UE5rEYdYrECaPJKj0IGoUyBLeKmpLotP+Iu+x4FTq7nX4SOrvleKsRd5c4
1LsOalmvey+j8M2F5dAb2Q5r51BFp4inelDe6fW7K6wBpbJRbRNEn4hBBVxdqnWl
HEg26Kyot2R2/CQfq1fgNeuM5u0LWsppF42W9pDbPkpma17BvEvYf2qJ721jvpyL
7apuOz8+5lQCivVWHL0W/bOuvFVFJX1u2jue6r+JmCKsH/PWJglZd+y5MRRyO9ED
I2YQT4xP9f5FGtcaK7I6ZiTP3t8l++7HoaTraZds2XZFbCWYgdUxobPGiozfjK1Z
Sssg0Iml1MmZrUjL32MLdlH+RXqq4tZRLhKrM7FL64Lbp2Kptmj3H78LDY0/FeGY
lHWlFWP+Bm9Ap4zs761H8sBxENxXK4+quC0+y2NltfGGxYagjLdwRdGqkeX2Mb2r
tmMYCOdYizaDdYeCgF7oUm8OU6ulZJAcuX7ykj+wca1OTUdNdQqZPY8i5OrdlUOo
zXs5cB6hTtojWEreU2e3zyGQfvGJmEGC+frbAjSD2ZVNJGAl5FTEhn4nZY7VA3kp
y1CFNvMKdKFEc9DC2xn5INbaZMoT9E/D0sA+CwCLg0vIKXaU6ZkIwtiBq1U/i5RF
dfs4O4WQhqPiP79yn+jdY0XZm4Glooo7uewlGsHxP3wa7pVjb7vpf1GFufEtzovh
eVnzXWNj9uipSxnAoxh72BYlDLVtulQRArbZkEx1xRo2ZUbu2LTYgKtbfLn33skd
rNHfYc2wN1/WlxYP3HGZAl86max5xmS722nCjlKxqwqzHkXOc4YINH1y1ShaAXrK
/2GL8CSvYb/8g22Stp3Nam4SPk+le6uGq735D8ENarUIp3pMhCJv4Pz+bY707gPV
gG2iFrUHlcl3bY0lwjM2M9i79ZiwaH8ulsNSpRQlr/ZbU8j6Kw3Ov/NMkPjZ1+fZ
gP6fxdQBOobTEgBssDmGfEat97zLxWTtl05avSx26Cf+9ZZRBEijyN7klKFwLdoc
kA8T7vgMfH4QbZ9cav1RZ1bvArf1rVzrwEXDzSALviFPAmCOyoUNEJb9QAtTFJaq
tRM6h4PnJ+icmPgYllsjW1obXct8sgZyKckHI1D3E2o2XaA7y6zl3EvLSjM14GjU
tXTRu3clWmlS4cgC0qLH+fjH2dK/LI54QV7BHxnTRake0+vPUnl2aO0dGt+sl3wK
5UfRlBbvSGj8+IXF21QW7+UIIbu9i/3br301XsqOSCSsN41jUcNT2Y4m3Iq6ukuK
JD9AYia8Gn9LtKfc6gLBjo4fqsVdecwd10mD89MrJqvO32VKx1syzmEopYMaQqzn
tXIOvHzHTSJHpsFDCOW7+aaK1klrgtyiaOYT2xRK6rS6KwGwAedzUS3hCbvYpkEo
x1xaFqLgcEF+EUTOcAm6nIdJAA4tF+Mfd0Gfx/BU4tx5ZRlT1Ums1FcuaxI53ha/
WXPhPz49XSsUNpIb1k91bKvf08jTkBAo4Qo0/RoWU3j8Ervkb7W6nZAIqESFKg8V
Je44yPZBb6qeEMd+JAglAz3exxW/k1tWAj0QdsrIEbuOsJ5JaA5hZ+JpNorfbm0o
d6d5u2uky2/URgrGechQ3Nt6N5Rv8KPnxLoObXCbRpAkAlzqTaxe2SG2jF1OIyRV
OiUwxMHKvKh5Ob/60jQwh2KRtipYkKGW1aQtONGBI9xtmI1H+c+ZBodkYQ3b4y8H
30m1nyVDWeBRF3TVVELOv8Le4D/sEmjuYwQldck6up3CrwDZX71j9i7dVpvJl/Db
/GpIXYADq7+sviK3uQ7XKNxLl6bjjvgO5wuvkGo8XRdhsMRVxy2xf9Qy2LVMBHah
To3CiaPkRvcgmHGoqZOqvElKTvH/dVAss2oN6ctpF8FQKJddOuDBVqaaPQOjmqSe
MI1cnNcuYqXLAI/P7Nunaohln/jHVnR9gRM91CSwgb1gjezoEtaw9IVbiiH8SC0/
vGgiM3MY+nsrr+AUyg5o2bFtDLwC1cw1tP36xYz8vS1ToYMgS5HGjUHE7BLv/IK8
grWKQIdIV63APNneRGDWv5YaIun2r68nHoXUTc9Jgtk3xQbZ/5o70H5K8fr1+wFE
CA/RDKIwceTKBNPhZuMzVnsgG6NA1z42o1HklDbMNg1uTwuMTRysvaA1fUOq4n5U
apb+DogLKsSmKAF0RVSq9PPC6hm6K9pJg0G2LliOMsxUHF+Qpo9qddaxFY37w4mg
7Dj7PerII+auP4OdFaKYyBlgj/EASLYYBZPjFncIf9B0KdJuFYiViyv5WoWBGx/b
TlDxhIovm+VE4dkYYTwoKJcvZG7cGCgb6N12fpiH0ZWHFSk4Ta0qLeDHE3j6Kxiq
l0Ii4x2IrXQD1C7J3EdZNhUrMbJoFbNrpBcdnqTx+2UENt9kqAvXNdYrXNDvH7qD
i8qLFA99br9uWxbmOOhB6khkfxoV3yzmjAU+xH2GgA0V8eb1yOny9rlWQr3PvaDo
VrzhS+G+oR+lEPE0nvMuqY96SDnec+Kg0lPE5c9qKU/PtipP1xoT5nniPAJTAKX4
zivRSviNykv8zWUaM94ng/JbA2a5t46CJB7WljUNtFldKJvIBLuZCAzXNF9joyRw
dHFsaVf3YK4CgGzgkNdHTyvWfR8wIUXLWv0njx3xF5On24OWZuN9c1HTjuK0DeB3
j6Ns4H1Mkl7uLkQ14M3VbJGHhlneCEHnPKBa/oIHHv0RsTHk3MYJy8dP0u/RF6Ps
BvDrMMwbaJLhMHWEXbQjVi19cXW9r08uErRzlUlG8lTH/Ah64BtOfdsKp3xitUDH
PZ53YJmPytaHcuY1CCvPd+YOnAhAp02BTzrbw71GC4opQffEgLbFlcrV4YQ9asJn
+qFxe44N4b2vzGAgME27vdepLhauBk7hgyY3dxysoqTRpI9HODMVFNp4ScfWmixb
mAP4LHMac67M9zzs23ljap/U4Kg7haaVihHdBbCN/j+QFoEyIFh/MctPKyz9Uj92
IAJcHkL1TpjPEZEd5g5c6m6LiFpbetbv5QeKuW08Eyqj0/v0tUuuKFq4XtTKJYt8
FVBnRYC/bULGwvF/dJnIG5EtdG2hZF+dF0k5unxjDSs4xmBpDLLaIUx/oKjJ6MUb
Nv8R4LW9/9A0LdpzQGq/04E0AzfI3BroSj04B56e0eRh9esja4b6TubEUOS7elq+
UIxHt4ZZxw/89NXDVRYV8a7Br+0m8jIm/+YDIjTztLXiswmA0RKiTBLKpVBIkuK5
d1vVDz5y/+lN19WnaY7YX6K98LXHh68Kt1PqGlQVzWVztirmvcGlryx0mSYcPsVf
CtpJesoF1n/Uq0yApF38b3PtAxwAvrMNW4h8+zYUfwOtZKn6lbrZ9bdS1h+pnEc0
zIOiSfqXpJgcuxkU/ExM38MqDaPUfcrLVYnoxVqLk2RxRxwzruiYGctUUxRn4ZWu
vqsAsNupxkIPr59cB4qDpA/ExDncCXo3vV5sbC5gCVRpxyR6xI6gNnho6dZGbgEK
2EhPWlqm6fliFBql1jkUVbzB1vKspPcKnqy94T7lwq4mRtbjUnZP76PSo2FBxKyT
1US2UihBznUlTO/lTxZ0cB2Vu/FhcPUwCQCRcvfw80tZFhfpBeMB7Jk+50LaambH
+tFCgRCfwhah6RW5DIrj5zjP/KcZlPoiyHiYTVz6Qfsq9kB4l9kVon4eSh/TySrx
IUfdg8CNDW/c2Hp7KmEu+ppxKV3o3LpnAeRvgKt7hXTPLoueMufzezZmxexLJ9b/
nu37rVA0d6XUgE4g3IwTWeKwBz3BC79zqqkm9c5hjBaj2r24Uh5K4zxTqb2Di1sl
tT4gV9bCoxKoyeXdZa3riDpMvON7L6TPAsdpPOefaD+XMrhhxQyz0wx9KdS0iyQ4
ej3pA7FGDxlPHm6nMdiICtO4cVZt1qMgETiL86xXJxAJJe0YWrNo+QCnCQzODyoc
HXxdNAcE+Gflvh4xtnnlA1oJy9dDXdh+ME13wzskYU39iw+GQ3t1BDSEMgSSgcVS
bJA3QpjIEJ5EY4+7OkRYcJSYgZlCpkyldYDELUxCNFyTdVBnXFxPbQaeh9oIKsYE
rUhJyYZeYNdkSwEr56Sd3ZqkGsz8VQcxH+Jwc2/PRLAjiby8oqJlP/dmUvBHIUFX
fSa2jkU+7hRu3MrwTptMqr33Ta3hxk+KxPdIbUHFuZPoVpzCJaxSsvDtdgQVy2Ga
cqo8jbvA33sKqqlQnR+9hFXqO+Qs+gwLs7dWvJfzQd+2H4FOxcwEkrilH6KvF3Ol
B6y9rZv3SvE+XBKfrI5jPD1Vrj6wPTOQ6UdPj0zUE7c497QtuApyjkUhBuecBPTW
XUMPn+/V5YkUt1Yj8aQlLlwLR3mma74MxvOQd1d1FQc+RyplS9UG04evasb/66mP
ZXeyJBZj53jDnrwr9kPgUn2KvnkaGMwpbPZtI0b0TtSu5wkSZJ9jXAaXb6LGCSJO
NUgYKRiCMfYpqIxGSb1n+l6oteuY3ZLK7YS2Xd6FOhVud9PeiNjf59HYGXieF89N
mcNNtVJjtUFTGGfF5WmpHHJW/bKrx8qV2fYVetTPI7x0vjQCtFnA3gtpgJEI0RyY
Bd1wSpX+SNstEhbJ29hbCsmU6uf0fJpW5C6HPKrWQl1O3IODb72W++7jzyj3B6JX
F38dmgtEKyE5jcfPQIjV2j1pVpoTZsC9dfY2jZR29gE++Odx0SAQVnWXrW05Yvqo
SDT/fai0iB0EaumeHtu9tLcZgFfmOKadTO6Vi21+Ql0ypgYXiGZlRZpycNgxRkd1
DQmknPU6wFx15/3CnDvI+bNtdNjlmNR+TkBLUdkuJOdxSjb3gaJTvpNpOfWW91WN
0BBG3coJxIRwEpxdZV++/o++AUlgoMB6co13EhWReAoQDOTZ/quwRvXAAS8bCAUs
AQvaBGqhbR+3oWITlIJ6ITOePEQaalKhA231frSMsB2kaBaRLOK9JCDc56riiivZ
8kYC+dWsVOpIkeJVx9UVmjrTB3lhCEtHEfkhkl1EyHFcL2ahIaC3OAeglqVdHM0z
rsK7qflaHF6h0bDCVuLAHGMy2rPn5hx9qb5xcx8lhynMAGLW0QQkflaNnf5K9YGr
Aawk8T5bVk/TQaMstCmW11ddJ46RKbq75RTXE0tKgVhMEA14QTXIxXMIKFehNZcx
ugbYP2uLU4aTCym/LEs5PTVTIhVI7Oy//u1y/A5zuZVA3Jo+q6G8xDSxWLKl60/x
Yb5vhGtGzSfJvg8wq5zPV2zSJNLAy/G/U7m3BV7LL4bs+PiHv6p806ME//c6BkPA
2RMqruYBgIqn17GZwNolo9+9yJke4qLIKka4eD0CHqcl4UCrs1LRePXlbAPmrmju
BxauCYpOwLMv4xI7+Q2X5lVCqfT/zwlPuyb+r/qMGn59CShq6/JmKfQpKGQCEbnB
37q5E1NSxmYNqH6lLEXzNMzBt9v9E5zVZH1Jx/PYZXPsJXiWKaXb1l+JyoVGb26q
U+gGJYsNrefcZ2hOW+RU6WaJEWkvSfg9+np7G79dFIzh+0avVFv24maDJ4zJ7pmu
0JfZwrKzb/8Ls9Gd03uYZJ4sj6gSuBN09Wld3LLTKPwvrHwhig0gCtgxMU0moFAN
/fyiXyTN5tJIXLnQhONxTkiDt/0qaIGXuWTgDTJqVXz9Iho2iUfRKWCuTClZLUi1
TCh/fqCW5gfhoxKGd3/iQzv+NTuy/o6BTvmeGes379z8J1zG+dfYXejRr0QwsgCg
LaW0e6XPd0fTttkbRViBwEW9bv6Qufe2FPxCKYo+qLoBeNSvwzq5Vm0RRQFKJXee
FQ2VSqBXkdtCJPv2WFXBHoUm5MsLrKhc5v2w5WCqEshno0faPEM0I9BYuvZjyfau
qd0QTAMZMbAFjkkUq4dbhgRX+ED8EAWOiOhy2wZZ4MY/1vrFkEiI/kmsqC9+LchI
YVLvIjFD8xda/MiK27L+luvozm5xR9VAJFUHnECft7rkcUf6iP6Q/cspECI0Yc/R
X5KZ33RmAH7lzgwzjxHpfUaXXynk608I+gcwYe/5WgMAClxaDRtM7SWCPCi9u8Qz
JMOxa8khwicyQ0czVHIBpu4bPtgu/YHphf9xY8qP079SqoyFRl94RQjGApdpuMxu
N1eAh5iYuFoBgf3WVaJbnbeXh6DsH/OkxIWpWkw5dV1xFWTo5NgjPW767gkQB7LJ
ApBqjouB0ugRyRxJZeEtf+syVPgPpOWGzWvIlI7c7xnQP0DQ4y2ccYvojoNVdiA3
Pp9u9ZbGKrrS7C+AwdQY4Jwqeb23qQVP0EbBCcJqFSFke2onejK4It5K+tBZrF5W
DgpsnzE8ExkRe8U3pfpo8ZRvjNC/ImT3NsghJOY8UNA04QGf4sWzIXDs7NzsW5yW
9cIwsdajiZmvI1BsiwN9SZES6WBQsLaQnNU1WMp/Jg40d/xm96gktKATwxiDw6Ir
v58hHZvSXuiy6HVnsxEG9opLgNmwm6nFm02XjIW63KM0VFS5z3ui+Yc/SjvlKpdC
NxhQD1D4ZqVavfD2jlb/VRaVXXwAvuatwLb8AyQ7/B14GX1DKYOnpIdOOorOLR8i
4UUHZxsy31MiK0WKYZ5UraoGWITN7Uu2sfwxUEXijrHdFWrkVUvNlhHIBYzpnY5v
J6J5xkKYu4sVLuKMTS5Et+UBrA4u7fmZ1jbUBch9uOyI8uQQA2zkjMjwdq78g96h
Sr/tQK8RnUs5OS7vQxl+qjvlEjNzpAjsVF4fDcit4AGxQ46vLOBKC6v9Klj2BS5M
RZYU8MnLZvZwq9bKG6ZTtrbCfd6Y/od2GoBHV7aTzuQHI1Krvo1YB8Z1rOrWTD8b
6rDWjnKIAZz5RaLq5f435QKB8IzhWwg3mXzuCI8JaFHlMc+sVXstnPti2zzGU2B6
YBntzPBKsaec+1t9sQ9afsWwRxgfIxZGndj428LZTvOwFu0ueHaS7oGZR7s4eC7A
7/5jaz1K24JHEvPVSXz8K5WOnaj4H0InU1QP8XT/DPEIQH42sMRqH67CETgQZrl4
JsawK/It4YPtlgLK9H+gNncz2xWTSmxE9iIGbinPY+dDJB2dVDAVCskHFdFnA+hZ
TSCgPUP0X4JoV8lV8q04njm2FliPb7MttePGbvTfQ3YBpz7R1ptHiWLFPQ+5GM1i
07sX0Fsg1xrx1DGH5i5NqNInU1BGnFWm/SFyMbnGrfLGxYZhj2wXWq5rhE8b2SLP
64DFhKCVJLOJ/Z9LOnc8iLZR5MDvti+75ZoMEG4HfSjI3qxZRHqh0h/jcLJA7i5k
WwJqWDjA6urId7FleA/ONwWuLFODJYZogHecm7jOTwJoRla21Uy8hSX1nwGwhXZk
O8mJS0g0GwImGAWK757J2o+hGtL9XRBa0CLAj+sUI7y7weQ5dx5mY2iIQ+D8Jl+Q
1oWsuaOwnrC4730vdVyiM1oEI7d53Bh2adrHikJIdP98Igtxpy9YT5Dd+7G3GjHJ
SjuMYT6QYf80Bg/xu7LX7Y0B3FT9e1rHL0a23eUYls+mjp8NlvjXUIpvFag31fDR
5cc2XN0z7d5VoTWuRXu9/Dqe8qG9rXM1YiG1I5FSBGFZi/IWWsiNooMf7ytC66Jw
aBZ5wDvYmz3CmLvgz0WFrMqMrQlUZxD6VV3uyqFxS4HrO+78RUyd2Ff/I1sMkCje
27BEVGWvmYD5OILotYzvTlqTxd8m9FF6VuL5071C8YPaj7bsX7PbciYXFu88I79z
yxK81k4KO1GKOsOPdPq2GJNmWgtNJXgHcEw5aCiNqPzi4LlYua4A5+mm+4uVqyfz
Kl88j8rGLhSb4u45/Cm4zFws04BTmViLk8SifQd+KQiVbxVITQKR39sk1+VHPD3u
82bX50otqbTLA+5hE5yHXzmxxepS7bEGl+ZESnTRRfiAS1Q1C2Kb5sEx7UxiIlyi
HvE8eGrMU31QSznCzjYdbvcWNpJCqXU1vmnaWTMCEYySR9AicDLJBAVoQVNJJUD3
Z1QZrFob/j/4g+E3vsIbCoiP5Eu1WNMuiL85XrnXE4sXrx7tlHWAnKUEPCaKxK/P
9aBs16KEFZ+30VFnvFoQY3foBmSfznHKZW1iVG9DngUFkjTD6C8tUuOb4h9b9ajb
nmk2HtTOa4mkLveYt+sZvlKjoYZ0R5tU6YERtC7x6/P/CqZlfeNc5/2uNa/DVuwb
PdM9LOdBIJffjDWWJdkzy8Ze5XD8JzUhVqUT9rcP7cfoDOpxi0DClQ0bLeVq+Qg3
MDgBNbrNTNIdeL1XVdV1c4P30DYdv4kopTsKBji/LUfeDq0w2Go9WoSqm0F5BDCc
8qW65iKUwWW7fOCLjgCuJhvnDX3fHmmE/lNmnFdl4exuDq8d8cfJoB/82FkXk1z1
Gk61jDfSwN6Z70oQaippNEimu+gLEVSgfhDcIx5k7E4YiE+dWeKSrf9FCtg8Snam
IOp08AJdHL8gUC4VlMi1/11GPyK8GLzsz9/XIJPtVbJelgusnw5IeI4lUZTkv8+3
8/8EEezp9X0wQkqikQtuq+AWYTaTypMAGDhsSA46t8X23yp3IBRrk8T2wy0LbAAM
c3v2YmWZcWiFmTP0/FV3BJVJU74vsD9iwZ9gOylll8Qguk6YjQBK2/LhiZdYRO0F
Yz9zRFzx76Qu5z273B4gGBrX12mEfOXfoOm16mk7HSkQjXFERyC7flwzapXEDkeW
eeMnpSEXneoqeamn02jwiGy5j5sGuer6FHqF3HdVzPMVU6TL899kq2g0ZOf6MxoV
y1k249FKueWE0Csmn/D+VeMcvHdxz9DbDOF8xGtx3dK3GKwJpfGiapj/SZSQ/xl2
RmQ0CL8qe6Wj+fdNni+27GT3/8EKULskIs4TmkS/8VmctVSSbEQx7uFfI74c+4wB
JrU30oU4adtROOAOBLkBEZL5xyUW78GAU4B9DXihOzhBig2DpWH7M6vftTq7H2xH
2gfdyGQ84pyKwXsLKdEDpnoXWaJiEyVTf2UgBb9KpJE4P31kosEvjCmeDvs5xOnu
KxMv7jexEfN84m8BY4k6ZnsD0H7ejB/4OuSLFgiJtbjSF8sOYaOF3CzrVOnCtVww
K7MxrABtmobkDKPv7gGOmLQ3HoUSNEJG59uLs1gyIoE0cNIb7tTltxmCwutnE1nE
Ut+GpGSO6HvcR3MW9K2lE7yeEwBhOfsQU+cSpo0gY9SCFY6oauR5+9VRaZGvSNXS
wTYYBc9jWwRwZgAWFrxK6lyEk+ul/egEyILvyrZ6w0QvzpsG7/lXZtpFDLcZCSmX
B0JZeQj9R1fa8EVqR80YRARsFxmo35g5PQaxy37htr6AMFrgM+0U4DuCipSCDont
PUxBy2Je/3SAj6xWS50a0vG64a0ghvy8kfyCZuOp1H5NIYNzAxtxxL/2mU3kNWhq
ikxTKQrJPwjtozI1jpanDkdJQ52jDUyN7WZvWFVr0B4BBgf6gzvpWfROUDoQeoyx
ksy3vLrjGU6oq5UHUx0w37thqPBhP7o3XIbVcmBD1D/gEvZbANUZo8aFxJfgwY/+
OD8kjWMKpkLXeUfBQyP50J+/ofHAJlHaXb1EOPneOWWgKGVw6jGGi/6bnS3lFNPB
Ud50+LPH79zddqWNGFu0FMKZE7U1RCZtI9ozfVb3AWWZbUzl3SdMcca2eg+ZRM0P
DUPyokBUVJCrHARq6AwZVzzw7l9ygZMiGxSXaXkDDFRm3xn5kZrDO2MhAk5FFOSg
hcdFhizTSdfXbKu/CtxxChQhffavh4h91WSLkkX/AYgmCtRJ+H6odvNnazZudiD+
EyLNdncMZag1+m+xGGMGlFxZIXghWx3+dnEWvWXWU5Qk9ZGsf5i6126D03fb8GK0
FgyPDgCDJVp5a6S8BO0eE4bW+pbuXhhVK5bJZeoXurmzeygFKUhFGMbucfga0JgQ
PzkARBy0f5P8mIPOfLgVh46Iisl4dgBYGpaSo4jkQM6AnROuRgUnJT9jO+bSrMh/
TkehO1+Vb1002I+QvYTgRflGlZksXNhG1nHpSNFPa5UKHBAxP7I5/57IHCYJtXuz
HO//eF72rAstUY/0Qh7n4NzkK1Fo0m4zmu+fTflEzxlqjwJgRUnE6es5YOk2UA0T
O3QnMzymyZWa2nWx8JA6XPFcRfGQu+QvcNkZiock4+ZW4CuWIB8aLLiKfy9uv2Zq
LW5I8Ot/aD8fc9QiTuaT7cDhsJmfVOefpkXsj09FmIO6ZwEJT3568KOnCGWLdkvJ
t0OaPQxDaM794No1QBlbVlv5XpbpprvGB6TMOfCzJo9rNa9JffUoQPJhf9mssrBJ
Fd19tyQD0bHouHpA/LoKe5/5l3ZdIzp+W3QHssVDAqARLuaycmsVNLw+mfLpok/G
j3a1t+0y4MBIxt1tr0K9xJD1Y6+wV6FboWrD4YVTVHo71wRAzbHvocBDOUOK84CR
K6eLKejekgz+CUZroXK4mB3rkab55RAWW5tbVG76iuEUspX9YNnKuqIr0KsY+WBr
IOBFDx9EGcWdWfc8Obt1Eej8zWF8iW4uflNn+oAUokmI5Fmk1WrJAl77ZKBFnG04
6R1CtzHmddLGSEUwQiQGxONuLTEOD691l/GDvD4vb8bYx+yVnEpttvV+dYN120hD
MrjxTCMcyeXwNM80nY9hzHqbCJf55xDZPlY7trgrb79IijVN8IA2mPMYyPiBMDeu
Pn8pl/RDE9ogNWc2LXyMH7BGKFB1u/h5S2ajsJxyB6e61F1ARbU6ABtLWUY5gJFS
zwHxNjXoghKf/6a5jkCCd87rDeHWHjNl75dhjsePopydgj4fVzjc/6KVZ++tWDYx
1EI0dTeLUuA6jbyXRMht6hDibbyNr0ZhG2yaG+MsajtU2hACz65v3SPiGWGxgSCY
ZmxX7ptq1iSNfWOzOCEPiPVF965ca9JJonHiAfe4eUa5gSlPU8hpzIv6WEdpz9l0
3xJ5nMg+4Wi31KSB39WtAiPjBgBJ6G04NznBld2WEAkoSx9tlYWeRT3AfgznZoOU
czjuiIclisKexMPg3YxZ4N0boU/9gCZpApkUbaS+9SG4MZTK/OkqkK7cvZ18ycfQ
nTWx/C0cSY3awqMiy8WjxqvSjJNsofCXhl8WAaG2YNJ3nDkqABXBlcxSBX/hMirU
LFD1ZNr/mCdLWfxXREjC3alFmOMW6hV6hIHiiwFHcBvC2iicwtcdeniPzVbAaTBi
H4dsNUQK8SIqjAqMJO1pDrA1oCMGdRwQ1IL2E+IA81VQAlQRQmTgFfZrYL2dwzrs
CHLDIiVuPWTLfcymVCbOUf4Hj/4kU2f58BiOl5LAvm1RPXv8SpYcVxealbFdcqwP
9/IoVF80e1VQrPma8OkjxAJOunkpWI9VEJtyOczJjaK8p6m2orutaycgCs9OKFSF
x/rFOpOD9aK6ybbEfij9fSEizzmygtfOBZlE2bUPb07mGOyHYpqEFUl5ZyFaWVar
3apqf+qZ4LOWkuMwx0G9Lz9oZq8uzYk2xjwZv2cbbq+h8lmEHRpcJwLuyx6jQ8oh
yMi9PwUpU6A0QyHn6gGyJ+wCcmcuTeh91LonG3gh4jV3aYwcrEJo3/mPXPC0lBWb
ygj+abt72YjYHfHxEkrR4UJRBKHJIpaec06P3kdF/BbmBUz2GExd9jXNlzhSxXDi
1So5S1AnNSsAQGQ27WJNvuVDD4g/FFszhOO+BuU5FNOfyyYnNb7gMMXHDJChPH8f
Ib6LQ4mDNmCfx8I/Z5ruovJ/HHW0l3+PNWHWsOGhGpBDpacxn30PtuNKQp8SWa+F
STWPAcWuCcUW2KFEQG/kM+yHyc5f5m+0vuBrwKpYFS+FXHuK/FMXdN5CqOFxxUX5
E6LRe3EYYGNPDHyeMWQPRob/lPg8Ph/qHhbUPRD45vYZgMhcgQ+tqLWdjMeVJnfJ
AF2Tio2gJkD+3PYjwQDWZ/v+hbj14q7K8rBETfU28YdzGBndPYE+a1Algb38VTU/
VASOzwhAFORLZ73PSEbKc+aQ0k3nx2wCTb+316fyBeBMKBkuQHuUsCpAmYd3lMde
4fgylvrJUXLyL/VvBUYAow7dbhPZrjWgaUQ+X6wiL/u9tDvMN8rDDzYSIgJl1x+L
celynkNpKEOlaLkvMXf8UgOHUkj6wPJK1E1WSOf3ZqB+P3aDRpuzq7r8BHAzq+iK
0NjYeBfQNUTicH8fHp8/Zx1sbN8uV8qO5HQwg4aytxoCICrBAqDcW2UTOq+r9fm+
ShU8gq4KBjHjrU7mA0pyYpZdbkqCWr3BZX0POyaD7PfW/5/Qcl/+6aTsERM9oAZf
fvyS1UA9yHwaGu0uhXGku6SFZOoPN/3tmDTAnhFDMgAMfIZ2X23S5xdbmK5vEgMW
a8U0FxHnGaImVibq2xHaz4j8zxhqO5hhAoHzRjVBC2T6QLXnDhP66uiQrU9/1O4r
MHAp3srrraoh6ilwEnZsKmETaRPvxpTG7wjqTpljeCEvsR3RkROXxolbcExaiOPy
jgnMUJfLnUphXgkbXQICFCoxiNimwiDYbIk7hQEwjRbNxoCowD7B5sdMxphMzVw/
CeVTGMPgwekAofQ0wTLZ0VSkC/yDFRaGMIDP/cBIQdUqS1aFr/dkFw/+RbfVnHqK
swK58m53hlj6MhYBLwTBd4JXQXxHIt0T2Ivbo8qqjQnwOvMbgD+KerFpfeiXVqgj
tHjtAQFAYEIcxdZ0JbygXEwei3SSIVkZE+fWHCxKAHr+HxsG8PQfYtSEVKqvlM3J
cvm1MCfHoMHEfopzezmTt6oWAMyreYeE30j5roeVuQGeKIAS/7H+hV62oJZOVo+g
mxMVmznsTRBuxt2axLtk3bRLv5ki0GqXpLcZPMSgCR5NBzK1QVQqevhPoYpXQ5zK
orbEZugu+dHMjeSwDZH0u5nv9M4uIiklZqu2u1/ijpJZZ3ByY9ZZ6kSXMKSvFU67
JG+2NGZoV6yaeg7Csm838apFc6ntNEOD0BJhTesSF9zFKLWDD2P3s4KC2Pp6NisQ
56A8DbFVKCHhjWfkkiPPI6RYYuVzSdZH4BZ75XywOQ4Dw91z2RjfaZi96xeUy1xh
50vHRPCAE/VfUVLQSXucCitjaeHw6Cnr6QwQttQjcqbGdebrUjUU4yqXkg0nTS7t
ylFMLXOlhutRqihE9mFNWFxVyKYf4Vn55TKDKzrKt3FX99TweANAk55PLB9mRpb3
NoJk3Fam9Cyv3l1xQSSaJWoctEiksQ/TFinhNbU1agGMOjEUpK1i8Nu7DIFLZ7mN
vLvh4NaC3GQ0we09QZ7eIIYnvsJKFthxKjwe6MM/SEALJMTxyLogCbIUiHNVgEX2
FRIxRNCvnZUjbVudj2F52oBxbTt4XfTNf3WMnLYtUSdhhmD4vyn4Y80LiiFQRU0m
Lbi59tpx2iFv6d5GyNfHcfzTp6ddZ/+4HVlj2TO1R2k5jUEEIe8R8mvePRuLG6A9
d93RrZIbkG3GegJYvpoM2iB170+l37aXNtNZBlo0cB5szE6+mpJIUMHwNjYlPMvI
hclDzx8YcxzOFfKdNWHnwqNMQJcGixlAf/65fHb17tVzZm3NAVcinq79gEGT020b
qCp9daca0DTy5CR++XhiF77J9yDJmI+eCuUK3W/4CB0PXVX3JhMGMHK5nUhlZIvq
fZDAMgsiJZ7pl3WvG7FFbfTuEMRmDPfFNPo299bwXR0erBEZL9KUaVpPIN0PkK8n
ATwR5axaFZ4vXCKa6bWs9f283W/ZXuf74E0xkKVCAjgmvWZ/L8/9Nr+MuHI4b6Pr
BXpDWYtWP8msVt7L2MSTFRaDBZZriGwHz3xQ9PiBcO0Ml/cFnpY5joLE7TBXnuo/
85cZVt1HnQjh4452nZvkyyiij23fX6/kc6qcMg9Z0MVwloEjWECpiV5ovo+XHhy+
AB8gAEisxpAtp9dLjDPTukzlAiM454cbTq0T//KmCOM9Tcvmurk9VwvggGQBo+aM
B0J2nz8OzpQ2ZksFxImrjD62sylPlHqHpvPONdTcTBqn0o03APDfuCvBXH6ZhNkX
pi4bhPGDgtuAPAqKPOXamb0DyiAMEJHYKwVTw1DWTnIUhwGfrCyNO7itvY2DDZfj
fUYPsssgRZhrL4r2YUmnySyvnCy6FQcXMoQNsum+aB4RAdhflbdpiEFaReqso+4v
6bL8QEADtZo8ekiXhXN8INV4ktn3RK9vkKd2NInOWvrBuBUZEAdEbOC68vSTabvf
dbEiAPv57uOemSu7rr6T87ymYBDC50gIzLt/FbwqaNgEHeW8yYtH2VdoBWwZmm+u
T6N0lWqEPZfCpNTO7XIqCl/QvknLND4Mhw08mnhHDjy7OWRlnODQJ3XjomvCJtxh
E3HMGfkVKoB7vEYIciQPkw27u7uAzUT7QkKb+WD0VuJB6xlj6OxdTP9r90I93gy6
diGMPN4mXXzz31O5QAMQJ9xX0hIU3xl04ZDXVz8tueHCMhPeZ90iLQMZXdV4z8u/
EaY1TKjonNWKBguGSA5DARhW9lkr58sV5B622ray3adch8O0FpEtEgXUkBeoggAr
w+ZzDqmfPj+p2d6YB8gplwgXoCkvRhBS8+AaibUSBjQv9bwYJq5MoqQZIVcUftc3
5PohI4IuAIn6tMm37SLPYu0XetWSOEZewbtq3KHNKGMsGCKg4ABR6GTFIU9wSHEZ
JiHiCHcH1JgBp6gyfcDpLxQhctN2Lm5MoCsU2wx64kif6JosLuqbE6zGsRlUYPl5
lxQdFnLBaCUhtGzJHYQMXTAtv7w3x08/zBPhqzTy0MGUgMLMIkFNnPBc2Oa9jsiC
avlqoDsLwOVyeltaqJh4JYie7iwM+/Qw+6W7Zjh/syh9QCZunNTSgwCz+K3SqkRi
fk7e7yTAlWkYt5uvKO2j40xd6xeEMYlNMLDZFxTzY9vsnmnUKjpDqb/O8qJ+MS4k
VkIuWiAfA4SSkgG9tIcasGyETkilUspJb6z28f0NJTtKW7Wk6Oadxw5TvfWnuzZy
EWjLVnI56SbtS8tuWpal44fcWe8xR02zSTdMhDSfyTGPMdTb3yzuA7elodfVnSmw
Vvu3j3MGQsvciBSkbiEnNMytjp0zbSEDMR70Th55QatNwKOl5wHPgOTX/6IcFA6J
SeOXf+dgdgL/Uhe4k5QGPPsQ/7sFsS+ljGS/E1rHLtMemlOVA3YTnWMRdJ3aLrUH
JcvBCSmNREitHzZ/WElMIkXGwfUzsOrCc7qRmhK2VCSGYT1c6/91QFN2xulD17iV
k1K+zhYNztbBsT07DmCzFkBt/RTMMBfz8Ir8TJoJ7sJ2OsBUxPqZIF44gNwe95/g
B1u8NiyjbmaMtwAgxOuAS2fmksgOggTLD5ab1RihETUnCKoZ4265IE6+r2aaROS7
qFwU205epOpErM/p/uEDqovZSsZXiGFhXELx55kjGRNs3/MXwYm5xHxPhTFO8PqT
bVawDJtkGKe4Fmtq+2mym7m79nlXdZQq8yQ3j8Td5pWC3D2smCusERe/31oDmiRW
fcwiLPgvff48lnvU/jvrohWW4ZpPfwMXbpxVU0FNA+FlGA3Hl5EYHHbFhTvGQK2t
lzXwVMiTFV0szTVS1MKp6yesRrHh1yVCCT7miUrXNMPzpRstPDBVEFbEY/8kfX8r
dCasgrSwoSr5jCszIGFqWPKwp00s4MC8Tzp+ZB8VGbcU6fc0ATNGuhAo2NM58Ok+
hJpHG7ei9FkZdusJ+FZLUy+PwDIM7D4S0z2pgM1FbuYvoCJ7H5acdeUWlzeFz/cO
j8GGbLk9L3yoJa4lXvmmzYN+gRcLTYsSlWWd1bA/IHPB1bSye9NcDJG9Eqt/9t4H
eH8AMwMQgdE5UBb0Esk3FamfDOR4sVQk6BvKN94uDT/IzTMwhGMvWtTPBNF6JJVb
EOb+FsW23S0+3lUvgKjs3Sov6vvnK6Fp3PztjDRcmmfwTgkikQDW1KwoaMynkssP
PnDDFdS7oRAZvr7GRDVugy6reL1DTAGCRnEqOOybYwZkdJxBHTfwY4MPf3+FBAlM
mMpadVjHd+8pVi4Yb93mTg2t9J5aLBOpSZurX9OFytfp4gw7vKcVN724Y3SV9VBs
GPOpafY2Cu52N1AzX7m1yhzaRT501WohZG+NXsBxWC7B7LxqKX4zJJFozsJrCHP9
9ON0TOOyUdI+o7H9ZeufzQGxnflMkt/x8dWkLOTp0Anv0maZ7IA8v4v0aDaY0Jw4
cZ6ukV0M7KAa+t736cSjGa26FnRg9kugrdUZhlbltBonaHd4Qaj3xQTVi/yu9RDk
6UyiqQFN9szknmlNx66OXwN0V4iZwfwNMQ5OQJhp8RruBHkrmGV5TBcn+6d7GDsP
wgC6/Qk3HYikP4Kf0iOn0qjBEsENDPCIC2itSslPoaLIDUclHtsttcmwjc7eorb8
XXxRw5RKaRgK3Q8Zr64rW3WcPNFmqOUNF6LfEwiG2KkKIV2MpCClegEQgOwSPCqB
DD1TWUTOfauvEqaJNDDkVKmB0svkjPpaS3HJvalTAfaUtlIhvifI+6Cns2U3LC7p
5lWcEiuda7BKsbmfxAEvfwKZVW5kQ5OX0ihMtxehtiMJuxBv1lSmavffMed6SyN0
DuYRZxGy3/WWWSGjdywcqkZpI0dOBvxMNbADlB6aF7acnYei40VE6qPyXb44N9v2
Pz6i/uaP5wf/OCq4gJlQof2C1UqhLh9VlHqwzrxriPLrK+tYS8cBn+14MxAJJlDI
oZZwopPImweircdo4hSoC4n95eGCZ0fyJyhU40uFMfY5W9UxkdRKd7oBgYK3Z7+N
R/FpxhJgGczwRXzQgpQ3kBgDWvPqh4G7iuLDIlmpFxvBvkwuHIs3gpdclxa0kpG8
lAMd/HZe7UW1ehzrPzHTXs0T4xuPCC82HfZcI+Uqp20W41NyUWpM69JPFUKjLaLP
ZkBljK8n9Vws6WMPwAcBwrlUd02Xfi9GWI13Fn96Wt7xM1Lb3SHQQ0PdFJGDdb+Q
R0+sovuUFOEW/VuJkiVyns2bhxzU/eVqC8VUnf1quLIffmB+VuDavSIr7AnwGdP3
L4/AAdtuPEmKMjBlW4IW040JtQ+F4ZPbW+BWYDY3t2VBJ7A7MV1vHi0EtqzLA5Gm
AsRA7ZiqI1gyBLnTZlcXbyjKvdBuKK9LQpu/gHmnFbRn70bsgo+/3pbq/d6IHlrY
JdilkW4UpdtzmO+lpD/UEWRiBZnqcISCeDNCjKXmxrpu6M6i3H4AXS5NTm3KbFP7
S00LD4s5dYPf9tfSmhxS0Kr3ppSIdcYEgVfkzHbTH2M3ESFgbgp/K22vhvaFnU70
DD2HEhG+w/P7eW5dbR+07/B6IGQEdQQEQAO3BSQ/DhoGez26m6GZ1PvulUsJMfVN
FcTW0HHWSNfulvVxJxDC3NMNesVBdxptTqH/qfk9yJtGdqpjn2LG63CB7MKbNwsM
fL0eS7GtE+f3LQZ9DBQG3t7R+KPbvinjoWzeAGkqeAfKrTSQ/r9nYoIQg8JpJN3k
LqH6W8WP7G4KAccr0jBUaHQX9srzqYfFRTghFBCUF9AS3V6B6gETWAj4Ik/K6VPK
BD9OKboHRNzrJTwJ/i/aoGuTr5YRi1suODbq4zrL9/Om41CFeZiiB4Im078y0BYZ
w0f8I1Mv3L2pWgorM1/nxwDLUyQU4tz96BYNeC6jtjyw1QDGr9WChDgW9Zu4qT4I
XJejunlMEbdinT8+cYjQngC/vCM8WKMbBWg4ux8ra18MALqF5ucx29iHMhw6jUvV
jNmT51UBgJ9hiL/iiwrNJg1nIkpWqkyIFsiZ3csUn2Bi+Ss0SZIfbqcfc1pJhX+a
Kdbkd5l78xr1+IJRNejxUtkCCNg+tD8UG+wWes+YLwhrHmyQKtU0heDnzSJ6d63c
i+/duQqrc5U+PPaVWQAiGDVEloYJCGPi+eZ2RLhMWztKx4c3Go/JDP996fjY/kF5
uxQSoC/QWpEOfkE3RkC642YKjUACufMBBqFUCViQYPyKJ1nJj2EUxw5TMiTBDhEA
mok406fAwUEMSAm9YKDKtY6/ajekD7/Zi9NlY/4KJaC9B9rX72QRB0IZ/fSg9xdf
cA+EGGhjx8U534yEWB5mcwzusyS9xjmDspUuubl8e4IzDRThNigNGHoPp8Smz3n5
2rZFtQuEQwItxkP3s2Fe3eL9vMyEKpfwwfYed80B5SWRZOsyztn604FD2/JlalNx
8JOBBqPBOtrzmWwDQK5ajpyUBRsyCRwz1rAt664Wmqd+G+5OygtDnoXeVTQojvFQ
PPNeT7BbV8o8l/HUaLQlCTq1twM7pBtJiQVcAyyFMoNUPV10AuseFCfItLCBeuSj
RQ4KMN+05sRbwkd/TmHGgpGjOw/zmwpnws8aWYsAl5vR3D0ApOlFDU+YQvsQihaO
RHjeU1i5ZqV9tgixv9MLfKCay6lAlIRaxzRSZGC4tFv4IObvVMd+Bue7kVxV5gYn
SaIjXiW5qcCmqOpxAdyMmzY1654skEEFJEaRgX+seF+xx7SwvCtHwmHxUeYYJ0IV
OQfHAy50zeU6EDaCWBwVeA9bUSVU90G7wCBoXw1nf5m0TvFBo4v77bGp4nJbwiyu
7bFrErn8gWBT0LDAKExRTN5Eh8juVGY4gQsaL771/cosyVg0XekBeW2SMG57v1t8
qQDfF8QX/Qk40OKFEwO0+8b8INZIlCGNy8iRlX49seAAXy3FUentI32FJ+bt7mSw
d/O30WacxiykOKVJkhhPUR5cx5bXUObHbViq83Rud4FzVa4zmb0XNzcDE9Ft3nQX
AAnW6D7u33fRAvnM6ta8pBgSpDMZEI2eo0bd0YwOYiH96R/9dSwHrjmnL4kgnBxr
Tdt8xkhbw3CHgiQfm/OqsQedmYOBXSQtdIq7Q+NTmAOg8ox45FXmW4Q2fYDeRUAl
R+5lslst3H/+UCeERImhMVJlIGZz9ItSugU97rHvzEK4GyTSpABFbq5biEFEF9XO
0wasnn1yBLeUZ9NL7RGsOKn7fkBvQubSbL9mqB49sc28M3plABjdGOTq+oZdNtep
FAnuMmDWHh0+9RvdXQWYIXmrSHq6Aktqr8dAO/wq4a3g6vR2qAfAQ3a0RQIj3UgW
7p7zhbD+gvbEhgpiP31ulVZVBGl0oF/nOnEqfS45oJ056ndN3cNUdEU5wA7noCnz
647qsaLL03kar1jbWjWOWOtFBAze4htfmOaSaL5Q2we+DtVaLagVo94r5D/Alxmz
9j3ErJ0LBq5NpgGClvy9O9gUJ8h1gjmvC72FJOIG0C4hS0mbqubcmpfjuNabLL/F
meP5CsqLKXiJYzxR/yrEPbH8r2P7Ea3ELF6LiS7YYyU+ZtDe7a+fXrm+Acg+1f1s
imERjS6BBOSK+o/cMYdO6M8PnxBvuSKCNzUwUUnVpS6OtIrriIyE6IoODpmxMVLo
jyQdeLsKLd/jDioreqJ0vJb+72UmaaY4iOXuvpmNkVQsJJPibezwurCoMObVi8lI
KMBtRaVujRzHsZdo9eQwS6BfZKRpQfC5ETflXXgOxEj26EGENquMaD+QtTyZTE3u
2XLO9sdvGYwRKrkqRpfjlCNlC39y/GweyP0rugJIenw0e24Ol6+ntlS+IVrI5Tz+
LrCVYKSekajQMKOpOQGZV5NsvpT2SNV5g3byxXpjwg14f6YqHl7ysaIZswZhYlMZ
FkYDi1wkDoaS6wbFhzfLCHXvrPi9fNNNUEJXHA/riwJwV2AAtlSwI2J3dtQG/csj
7tZBitg9jg39RlvWhKaC/nASfS5bFH+Ky9a7IatZqc52tFhcYaOZPlDorowYK2LW
fWkBRE217Wd9DxfPpG7/6BN+kanSguzhU/0YhepyFCQhOVYPiJJpU+xgYkN1Pooa
d/d3Z2rr+IgdA9zY2Gh6ny9aukRW3dqY1KrzPeQRxf2Au8j5YuYh2TKCqu7P1gBj
pzlVq7d1VmcK6CMVIayGQIaS5GodWsvSFELvOk4nfowA4JrOdj/G/Pr6/0TEBXG3
e8bURO6NsMAqWvBf1JKX+tRLiznFHyBx6Oc0musaAjV33UOr8TN078R19Txoa7wA
d6tFR3pxl9wUouVZGgFZYg0hD+kHwmnv5LWKY9cZUBmGFzEAnOEwh8sKmu+tHCq6
edL4ieYqHs2+S2Nb0JZNyPVpuECiOk8w5+3mzYnldILsMKHcnlgNp9DjHjr/pDlZ
6XnRLCGdW0zjMr1PE+3JuBUxil7gSKTfMTCJYcCzEtMWWwtanKS2AlKabxfLdyFy
/T2a4Vl06GLZ8/fGVnLVCeIvj0U2rNcPGPRjfH+7hiS0Vbj9Adck8rcox8Yaa4GN
WmR37IaSFWfinrYF6xhAlwIRTV4uhimxnf1M4lSIWclP71EHm78n2OZYmPA++eOO
xPast9LXZBwgO4UUz9AEvR85rLQnwF6Ch+t+gK7Yw95HceaG4A4jwNTsIgtAjpJ5
FXMrhPWaiY+4mvmIhS6he2xpaCPwBgrKHiG/Ss5P4/H9d72AiyosZ2FBA0wAJxIS
kR/kgcJ+Hk+821XUQOAJv4M/9vgJd2ZYxxXYUBdYkgMyNAytSaJTxgn4pEUWdw1S
XYw4dTV3TxqemJ3gdhO1F2H9ObWmrGAl9fLo7OrpZybYpm58VImFHsAULZWu2b5U
OsuOk6fq6nKlgRNlJGyiFbgaws3wqpplzqjqHkFqbNCi0dO++Xjw8vwvsHSPf9nM
YbRtJ7MFppXGVJY7sQjChkc9v9u7puog1vs/G08GU8rTtEo9eKgKNL4aGxd5bTp9
1OAJ0N7PiRQw31AI2uFpVsTee0Gsk2Z6OOrcPCrl+0USiiCZJSe6jCPBk3aDx9Wi
1vu2jgg+ZrjNyvwGct2B5g7H0IOkbxalCVD9WirrPuEG8GZO6dGZog+S66cQGnX4
QrjhijSDKM8wjDKnzRNYizEalG8AY63jfUH5LKw3htcpI9DBoAvKSXaXYmPWFTBX
vFqJZj56yMycNPlNUDg38qofowcx76hASsyUOSIofZTR8lqnyM6BrUYFFcVt9JPr
hNy0F+pC7YctIFEIB16cy44KpIMH6tNJM7/eP77ethRJf3XbyMVhgsemXYvShSyV
NflZazQJaBPsD/o+Jbg8RKdiKQNqrRHzKrAtLeV+otaS5RbiP9ssM/2nTgF1Am/s
W7bK/lJv9Og7nq0cnrJ2bAeVwYqFiBQnXH3DIymp+ZZwUlUmN2eBqZbDH+CsxNA3
o+7XbfWoxBIyeL8IPWpl7Bpp92KxHTkNn6xo9AXnqT2McQC/lXBZw1FCyToyjPuG
weEeH7hTtF1zArM5oBVHdvPlB5AH/rt6cvKPWyULONtgwyOP/Erm7gBudRX96KPi
GW+o+XOOMW8zcEerMGsS1Flx9pM3m89/2ByJGYUko7MdmsJwSwl/LvW0JRkquPQS
ImFMP6HNfPLjcn45ktj8V5jIbGTBpVkecEaX3t+Xi1QmccYCX+bwul/AjMJJJbK1
XIv1g3qLCNeBCyy6mpESW/XsFbxQBpXLr6DBtW2+2qwGQb48DaleDQPg3m/1Oigr
1FlxfWLBZqpEpZtdCJVb9O3CtVA25YmmODCr6xzL15FGXY3tu0MEubmlrVT0gXd8
xOve/3azZf5V18XJNHFPDGsY6ONwcaV3exSvvond00sw/P437EhgGKKH/xIGcteU
UgnDNM8YhMfrPAvyfXAJ7JCeYRelkPI534lnFvNtxhEsybKldubYQ9Hh+5Qm5Frf
ovdU23C/5kJRA6fMbTy61eJmD9iKnrFLf6vMttHydDcF3RoT7eLufprL2Lf+sBBY
bhophZNFPuhWLE1WcTozWM1Yfz9ckruuULtwkuSM2jYBivW+G4pfQ39raGGeKROg
1C2TI4D/gkOJ5DXsoiVflBhANpbwxeZiJ1KeAn1UZVVCVxB0kVV9GWfrz7zv+bcH
KmtVIiqkzAOZzVhwclIFhdnTXgDyZWb6u6dv74hOH0rm1n/xycyDjuW1NfFXPoOg
fvjYaTNQgfHXfR7LriyJhcDWIdg0UGmjmkNn6cT0jK8Bz+O/0uYXloDFVlSKtJBI
EUPwV3x3NOcHUGGeqY4yVJypAHmphlQ6jY1XaeJGgBibHrPpH5QH/X3ikbA5mrZf
TZsRUAQWgWXgDqy5u1QNkOmhljf8jyLfmZq+DBAcc5RtnXSFRM0/baipdZildzzK
WSjqFh/sZxQE7ubd3vvlp0tf7qJl6XxpHDPLG0oGurX6PPU3cCPnx0KEBH0aoklt
oQ530JZTKqIwJ5WVC1QVg5kDqePofp8FRIRZ5B+QiY4fOvq0f6modN18k1XhL+Rk
pgZSusd9E6ZwQF1h2lLfK1FOXv3TPmfiFXp67vC4mJDP4jHtsig8ognvEXlzVoNn
LTdWOnYipXUpqrz3N+OPlRLI1Li1oePvQZD79Jx1jjV2bDSMTMFTq3vw4vCjxEGG
/3iSumbxmXO9icgJesRMDVsNe05pBhwQ+cI4IW6gmZX9l7JwBJjG9PY+IEuBlPDf
Qk5/z/Jo+bO775JUyALzwwbwk9HYPrAdBMpWvHpMONXszGqckaLBJZAlETpHurBq
j4ihdPQ5rBNfKITcRt7nV+OJbsrabGRrnd4HnKxpYTobneggRHRw+QVn9WP2C3gv
YsqlF2TmEsPiXkqap7SRx9SHPwN2FeBZ7p35I6XucG7jbC3TZ9Af+YLdRrwjNX8k
+qtmR+2B/rcSKWDQn/ppkdfVu1FMZDjqrKHWYKNCAOsYRwiEpKYKNaTlWvdQynBk
qNR65WSSm/xS4zZzPWEscQCtDZN7TeEjbo40O98FIHfbhCSzFOF7AtaAIOOlxw6G
ttqfS7s2/+Ku005ANOZ+RnDDyBGvly5cvS30jAFb3ffSW9KEbdOmDqprGsKAzUn5
i/OXqC6PFRSZ4A09E3Fo2LSperL6p5aQPLRo7ILqe1VswpI3hLayeQfQQqNM6W/E
yamx0Hkscbg+y1e5KbCJ1itwMkTK8+7CuCqa/yf9pqRPMOZud1dVvRPBzuPk3S3t
jdYeTcaE8JJKrqSqrTXI1Bqxhft1/6Xfqih1TMIwg857VOypfbkY6kRXAT7wNEX+
ikT6u+SOiN29bNiKyxeGA6JMfChPHcEJcjdYabgy3+rsrPnlSuDiNtyr5LsjlCy8
MWmKRrhaTxhPQ3DfMOGpZZyqAsOIswc0pbXNrm1NbopNurQEPcO8C0DiwQTuvr9Z
Asa64TPJWIlFJ3GuYoPj3ibQPcgyyVkDlDL787ZaOY35jaUQl6ATkKR+HesJyYKG
WJ6ZxWm6CTxeZdSrMQurVh70LWEtuRUB0NH0HI1dHact/Z3sY6QSNN9IC6Ps/asY
HWQjUOlz5FYjIa0bovFzpaASjN85wpQvFB28wzqXcYQv3Gg+NTTJrHOYlzlKxJ72
4RlOh8LMTqrITpr7bfwRjPA9AY8o1IdwW2cq/FydQ1Mf2rsaeSTyxIi4rSUoA4ul
KAn9RJXl7HopiOEe+S4VWkrxtcIUaYoLuUSwSwZEbAqwxQFI4AUiTatdt4BmhJax
wljRYfymCAyBLCZ1ZqTlVJetYIVI+V1rvMEAEtStWRoAOhpmVhfnSpbYT27rQAig
wK7GkAvjGJqk9tAT2PUaMLL6kRmbpq58vuS7X4i9z51HoD3jWOXy4otg7Oel7b2D
HpiuAVmrnnuNCCmRCnJJxbBBPFITFQaUxy6ziky4JAyNey6048xH3nahETb1RzDe
ncF5HHJLAe3sPJmCV+PNaFdUibkEtNWFCaeZVbVT77V47A03BRLhvkb1GR8hYVBf
wrirdd3B2f7xuihhfKOTKkW2ZXfkypHhg5q0/6aHcZ6XTZW1N/O4Zix64zetQ4nq
EL7BcuhQ0FUb9VjpvswMtGYq2IecRv0LKZUeDgZWZ7vgpjIt2z/UlEA0wXHga352
cfxYDcYVc6TXnEaPrpoP/cMya6u0XY2IIO2mJeI/JEDqoXRpcC17gKTCuAiOUWyE
FIDGxci2T9dxtx02t43yaM9eZ4rPJMBzeAhGAgVPzmqjt+NWW4XTsADMG4GFOWLS
JVNiGssjpTAJsIVLCUvj3ORPj1qLowjPyexMLcuGD20SQ+qdol6nt/ROqRW/KLbA
7/B7Vr0KU53JHZK425fjt/dCMLcBA1cJl1DQA1v9J/y+NDij04zfKxZk/7hIM0Z6
TxFrNO/3q+3gbFgjTqKp42bq+JqkGQOqqNz20xIHJE7/4hO+tj+6/Xyahm3vbOGs
OO8xFpIcC4Hdo9DjhDJh/xNVis5QvJWOQAsa/fmw+ATfqVDM7xQIHIqfTs0KijN/
yE8SqicxwaQ90hXdmwYakmsi/1IahONW1rzfeyTifnplAOnJfmaHBQbfzjVhTncd
Y9eq12uYt/A0USSYAb67uuU95pF7jDk+8UtkHfRMKaqEVOEIXF2DK846Ccpbk+v9
/J7kKl0MjPsyTu36qnLa70wqdJvN4mQERqgysU4i9wzQ6zjuhkEdaq35cm/jTXjI
4Var6Sy8Uvy20kqlYpHywyXJJlIMJ3bJ/ZD+jGVGSnzP1iIe1n1edkcaHkSTfSKX
HXq3OejvH/41us9ldPkF+b6JPmxY935k3iAF9HbcuyAkPc2aRUihIpgMYkUd5TjZ
c266q7Bxov91cVhFVN/kHCkedy5uu6j8oIS3f4ZkAdEv+tb3wPsl/9asGaFVS7PX
/Dh749q4DZOtjRATv6lMdlrKZWKxgLGjflmfysSn5CAIVUfVuWHVe1lVTBINXDxi
PcJP6PkPLjuUI67O5yFgiBFxn2fHAwJ9z5llaUg8M3XO5bOUkVOdn0ojlTQjSaJP
7mcR4PPil5GGM0qqSVTUCcSrxVXTw6VtqhYIR67TEyh9WpgP4RJO9YSlYTfM1qwY
N6g6Sq+48s1n8MRVzTfpciTP2rnN+WgzYrobuP88xGHoTxtpe2CFiBBoS3O0LAK5
mz+RTUn96EEhjb9RKrcAlla9WvM+MuBeVdSSuSGSyx1tN+pk75sRr+eJpsx88hXD
4ja2a7xd9a3yJ6d5Whit90Ir8twmjBdI9ZauNZ1ec//Jv1p4+PsBVa6jgRKAVwbh
2DxmsVz8Om28Z6YaRC7OjsYUzwQu3f4E75Xd2vRvkAf0Jv+j/EWGu1ah6kAlZZlh
2zlrmYPvvatXzb3lbFvWpJj90ATXTUcGv6I9zJqCwIoxWage13/sO4ZNFsQfia5d
s/ciSBaHsMMbqBpvkaeEUZT+V7rIadR09xcXhyLibYSs2Dh9gVauC6Ig9VWHwAW4
FtxM85DpHv/6+j6MBLkzXTCTW8axVXGof1AfW6SQ0uVhQQvzKXdlddCoaGzI3Zvz
FI3AmHUjTmTFM0wEGiPOgHzbRraMRvk706PzPE2iSRgn3MiMtKA5bvENelWK9e6p
k5/mwEqYXDh352IP6V5hdhQwQbvR9bdGmdhUMHsew/u2W0NXAvQylfEu4ZRX91p1
0O44LYWNuAWwmDsU+YZ9hS/FJtgB1BijF866695OmJHJbfxPBLblKG1BVuXSP3hN
FFGBSPDm0X+SbyorPTUrCCVzpSHo9uEig53mPhD+WUFzzVAPstcURkEHmA7K8C45
V40At7gBWamyCaFJwdAalmL5Qs5gL3+eH18Vfx5ftukTzf2mKgMwkqXLU1QAcqQH
SLEX1DRb0PxFthGbo3jSazhYubaRZtWvb000BLAbt5QwyfhAZ/smZxa/5x2C4ChG
R2qdzVldNhqmwYKKScMAJKQjCadLscru2nsnyqmeLFFzd1723ezy7w2j/DPxNZME
uCpqpMPOBQcpMklDPhv1jHE2NE++9euyOYP0FO3slMBXEg3JD06DcjJt5IXaMgas
xt8ELwCMtrQYF9O3Y2B/6j6+BO1++44uCiMKBIxeIB/kj34u6BI3a4Ty2fNBKNhV
KrAObwigBb5NUUXUedPFi8TA0SJ9RxizKgZrE5uKMFmMuMgm+WVvw9tt/POoJUB4
4OgJ6stYo5ZpEd/FyR5PqRHeWGMvl/TxraqlaPK99hfwA3miSaIuyjL1cYcteMCi
cBzkeE/DTl66WU1Wy6XsDAMfyVDJNtUVGfjDo9QlVZH/rQtjdofgj8woyMWIjAWD
ZHYt+Fk4xCnKNhcReur8pdJWnv+hos4NzbGxfpgbyBFV8xK1quf7KxBQMz6QjkF3
smPX6nI3ZbkBfNXnns3SbrVSbQQyuns1U8W1yBd6q5LqvujjHSnJBNnXn07irblk
TD9RkYHF9+2n8uI7x5pBfmKprEjXovtAwKRgdQXDVlkRtViWMa1n0R9FuR16++jd
UvUmeHrdxvZfXA3fUV4qdoKmDJbjzLLM0zVbeGmFYWikAcFXeWD4mVB2QpmgAQSo
NASpUc1FbCBvxhfZIugcSxFauDrkvW85gw7mMQtM8yEjvgzqxhiudL65w3m/4ExS
QUzWCUPP+VU8kYWJRv4VGLoqRh65sV4opGU5qEC4eYiF1xXLQu1YZa0M9qTtXoN3
X4m83N3aOFkZH5gVmsdoqObDEFP2ht3XiZElFWr7HFFQQlwOSGk6Jk+1Kf6mXO7Y
7/QyodI/wyw+WFT15rP4vkTrP+3xKtrSwP56z6G0aIMQAKfFCirSo/NlnbJHktrb
oyBlC7reP7LMUpXuojEtkjGrq8rfn2EpvRBvASZedt+rEk1s5Ukg4kp7lbhfJNVv
e62paaeYUACNPc0uvHSaKzv4eqr17GbiARkzAsJzGPCM4Bv73oAwNwJAm+p1h7tg
x256abztlIL+HR+fM1+OD6wQ1JHImh3CeTo3VY+256d4Rufblke7WEumjUAW5oBy
MY1fkQzdwXr3aspyS3wcPMzghdcmauTNOAozSO7nMUKT4yiaUx/vuHQyJS8TVxeM
Kh/BkeQ+wujSQXSXO/8PK4X6m2CQd+n6sPDJ8+nbgfd/45L+qnXaR/hBpgKSIG/f
GWDhu5l4psyhRfvr6QLW7+XoEJ3aEBrBLYnrLd4BJ5XG1MHA4iCbIlodJ8UoL1nc
k+bKAqKVYLB+qAMprWM+liPv+FFJ+tvQAOUltYGUcz4KM/tYurMpDUS/MGNGNF2F
mkmJcC63qoIufJI3XeQ0joopL4R5kmz+roLeyOwHTDc+J9YoGZcqx9RmugQbZomf
N/mX1o/wzUZ2dPMz6kB90Ep8fbAqt4H14CI/IA9ZgBG5t+FnweEHWUSsayYtJuea
lKB34NQOmw261scM3mFMrxBph/oEm6kU5p5Tbt+ybStvo4NbILT5HHdInvoQ4Huv
FVs4lY1zEk8nB9Gs3WizYGe3jZN+JQT4V6ctztn4M74nSh2C+DVPoL351BmkOkt/
AiX5JSTCTD+fESIddXjTk15AzGmbbx6YJMa008nPlhePEBj8dOufQX/OThIUAacY
zmGe1xbmi5DXPUL4TCM8U21O/1s+jzAZ0cazi+5GFJWsm9i25CEgTEZ+FflJbah+
db4O7Gc+jEFa3ONIfxD+xfZLoFroGo2WAbWNC74Nk7PFs0qgTCPIV0NcEe/OOljg
y3HRz84ruU8g+RMKiGXFxZLsP/fE240uY5/dD/HJqqSF6BOgAAjrIhrZhN+FdPym
f4komm1q3/EINB5vKXmPMr+EiYwsYyXsCc/R8KF1pssaRqY7rnxidlEU4ATHlPws
g/U4GZmtRUO9epgYqoI9V48GMEvWVMi5WUJpZU+KO5Y9Whi16SJOW5eFCGim+FTL
/Tvdzlr+AhpLpLsIP2TljxgVEg6UA2Zxa6CL037hKU30RPhFxOXzWiCOuA4pHYDj
VlbBr8qHZKJK9+KL9hFpWnLuGler3P3qXuTrXcf34HRBIaof0OCzLvCgkkwFSxc0
muJQN5EEcj+LChS2iBjC6xYIC24cTnBH1opNzMqIU/bjRmxDlCFk4CLXxEX08dXs
lwrxnnczle4/DR6J9BwB927lVXbpaWbSeGZT2TgZgUCY8t83amvKus/RpJhBXUYA
Pu/QznrNDeTTm/JhZKPEX4/oJr9qXJgJMjnav1JkSOIDunfnIvVnAUbhEXsKwRyp
W7Tet8/1bkAoJBbYY7bvI6im9frL0c4LEzn/Ai+k6ai8rzXNPt9dWD+PSkFmwOuD
bhXhMCUixa1pJMp8XdgvI9armUEDE1sDC2Afa1HuhaeMiHUullOaUwDx7GoP5o0W
ROyfjgUsRGGBLjChiIKOr1Au0Q8znQ9PHTpnlYnRO5PrqMywJqKMXej8aLvzyXU4
gq1Dw9rUk5whSzdoh2fH6mm1ag1UA0ZHdeL8EY9miVYJeW8u6UQKpnnEV2q70i4Z
mi2s6273deEGRoP8ausbaZIHUoDHmKFf5QpjIpMZIs+5Hd2MTo+JhlqiVTPCE+Tk
HSrtT66fmso1HrwrUpeHJ0usvwCAShDugH4xFXclMHeGwcVAH1zOCOkUz54cp+rP
/Za8QvBMVQqK5gAjEJ6jhWDSpmMAPX7nA53rVXMzUWwt2KOqUhH0f6ICHd5EY7gy
OoxB0zHd+6npUmpgtYJf3/aVUPzpOG1AZjOTJbxGt6OG28TSi5MJXgJlhhqtFyqH
bP3p83hpHdW/NctW1e2Av6BZnQ3SmJwuN2PuufpS3mtYGhCSXl2LX78z5SKxebSY
30e4SJUh6960p3TlQWXiqu1pspcc/2eAcC6+yU23aUf78SrhRx3hjRUovlFadJQ1
WWwO+ej5jjAoqOC9GNhfo9c5b7ifvzITvNHQNvlBe1Dnj6+XUD/VvA4zyBnkQZOo
7fd5pn8Q3cF2OccCmB+q1PEvZEy6xi5kIRughS52RHD4drwBop6INqgISxl7XnXU
wnJlS9HkSkH4s7yAnlhfE9GhFL6ti3Uw7PmkOaKWylBCT6lumiuIEiWintKSnqD9
XcYjniVZRQZ/WWVS6X2JXy3490rjCEBtWA9bXgl04jNduMgsPYROEsA6MTOnIkt6
8oW1IXo+lItkCrmQQPiqM+dGaUVSt5FMPGwlP1wv80sQ7ml5fiSiGXBobqBgq6gs
co+Z33vQLiNsg/6tli8mLf9tojld9Vt8Pzc1OaMnHY/VoZfS62jCxefZew/PKBt6
VGXKfb6hx1txiwrWzXMbDInE1yhinmNdj5fz5LpLrlsbhOelpCPZzsvZVk4ZoInt
U3eBSqYO5KlBnBf+tfItveDcZ6z7DTPV55HAvcsAWobilGuG8QpR0dF8et9bdFRj
bqo1gm3cmqFVARQRtA3UOt68D1iSgJ/99tuFs5ykZ3WHr/UeEqLqkcV8M4iINoGh
2JukUHJbPR0n6UmvFTtz42KtVExLhSJyBHxeqt09JezAwxnCjQnwMeyuo5dwPqGJ
qZiF4JAdCEP1f6/aNDe3xnK6domgTAK6DTa/W6dkAS2srIm56d20QB4PzUOJ/tq5
qae2T8lKsFucyGVBA/oSQDFieRf+yYohytIYoWGUc0Ajk2AHtc1Td95Gqy5RI5yR
+zSCs0F15InfNBBZrAn2uD5kQPiSV12bVMAZQlGc7MZTK862BJSB9NE1DMmzkOpu
vKEwcNCBj1Uhi3nxryOg/47SAQfcHzhRknA2aAWNnge+mHF8L+Z0KrwFqAdga7UA
p9896XkV//F2pVLgYzEj71g5cRtr73PtwzigTJ1B75EzvJ2a3S5Nw2GO0mYRt9Rb
ZjU3DmUXbWxvFZaOEdG9O+ousR2kycfXSWN8f9QT5mx3cF2RybTqyGL1LrWQCLs7
KAstUmgAlbLEM2Y5ojlAr+99AQfSGMjfQ1sFIAIA6mrKcmm6rT6CDxUAv/n9YHeC
Wp/vD+EKq6il9S+tqz4tN5pVGKjLYI8J0fShqejgrD63eun+l81n2k73sYSUOE6R
6BfZHUYcEaYUcnjBiruhqMkR7v/2NB17DIs+Tl8DFiSkUB4tlqTfBJ+nFsvbBel1
3uwvrb5vEVbzelxwoqKyfKUOoBDAvRXv2rTeYvRKx03Y5ijqlgvVq+XrDENnR62B
kqID9Y89wCiklWMsoQWHje5BtpKhZv1vQyaY1y7yBuPbsohE+BPTG5G7s74iZ6F4
7q3uV7b4FHoOdonFF+KDQwsfYiFv+GjojlsJfpSGAdKiUg3YNXBzM7/0bC0wrwaO
5hR9a2ye8ZxTH/4X8YIapzzFQP/yZA3t9wFSY9Mhv9iAZ2aOHtPkDA4NuBbglbah
f7Ww8BlgujPG2puutMzCIjBUjmhe3JnWGPZGBYcK9BsbHUsouicnXAW6HfcPMqK4
A50taHUAKdcSOMNK6nnQ/w1qJH7sMBD5avewOFSnWakBWVddBosF4ENKXExB28Bk
FdXoxLcksIpqBbQzi4zY6wPobTHn9Y5CXeCaqXHzCYXTLRjuSmPmLpKQywK7GiFM
/W8gSAfbOoppkewGrxqKD/nYPdLkiOg6dOH/gPGtbNNr3jA5mFtt69hww2c/V7Zz
c9AFdHTXvtYUhrexvkhBnIeS3nbwKtDPuISX4ZPDZgMewCGML90AxtTaUpB8eigh
WXzNLsUHxi2AC3JhJNfBN2nR2ILv86GDRZXJ3DOVc/YA4sx5FdC8NTWm3yfrxt4p
Y5eKARt9x59zw6Te6FfSgThpSmeAbCJzOL4YvcGKFdUftztHOeKNP7EAeM1iJFY8
Hl5TbC5YFN4n0Psup9EuSmCYvcM1m5mz+RFDU/SDNTdykJkaLG7fRsecqpOT13GM
KwWYZkTULTfGfBWD8JkX0H+taJt6InJ32BMXDj/VOXqnxRpkk/LlChqqULDTTK6q
QOAD2Q/n3bWotWHKL1RQdarhARJ1A8+W9JIZOPBJ5gJTUYTRuT2hf4Nffx47h5hQ
tMbg+CshnPYXx0P9pqT534VzSoxBfcJWTWuj6MqTv1G0MumpSeALP1uep0hR3GNt
jlQnePVLP1oeIRGtRfmvxrDAcjEF2ftWFfQTUtOZ2S1mlWM0pzsvS25j0UF/SUGY
0VE8to544sG2FFvCzd6gcJcQJTc6RDWR8u38c2pq21QFHDcDZHWwejflYgagX+gb
BTIP7KM5Q3sa7ZpLA0OzJsFwoi3zmZMpMvwZgfwCvnyxAxFm/3Xd5/JbTAwxNM2I
Sf8fomyeNlm5MeQQp8wV6cKKmJYJwEIuaVkTp2rvogkcWK/8GR4xV2NaemkKNObX
yQOK9tN0FZEenVdLIqmcFbnfXQKt0x+sXYGwxM9RJWgUBi/iImH9HGXWwzxaaLqz
6EEHODVRo8yQi9S7v7sUkcZjS80OuCF8BcSc8bExn5h8XRfIkMShh7UILcu9fJSW
az3yW8xwd+RN24AGn0LgiWNwuI1yoZ+6D+L4d1u6aWpHCohvegD3zlntTcsVfl4l
bHkprfGw6z97Fi8vVGVnSqNRfxaOJfQ//Pv/P1+q4lsEDVH6qtFZ5K+cUHpDqMDz
JPKsMSeR+4pcbd3FR3EkECeI1470aRRBaIzm6jC5FtP7JTc/mNtRyuQm+8JEyvVH
7vTpV6OUwkS0yHN87SEdFYmpTZtSBOmc4WBCC7LdTs5d+Sm2IIPnl6Q8g6TzdQzJ
Kq5i9Q3nJ7Y3B6Yfmue2/X3vIhyHRvThao6wwcbaI6otC8nWn04EALJSz08b7Yly
AJ1uhXkRftRFeDoBe9sMn98WGpe14hAy1M1HK8llG34xMb6zW6upQSpagbCIBYx0
lUdeTUNXcotqBRIFeJMGoQ+W6z9FTp7AL5cQXFAUDnvKed4gu4sRS4EFA5fL6Zjg
oqM6/P7rbrcXvMEsuYEr4OOcwtFYpBMTNEHfYDF9xF/l46W1QcsoD2JUNIvHVKf3
ho/WCjlWQkWSfHELVKMrQiZl1FREJAst1Fq8LdrsnLASMvkz1uDxufLK8XEODDWh
A6S6+VUk+TPBmddMurpzpHwX1sfy0RHtuxh53y9y8eHbDNQ8m8PHwvOqLLyYK+qZ
nPXvz/VMbLnhLIqCRp/3NdIhckoTrVOkTJKX4tnkHrjKrUeaDNMSdO+5jN3mTOVS
3jkJhWQ5ZtiawosJpUEhc8sDNgH4Ry2EHSqzZLlPJ6qiVlThFN0GVM2LkNkvJRMj
U7WtwGVUMX+u2o7Rulqzb7I6L5HC34ngnd5EMazO5dE1x50KDqdUZwxxIcLoQ5nE
EvKEHdavN+nNGUtBRtqCqKKWgwONpS/psqbvWZRcdYOGjJwHxlrzDTjucPHCJox9
P3Nh0OXGQKB9qYm+mvS4WaVI17X/yWYrwBsnotBLnM6utz6qOKnu8H5ukom6Tfku
WOAcbGCb59A9Y9Yo6XIdu2ckzo98h/x00eJrEJBsoR3VSEc5w02Ic2aNXIfWlhOf
W8JSr4MM7Ep6Rf6Rq5Dw80uThWUA3YySECKh68Qa9JwZTu4P2WV4vOQC5weDegLl
fSnLHjQk68+1Gnqrh65ByV18CkVa0LfoHU53DzAZduEuKQ++w+gcTDmp/ssnWs+g
MhcMsjFhmOXkxK0ZSjod3FVoiKlrh240hWs4OdRWJom3SgWTn7dzReQEUlGozrk7
EWguGbaxttPUIAobNoNU1cO4Oky63LNmdThd86RtsdQg1SHjAvc3JolCAEQ3NH7a
pZIdv81Z0uVm9Jb2fIqUlRsubBmZOGC8SqzYYsqtKghNPvTtvZaTRsKwprt0drP0
W1Pyn3f5ED9OI1A+55Ml5UW3JOwSixn5N3xs6AGkAp5tbvGbXxj5+YpE0oqUllYr
JNwk9LtS8REjs74LXwGuybj9/Z7niEHU/bJ1zpQY9KQ88NSs0G2qorigH5RA6Cf2
D77M+f016Gfzbpuo/yIsN/TuWVXOXMH64YIQ2AwgK+1ljODLZ3dMa9CrB0HHE61p
y+ZnUfkEXiu+0SdXCTEAb3PoMUtTmzOZRX6GAXKBCIPY5z5bcn2T9C0bBNaPq5SL
UaF0r+UGrH0u3NAKAoCi81QAQd1sDilza9VDHDxLiwqw52+sMykrJi1ztsMPxLzC
utQhvbatyqUIzzc8Cereg4NLscJyfQhcQyFMLL5vbIdST/wdIjmTFDUTvnqe41mq
2sRmaL+xqB8lYhYsZSuKg3xCrv9F5OT/wpCitawHJiAprP3NiffjwEMLR6CHgMjP
MHY+YW0I7saJcYnC2ZGKfJgX+BkEEObP0qLFrrxoIDVMF0gOa0f3OJaPrIc7rkHW
oRLq1aBr1I7fciSrUHFLDVVaTW+m1gwNqRAWzgPZzWt0c3VKRr5yDfZWzdMcleyT
DXJR3nMObxPPNKs+JBJU6B2fNVcgc1AKByHja2X73vhoSVKTRb+NzM9iAYpa280p
JPhvAkljGEAIQqPAF1cbGdGNh+dOInVqKhI4nOKwd1qWpbgivXFjVyjRwFNjIwLp
wkXE8kESlzl7iTN7x+Fdx8R4nJGtLFdNXFzKZI1y6kc8yzG82eEWswRYxTUDvpCp
YJJkRiqVuxGg89PnB/XMwbiVLtMcsR5cQIH8JxqfZty5cUCBKrXwO2U4DOQtZV6L
dIFFPv9E1V8bYbMQn0CV8rm9ce4o/nCmokdgk/K8QAZ9ut4PP0qFEzf3E3dtLjcW
INXgiR1G0wa4yhGg32NCIT5hVkWfxhfXgZR4UsX4r0yb/R6n1GfsffO1ko23GSm6
3fl3Ss9DV3cS8Il6AfF5cslAm2FLwfoVMWKMOXr9CG/ps9fj3Q8JCnbMw0VNdryx
Al3hrojxjGH4SIb/ODPD0z2F7ENkY2ht4xQL1dDDwaeE26kT6+BJEZTc/HqryBnH
zpecPf8Qer+z962WkG24gJgYxOsAoheUYTx478RMYwSevC5cZ4wAUrha7PqFRVam
Q5kWHYNTN7L/iuiCUhiyR+qfLOTEs5drcawXgR5qsepUuES0gNUY5W/gHDck2gDq
rBSwgpZTx5wjseTvITkYwlYe1K4R7VP+SUxstMkNbi7ClRJ+redjW1Mr+THBgn13
VmPvXBfLxEXXsek/z0mYKq9sjxSWdnaC5FL9uFdYXCpWum21XtGMmKr5mDuHuf9/
qmqvWTmgGPyIjJ2iNXoSYgY838r2AILdFzpGFwfiDAJK2qwO2z8CGAKvEu95EXrf
rAXpi8/Crw5SpMjThVl9dpBeOfEA8beUK+NBcrcQvquH71D+CCVRAD5acKS4NnhW
Y/rZSj536MbUEAQTS8wivfuczNydqRkeC6lBW8Y+M/KAv+XKiAjBVzCGSnTxVzEU
ds5WgnbyfrOX0FIm4oe2wUZ1xhS+oGgbO6RShRJZwO7/Mt5SFpN5zg9BZPcsZ43e
dMkbB4Y5MZrsTELZCKyILx3AmoA8r+knTigU3nr+jWmRBn6ecCRgLS61fdPhk2/R
iGUUXpyF3ndwvfqw+/4PSjmD5mP1vlr0MrERvc2nYkejY1K8Mg/+DLotLVUeE1lR
UT+8ulxwWwya6Vnx4kVIs/L1IuDDDwQptAm2haoZ1A2KQnUdFLZZvyU/tMm03zUR
PiZMK42qMvoK4zRbACKZOYG+cWk0RneQr9UGhPvAM/2th4jYCODBb8RIwX74zv8f
OJPwRPwIS22wq2+GP2ptjr05x7J2A7Ow0RRZEAP6d/7jBIKNfbejKa7BlWd9PvAv
I5ieL4T7C1sLM3hA9aEtcnK8FwGL8NMpH2Kqn2jewRTm2a91RadiQq6ig+59D0+r
M0CxmMUXK+XY/A+G2c4eW+C2cr1jCb4IXksRpZIuS9QkRDAo16dRSidDW3q9X9Rz
rEVp1tNxYwmsgHK79QPAwvYbEP7DYCUa26uiO6/iFhZSmWpEZO9IC6zz3Uaq3Ape
HzzAbZzhCu6L3QxJfK2+iXhFI/LFPEoJfQuRthEGeLt+7XnB778zLuB9yFOnFgpG
gC7Zi2nf1Kbc47zy6mK6BjB2wYUk6KVXTa373gjlybSexqZXmz85vgqqoY4ClNJf
rgxL2cJ6cEwv0sDLzPPTQesXakDcFNuD9QAttK7bXkRZM5ShI+7dBNUe1skuNq/w
qSOqziDRgea7OqI9rFoZwSozaefsqED2rMBEZ1t8v7bwDgVo5GsyuYSlzN9EbgoO
cJf17LRMrO50IUD1c6Tmn75+IV0diAugsv7C2vSyfXlqxapIDZ25UwpcXpFGgEMN
u0n58iihcBG7ugOkgCkMomcdJ1WRUI+CNdRxNkJ9jiqG0wWXfzVxa8dmXeS63T6y
fjlr5lKcvYpQCq98ZHd/EQ19M/aCtt+/5+8wg2MirtG4ZVdz2XRhI6dSiqeWGqbm
a4WD5M0HrMvjvEvNscV+s7OgFF3KpngMKpY1UR7xC/+iCsx3TVi5AnaKzG2iarJF
TvOA1IzMTJK+1eF9L0zNsDS6iw8U2ouKS46B91qiDqjn9ckB42ARbUv/CcgjwoqQ
2A2cMuEmPtyfWdoe+s3FRAYGnVIc1scdbjqf646Y5Hss/12PsxBnuELq/CzWglrS
dyK6MS2Hd5V5kue5Bp12nlrx5o5SVc6dwzS9TEUX4d/VUS2YkUV9Bx2hDGeaNOpJ
SZhzbH6bBnGBx5m2F3ZsPBXOXnzEnTHkFCB95q7B4J7/kn5ZTVu51IBNhXpnk/8l
Fs+eHvHOQPFolY4XOskcf5kPjp1/xIecEj5TXTtizBTFoB+0mlkrWVUQhdjfYuUi
rpDvg/I6cJNTrDdx5m4lIm9yNn23D7+xlIiY9CMYN9E6FxRr5h9xnqt+4fo1dOGs
nynbJ7KJdBvVpyWzP3ECzsK1nGaG3xa5toKux4xcUeFtZ5fHkw9R6BOrj0vD6gD2
1PAy0PQ5wK2XDCn/N9W9FJnuw9gLi1jw57aBXZQyyz0NHxh+3b25sSs9IAaELDhp
81zhE0gaycLi7D6T2VYdt7QYIt6Fls8qU3J/dy2TPbgFg8IJLyIXXQKkpnVctGCw
eh9dSf0wpMC79loTXR2mtGY7TF/TZSL6/remCZS0tlMxH0B5dsdliv4mGhH5PM/l
Bq2mMf9mtyaPoiEv1AhFFI7JmF+oDJLg46J7cg+r1jwoFH24jTZaPKm1y7sl2OgY
33T3jZFUL1YINjfLPxW+/ox7fnzip5238EMAJZQG4czeIwIrvcybayAsrCAgyofF
vMSAEDIfO/xrPLMlPZ4k0G4SW63jE3hU/oZKq1co7071RYCrSXHm6HYyNxGT1jEj
DyRr2e8c/iOP7u25HNA2y2auBoQJkHvkn2VBQzt1/FvMbEqbdY5QfG2czCK066Qo
/eQOBA8RLar1vAzW/9h1hzhH4QceImhrNx93HKURqkKoZ691NK7dvuOe+/w3KaB3
yY/rBqYvJTc6MebPQp6vfd5jhl4PqsS7DNRrXRVAzuT2ol9EBZTsGvxgJNo7tHzG
vN5pgFmw7GOfx0759TXayoka9pmNNeZcS7NDOp1AeS+uoWw9mRF1aI9sVaOJsrvR
uyQRCzWooD91yAACW0Esrw7h3MatCDewDMsGjKeSMO/8trn5uzOTCdR0GckwOoVM
sb/ZHWC7JxCCqCyUdKdVirwl5sJszW5/KtJKWmqHixfeTU3mSrbRY3wBWTjmnWaQ
VusWWTMktW86VuHzoGvlBGP0es8duNxGAZQVM0/IMnYETgvBobRUBT0FSbYMWacl
5KufmGT94SxphuAPDaFDmLhQt8VBtWkfn+njHfzpbMM4Kn5rEF79oC5YpaN19Wx9
LCvqN08GLbqUph6aFqiTFw1GZH19p9xQxCr2kdINC1TX4jnRzP+o/j9RrYns2F5K
PUeKiXMsDYic3kfgBOWh4dpG3gnkfIjLNrGBON6gYJcekXR8Gb+2JIzw+OB95eAP
K23vX0VKTybmlY+SToW9m3kNV0nt6y8kelrSsV5DqG6c7p3YwVwP6jTISTiH19U1
AHA4cqLdmamEZbTVvt9p09jBhIDpJHB1gVFdIo3HHa3EUscImV3IPQHgPqQ/owJA
w63ww9L+sNzLBd5/WE3qbsgGIRMxo/0R+P4gjleIJU0RJGh4soWA91xVDzBL0C+Y
TsB7rMqqDc/GiIu+ApmZuMXI6pEnElsp0OYiDZ1ylYYkhYbTy6mQE8e3v1H5xfq0
dW+VFoJUCykeeQlldUMabctk+AX31PsIbIT3Y84c8Yrv3RdXN6g/UJEA3mgP/xvy
tUjd7pDAUQ0g1ybRKIXflvnhih5ag+ItxrNtSOuW6BU5zNz2KjOZ/44BlCth6MuA
mzcTn+3RZmBZBnrJvAioGLoQ6cPVc9ASJWGI3eEbUOMEwFOjP0qmGlOZNFKqOVgW
N5L9oroLRkP1HT7RixIaKjwnoxRDn0m1mIZHCw4BeROznYeMJznE2fk9dTuEOJwh
8ophs3gCfysnZBenbkCpF3euN2s08/jcLUUQS2LAiUAAeADRKcopg84aWYtWdXlb
wz7C0BxXl0opUt1uqfG0Tr2IYItPXzvqKGdCNSYyvAZZaMD3wbY001QXylvd7a/e
eSmaWS1BSyOVTF4uGeADYvYuaWxqYclCe9EC5yZxnEf4LBzRFVsIVF6vpnxaMpHs
j3W+KxwWJMozuPi5YZVn+xfE8a73PUQdJZJDRIEX7DFDz3AHIHmA8QK0AxDRu0pK
sRXhBcOlzPK35gknVbMcBQ8pIMwtEISLF+y9OdFCgHFdaX26TKRFoiyEpd34cY+J
7TcP0z6cqGMZBlFUTbHxMPOM9c0InR46Q6Pe2C1q80Ezm6nY9sG/uxYcy6sIWQ77
EaHuTeNlUu6SYBtJWIfdI3abh46kyAkbWp0bxwmy43uEzP2tJ8A2G2qtRBQwOLXG
rhHq0bxx4E9ZeehZwx+UADH5iDrRKOmVaZXVDh66MKzBXhYvrPP5ui5Ci9eqERZ6
4EMm8toO4/a7IykNjtvebZd7leTaLPbEItva3vfBKTdnAjVH4WMExs8V3gleJPNl
B72n+xCFbyIlGvy3TmFI9d7s+CZZ6e17oy9daP+pXTv9IUpsVhxUtSvBw5OAPZ1S
DJu23nT5eBZYym7OaOu51HDqphT6y0FGDMGCo26PgX7NwTY12NIrUePitphQw34S
Sdoym9Zmc2W7gwJUCxqlLqbl0xERgyby7OzLFNlRZeUV/ABkBlHq2IjCCiZeUO1v
yOPcL7wJhCXkraqm0FZd1CUCOUl3+uQa8sv4ZTPTNZFqWb1keAyuSHTarTXUIxBm
uqwH2GhPT1mlMgpSF4PnJdN1QVShE99ILeXCLCjPt1rdb5uuLauTzBcVE2aI5H1i
52i6zK8QS+j/XWmsB6zCMGlumywMlfRN9sss+/tzKG+2f6lHjLjyHpf6ejDT4eFG
rxZCCx4RrDtQWnLYHwc8sNIAneoV3QoJH/xtGg26ieDTLJI9vnudMUGTbIeRID54
B3gK4RqyE3eUUmxUrf1oqYBo/bAykQNqg1pSg2n4p5Um7/4wHoyoN4FmTCS5igu7
PwkyyoJAMXhbqCsUoTMNXvdAW2YD3LHkaqITJ0LJiMGccbWg8HUWcP47JfFOoM+E
0p0tRbbWus8QDhI2JoBy1a05qovrOEoaloHj2PZhATx0bA1SXnXTo+n1+EYdJ0Ph
KeZZKnlHkZmkmp3MaJpolhP605jCfbtgV2F8E9dXN2KVHREVedzy4PBWlsMMG6Qa
EGVdzFgX2KPvw0kOx7r+DZsyG01R2Pbd3mYHLyRiP7YrPG3Pqy7rjkFDVwWj7hSH
mldwgU6wkWTlWN7PMqoIuJ6UsLmqAhK63qNWTpGq5susReAna13km1eDkzu8kToO
DXtApDJ3Q9OV3vIYm0avQpLU9/JC4U9czDM6WN/ZphJU8Mq1WAkqOiz9R+2RhkfT
DOB2mUSKT7kTVfHF3z49TM8PXE4RhkYSaOB5e6q8IGH4YrHcWAKwLXJ3a+R52s3q
qFiywmK+wnxd++6HIvvwFcZBz952SzRR6EDuO+CNDiemPVsrom5YEvQhnSXJ9C8E
Gu5pjpSSWUIGL1+lWac0xQRI3ti+s8hythSpFyoUvJu8Npdg3E+FB6BPP58UTgGU
yCRd9ENUHn/ZikPTVB+g3nNNk267YijOaL8SJJ2qLlCf5AD11Pf4cVvbVtF7dVjr
ExSeQidykXeAgIhS66bfW7w29rzuIlgKy32LkLXNTA+2+FrLYZMRVZqMSzYSRqmR
TgmxG7eTLc7Nh/HsZlDaxXp3WTVC1vGbxxLEcUIILMxHj8xCvFl9TNoiHfT9hUqD
akcJcvHd73E1b0mWF0RYJLI7s6vAG6igsvpTKFOhnYwQbiaigQaU/SnyfT54bGJ9
8Ioaate2kgAzj7di0kQi9w9lX/HRwSFDWS7DoL95vPKjkGHFObu97z1cSGZSvO+E
72Ak/IhTrvi7KOcZFOB6aXCfgpaGXkkqTctwppjqn0nU/rFcUIkdUYDO05JGiG33
u6b2zSw8vJmUvdGSCvZoPbQ6DUxjy4aX9zSLrpyh1HwW1wnchrMl0NQqcSr/yLGA
DiMTLcS/bzR+9ZprlXlXyWmjV8DkZGuS6YyivMH3usisNVcQPjBwa8bWNV/zUhm5
SfZQDSJ9yNkH3wmu2FZbyGNc9ZaHg535CwHK6M9KTrSVifSF82a9zueTey9WIj/8
A8jI2KHfLDmuzbaeNbiccTWqiJD7oui63Ww/xR2Ts8+3Dp7Z0KfHtQpzOqrHSWwA
Mkf4aPgnsD56gllMASzTpLiYvBP/t7XyDtOV3TJTXw/rXDSwyxwJFQHsVQdxogQd
dENV7VuclpWWaQ2mzc6Ue01jOpzi9dp01RyoqAm2J5bzJJ95CBGBwxmF7tZ6Bss7
sgcdOtj3eIvKBWfuVYJLLfi3UMPm56qBS7GHbQMSGmmJimphIIQM+VJDnDEXKSjW
CFEiGBg5o2EBecZHSs/5fxdU73yrjNkU13u5ppRRg7/AchlvJ71d+kD2Vd+/XUKe
xYBpWIwGkzMc311er738/F+Y12ev1PlxVZN3WXF3e7gAjgzArgUhSgHUXeYgkMdA
+mDZ+PWqJ6ule6SrznHunMVXRFOfTLWz6FjfR8QoKCTdYrYDg0i385z/WjORi4QW
shDd3X2zSLVc36vyFXZ4iWPIH9wVsZ3itJRXnZ6CYCUmMQ+Sxk9D6+vDUdRySdWA
PhH8qFRaSW9IvU4aBCobIY3+4lWW3i/DY4wJYeVPv7pH5oMkIdsZk4TOEcHlv7Y6
CVG42Z62TPGG3vpL2pMBhs0C6IRTxrDLj124C88EbqMp5qIaowhz8EJQkRw16wlV
GcQr0ohy0FpNSPYey5dao11j1/Rc9erGZWwN6R14VzSdnZP1OLRQ4m8d/TEbgWe4
S3S1SdBubuAmQBcvo0wAObrLMHy4fZYZJPRYfm9taSop8Pza1gPpOokX1C3920Cs
oG+DtYijPhCJNMc2ygDhi7pZREVK/VdAJ4DXqVhuvD66NpmgyA/MBzqjjebTNVch
/TssFoaCAj3KMKPjZ33FpeLZywglcR2ummWCniE71l0UHt7YYOeuHnbCuaszkyvv
jArkizrciX565a0fSKVhu2IE0StTj8BOmNLUfDuJrhqILva6AD250nbfeMQrDWEg
/t5DvIwhWU5lccL7Xj2CIK7e51MzyDviqDhq0DzcibIwbHteQaHCJLuDrBvqpxbt
p4e71UsnxUq5DvFYIOTIsvUBsTJwFonqvfmdn1pfl5Pr2UnnbiT7HpP5prUyu7h9
qNGuKX0DaK1xMlGZricrV3j8UY85FVI6PaR2twErriFMqXssUqwehtqgdNBfhRTd
c9R0+FUR0nLNaEYBvRq8WufBF5297FJc3h+kTEzIqbxDy5Gh0EhYJ0mLQAI3ofRk
TPSw4wUItLxQXyeHn11fq18fIF0Mc/Rv1qPJ248pHhrYBkHg1P13PK1w0gysl+zr
QhZk8OfjLQzr/XdtGASrDH4h5FTyPuVZqFREjNJDl6zORLyl6Tr4uv/YLmeq2Rfq
z/hDXvnysaDLfjf7omaT/YJZuHSyoE5w5tlu/n/en1SXE/g3We2KOhCDLyHSZGAJ
Wi0NRrAUwFMoi9tc3Nfl45/WZku0kVmMEtu98IHM4eblTiILAHZiQzHODboGSebe
Jf46jVOxreTYSQiUZx/V8IXCpoDVTTUb1XlhZfSGJr7fyQz1++hY7VM5qn2sG+9X
EDzPW/hlE8gG/O7AQTmWaJAPha+l8KNhOKLSNCePlym9Etw4IHtCfcEPjMmfXkdp
ktKm9kJDelhvC+YtZZLD0HKtT04xCfaS2O6xytkazrBr821NJra+0v7ChfDx4NwS
lbbwk68h57Fmw+vL0QafxEw8m2K25zFzb0h4aanfIm+TPwT6muLFtUREL7euP3wp
Ige+azylzWjSfaRU+ck3auC1EQOiCEjkrNVUHnOY+BVGOycH50B0EqjvCRyhwneg
81JCdCriLcK/JfKBsOLl7d0iFy3OGbJs2YhmffJ1tPy+kSxyxr0gQZaanQ1mqtbO
BTWSq/bNwYznLhNSqKaBlCCXPkU4njK6HPmG3ApYQCfjaDy6lY3t8RMR8L8JAJn0
V+1246TiAE6A/ZCN280cMIi3D24TCgBTuy7GpjW5ch/HsmNbvV9dklj0ahwRHjHq
fNnM8KuOLzUiDdZ3OS0PzhAywayNOCc5lcnNo4Y9BJPLDVdIDxUsYwow2uiGDmr2
LDafJwCGLFx/09IAakdBxezEEhdLKynnHENFz7pPLUF9RTwAqdeOphTdZHtPFJ8W
CZtni7in/34LYgG21WM8ag+d/e1Ga7dVggjN+PqZ11OVuNkUf1fhJU4srUs3RxoN
DUwCQPR264XSlWoZmNYI+gEWIKChioDRH0pA7dfRdwcPyhflAS87k59CvNm0nLqU
sZ3+juNX0jknFuLyj8yftomlFHF6x5DJqt9m37UkLG+tjl1eUj6yq9TebEt6qGvw
lRVUtHsHbyJfKlw1d1HqOm/C1teHZxE3iCFm1vC5xxQHHfsK7MTMV8nW+qUUpUI+
ikWF2HuH3Xw6+5AdEOc5oNhHd+B/xk3gtYuw8L2uLTsPyYS7AZ03kZX3cxVYs/8K
bg2rg+2Jwzcajt3X45npJN/SZkwjZxH7dHYrYOKgXBSd67gBJCjK/YaKccy4eXbb
6YTindoNzOKRTLucXzKYMOaGUX//IwV4U9c/aprxeAuK1u+wnB+ojSGVFLWGx0ey
4e0Xza9HgtYpcEmjB3sXy+eGhEEPBOUE9Idu40RNRtQqxAKbHx5DVrhNUPNrcaYU
zJ45r6hoRYv0RtuzGql9zco2cyNJaC7Wv95DGr9W8Y8Vc3zdrTibfqcU51MMpTg2
I0UMYOck53GDYua9qD4HBsZVjB+PSOrETlbgakSQQKHoTBzqlqS9oTytanQ4IbgL
L5iq8sYenzALSvoG3rX6Rnhf0mqP34Z4Q41iYgQh+bNYhYR98MTZ0y8dFpgUXRJk
HObQi1usZoPLjgwOH3/JcIcF6cTYD7pL9mgtww8ff27qkQ1k3N6Q5D+uMz9PSZ8s
SZDI6eGuGjpBDvNwfUdTbIJv6Ox12gfpnTLGLAG1Jv+UCjMNyBRYgrziOai9aSlA
owv/XAfGMRJdilC9f+shmIc5VSybxV3CMlAjuajACG8ZIgFvNfhRghUXnG7N7XKd
C69416xEVTzVmHTeYHBAOD3BJQBJNvLO70Q5Pa+1Jm+MT0yUbOVjYHBmdvxAJKJV
oBvx9qOtsEvop+1elecRB7QcstHTFiNyP/bbw0EU9HZGdB5ER61vh6ZZyUiVZz8H
5dldMJspeghyHsrb9pxdByQmwEbqvGCuqURbWA8ZOV0UOFqxcWezYEdXMSeiteHC
havbROA2TuqYhEEb9ezhNVo6XCU0hnF8z45KgZI08yeWPFuF+cshP1BGoznCBby4
ukkcgrAqXYrp8v6BspljuH871e/RIJT26a4Rt5Trev/jip4uhYO1sksP+PMhkttd
6DseIgbb2eGI2Kz3pmFmi0ek9/3MNtsQzd+FdfIfYkgDn3nYm8j/sBpI92HQRegV
+gCRFqDh9V5zb3ZzyH3vKMfxekzJYzLO4UYncGR6Jc/fWbKUCPbKn8BkIpWkL57w
JFRWevtuuFOIP7UV7PXgoiEnGq7zEoNsMN2oolPKNmgSOV35gg2naAzIeokQdIel
4Zw6I6vS2v0O0lYcd9t42qkiHfyopSSSxml9QxAIZye6FIQrU0kBoCSelDP56rOK
A2dtY/RwePDLxdfaAuQx1+vgPMyimT1++RfzOkOmE5PwJYx69tgeMb38G8qMk4AG
mSXpMP2Ti85dtCEsqU+s9ovD5k9jF9VDpf3YF7k5bET39PQ2ceH185GEDKUr2bqh
8aXP2g/eauUaeHPrtmrip5Tqn30hkv9aFNpZ6Lc6Jfq5NlGlWfdSkBIYDMeX7fzt
QBOZGAaQ+EId05xflVCdYkljrob0McHTWrO7JcqPib3o1vhOkoBGUa2RezEnJg1G
xVDWR4tjVJ6oTFOKphaW6m8jHVH0F0lCGTsMx64t6BbjcUuhkdaTBsVibSHvjE7x
u2wDTdnnYceaAzQtKG0UsQV7LD/VLXIDD5+wk79iuNiVxfgapltFDuiHZln0cf2j
wDDciOMkHiyITnrwJqzL8I7G2JwbzAuDbOxK0DfgWCUIRoPKtrMAGCDaCH5Y35W4
gL50LdEynUDVk204jTRqm8MrV74CVFK9jMUKzCUK8Wgk+apawgju9dP9fsNwiDWT
u7usP30ogcGBG6sgVX8+DK0jci5EFx0ZY4RLry5FUUeMtHZlCImyjj0r7dM65R2O
8fkdX1WxAvKqIqnLlQVAFgrb7TZU68tuDz4MRVuE8VPY8GsyhZDr4alnujOrkifq
JR5euKDFslt2F2g93MlEbehQkihy/EdYrExbXcbz8lB6yfkyytVIqAv0bixDNbB6
XKMbKOc4zE1x1CVm+V+91vlO5aoeW/DwORyU4qze1g8wRbyEAey9XFTQyp67Gijp
fl2N2nCEJ7IdcDjHk0Jm9BQet6ykBja9jKifOwnbfdQT7pLFuSlCbNNl29xtRU1p
Gn62NSw49umDHZMKVzZGMVApxk3tq0d0ni//koH0kzCyrwoQA9W4VAwYAtK7luv5
eX5zTQnVrHMxces1pExoeOIyrdiCN/hPomfPxW3ejOvrr6yesfS96DyN4PlyCU4f
M4Q8vWsIiQwqHDQgAAiWSxOHDR6tvEs3ldDwfn2626OpwOTdSmWLiCFYf9ptiJae
Qip0d5EimEC3JvC5X45K9TRmtiILMHV+K7cf7Smyr2HLW+/lYayZr6AYSihiwuMr
3+LTsaUKy1/9PL/qXzCL3nnd3MZ0MhbNCHdTHOLj4Jra3YYsqyErN9/AY/MB2i3k
TuJNU4MLlTQjsNdxeyJINHRPfAyZt5eoGkqgYn1E3Zy1e+IXTL5XaQCuTIsnZ43P
oO45mOfJwvHCOEkGcSud89kKsQ3sVjyFNLg9EwHOMzUmPTJrlFTGB3ZdIUtV0yK9
uodfiay6HIy8mNRg2Yk2BWQvhlV+D6BlLcHzRRDIE4v3VSi6CVRJuE9AyTgnonKY
aSrxOfasrh+5COfJs748GB+sgK2DKR69ZS2r2gy3anvI/RGz6GTAwk1E2rwY6N6t
gkrJj36iRiO19tAvv3i0U8ZWmJG7/JUIcxsKNjwz9vNy59JiQS956d8Li2Gtp5aa
0Et6Sa6Za6vdJkpoAC2SGhsUFcqlyANDrbWXTY63lbzWe4qLn5dLNN1fAQA9cf62
XAE6H8EpjqHUIf9DDOBLP5Fw9RpVRI9VPF3durKZqas1VyQ4gk3Jim/nlxlyghZ+
Jm4QXepgd4aaUtl8g/ni5W0vXQIfWcJNXOS5/NGdnao2G6Pg02Iov58tFKxgzxlJ
rFNHs+4/3OKjSW/v4ajHpvAJI0y/AOib9H2xyVKZiUe5RJ1iCAaF5+0n0xZUl18s
Y5Cw1G35HzeBBfxJrdhFBYhPUCcRhagsPzWGXUhthZ3e071MvMakRD0UpyQy593X
1EKkadN/8nS+3AUHYQnXDgo1gZeAsxBVsWlXmsR5dNmslfJJ4m0fCb2glop085ls
Q78B3Z3hrB00V5pPwDaoOeujdZybK47c3Qpdv3LQjBcMZj+LEfyybb6Yn1HEPt1U
o8uXbxLHd1hPXtQ6F6sgUo7NNgiRbDGK9b3qh53svXGHI74vbMZIAno3CO3ZQ730
4nOlJ+9hyc2WycjD4LbgjrsAemCugRRE9ZZ5sUuCeFPiBoKy0CbT2MVxGnHa5lW5
+JvZqsCck+vnmesXbz3HHnxdL+J4ipDxoKFLbH0gW33gLiRFr/7PUYUvGKunv51L
aBe+g2SbW9EKizMBAntERNJT/B9h8anSAhCA/JUH66ULRrhUygz/GwvZe6cmFHiS
VOeWTzvu9SoyB9K83XFAcP8rJ7byb6KsLd6QqUI/w9H6gGLhU+DZDWi+o9SERmPE
wXp9d+nEnaY8C6mGQoKZsb0YVKmib/FnTk0krOmozQJ1aU5XydeJ8Cu5UP+dh0To
6mmRy2rhv80S1vAPOImANG4FS9VfFqRdsU8SWo8CFhRx4a/R9nO636jKuEPW+aJ9
vnBmO9HdYw0gPCH+F4QcY4hUpuwTaxAQh30aDya2hOsqUluI+TZy5kc0app+UqYR
WvDWgk3jZRJcA+0+j7Yzv+zyVv/oBlQDYQrynn52OGV5r3LO1eA+kwsDlzZ6zvfJ
SS7qd9Uxs6F/elAeVyUB9xlpxpxuH5isCNR6nFCTiApi7GgMOgALmWTskijP0F30
YdunB7mQb9NfRYKZlNRxHtm22MnECC0wfkZTEgeb0u8ytLNBzok3mWVT52hFdGNN
BV6bQpipUoAeYDEyp8QUql6NFeb5pmsV0m0VYRvSUJIr7ay8AXZ4XcUDDwxsXQ+6
LGh9vgwcpSeMheiNcZmeHPWTpfx6T5qiavxu0j/uCgbw5wHsJZglNfbuzxvkW+y0
A4dFLqI0C9o4sAyILB9CMcMeJ/YHYdOma+GHmm8zuyPXLT630/fcalL9OieQ+nqr
msCHqtdLs+0KwnXRUuDGUULDmPy5Kk1TNH6zCxhygpK4UUHaoRxTx8GLdXoluzKL
LDrCiSxV5dUh0kNjHhfYgihhWzfKV8sRlcarL97sVzK5E5FCqtDEvyi2mfl+17sO
iSlkjTaVHkMmPLvTk0sWLgZ3MmgeVaVDBs2k77zxWlfhoyUiM8344WyaM5P4CPNe
6Uok8BIjnhktY7eHYLC4FmWIAOokaLOfF4aMj8O4ZaSb5gWlnhOVT4OoNwI1S51C
HwpxYjKuRezOlsv11qHSmQ0F+NTB/7l/l3YIIfsHa87cz9PTYWK/ihBy9bHNdk/C
BZNzXtcoibO4BLTlVoZwKaiJUC6pgoMEuwynwZii9xI7U8eH5we1rEH9x1FsZ5nV
DgSE+yKmfgFH0oC+ZXkUlCVolBan1NMXR2VytgX7QoKnM4e+WGQb8pGMQmMz4UeK
MQiM5nn6Ayg8xjAnbqS8b9/TMWfEwsWWJz2PedZMgW6j5QBPMErxLe1a6/lS2r0k
vwMGMm238YQO8JX9FZKQIuPJRbP8QHCeNeVJrllfnWruVtfauxdZpd7jvsJzYaJ7
XKRIyPU1SuqbkeBWhRjWg9umK5ml6hdvpM9obHVRPyZZhTWl9o6+rNFMUJiOL1wM
B+sVjeUvs36fD3EoK7BARxTxSlaBOeC4z+o2cbSsJwOpi7456xdYVhUHc5N0stEh
MXWbB/bzj0PsMujDvz1k1Fic0lEAtH4EkaMiKw+eLhOMXiK296U6T4y7n96HsLrJ
WhgF8tKTlVaUDdxwxQlc1c9atlXg+oN8usZHTBtxYppM9FihKFohRP3ysYnccme8
LEDMAr4fQKd/4eMdzySK6vOgpqO9GJps0xkUykWYUOmPT+CAyjltH4fWjzbqbUTh
gKriDfWZH8+eWcTOTd3nXjokBsR60yxBu7hsWAJQm9AikhaA1xI6BBYVIW+JcRHr
43H2QkkMO0ijxrI5Xr+zu/Jw2aNxy8Vir+CY/b6orXfI0KozVAx4HQBv+J3DsufM
8+/Ce7D79oGF/e6Lj/0+Xn+GyDxIIrGA4tmyYTpH7K3PJkSOji++L6I3TFuWX2g1
lZjoVQ/02+kTaW9v9L3z7ThikreAiA6KgDj7Oe7i1nGoG9bGK6gf8TXsiWWqZLnT
8qJYHQjPCWCuZxvzThy8JBzFUtOgt+ROyAOx2KdI/gSwxbQ0w0KgsTGD0kzo/pyC
K6DEpovuoFhz0qZkdLrnG5vIt+Dh44th9NbCH0WCzkUw/86s0gxlPb/IlhmMk5+X
YldFMknKv5ReF9zq2xuoZkI+YUaTho4s/8xymS1xl1ljKiuTZsWGJsrDB0Kf3ixk
u12RmW4ZhmwctZJv1Xrv/6Vh71lpKS3jdj/9ap5Zml835jXSTAlc3kWXxftfiq4G
8+hx0Veg5JPDtUATqvEAYd9rltSh+EGxuzw+cKkuz6WWkdsBpL9fPBu3syKS4KKs
UsVCz6+jfVTEEYn6LSAp5km/kJi+6/rpAyGkZgaLl99Wog+8s462Yxz0idfBUzgm
3j3b0HNT3vB70nelnEbhUQy382OeEYI8VSTM8m4NPIxsFoDh60kKAh3SyM+MOG0c
2+5bjL2bqgezb3FivJ2Zn9SDMFPXPHwEwdjpnmAmvNsHCzzgKVejP/3u9GWyz0qc
G6DehOPhBXWEIs6fTENsGyFzJwZXAURLEgusQT1J9SlkM2xMGYzWxPmVBBai15LL
Dv19+c38PPQ8kRB9Czrp2rQSe+T171uTDZlbouq2mHEK5lIflCGwWdUtxpzGW16d
wrEMYNlTCMv/TytsF1Pu2JrMbGjpcZWgw+TD5VDmrL/VB9cub6DjL1UXW8H2VcJy
ZN7T0IUhO8wMcf8/NU9t6VXd78c2a85af0WOMgseHXYkMx7C3Af5FK3/hwlcfesV
gKxmW8oHd9N3oxvHEc0p6kb5urL1XS0xLq44e8oJBhPOaEiRRs22qfVtHsSD6V64
lzoChcerUnQYyaXJ5RHJCHWXe1JJH4Z8Wpc43X87GZnxaHm+3ymBi1hhwFYwa0ZU
0LriSXbyqhqpmFyCWO43aud2eX4vkSpDqK+dbBqp8aHLkfbpY8qskBXVzKGRkuhz
j00CJoDFJf2CPqv0pxw5GCocm6Hi9krK5BZ98fIS+IkqmvQ5b+2gXBujx339qaM+
htN9NKOPyfO7386sokSUn3aupiomJWTvTyEZUwdXzsxwyuJsk4rG648EkbYk9vr3
bzgWW+ib2aEBXZy+7idXa7AoEu10SKYUZkrJE3fitwG/CyJetPfVFTsPimZdaJgt
IFztgrYtIJ2t/LlbCs/f02phOPVGORlZ9L9A+Y5vYN1lWYNZ7vHh14QqrEp2Wolu
nX2AiYwxtdBcq7hk8iceySktyY6Ly0vNK7Vn43JxmIvdxnDGP0NCTy6BAwxS73gu
Ib0iaiZFCZDG+u8kBQe5wuXCvdanbm0aWMgahd2a7askC4707RtIRj+VBr0I0e4c
rDYlCCZqMUSPjIkf4JcKGFC2ho4CKvyEu2uheqeDRdHpcsnwF+FhdXLCWYnFkIrS
aN50jl1IyBXdUSI7yzUQLRWIgxvjnEORcN+Hb9ICb3bVp9cM7G+160cyAv4j/Og6
xO6EHfUoBVHwzwc1tnG0iHIMmNCDTU8b1vtncf/FCJDHgkA+UFnSf3rtUJa3CGAN
VcQiLxFWF33MEcMFNLnNay8+NlY+gl0LOiKWn3DlL5I1iNjIqa36YIbvT9LZL9R0
p4IMsT7lMoNNOpCHljIOq2xYFZ4VWwgm50pBJwuN/5x5phEXo5/ZTFhVI8J5nfSn
tBF18f1145nh3hbh1L6IZw4L8hSe8GhE9Oq2R/db9m3Y5dVhG91B4udkgYoc01po
OrEd+JHM3wTGQ8HHJgO+p4mlN4ItGlJ5XZpVvQGSpzIW5rsIY3swDy5pSj13rAXl
eyMHxHF1mJj1VsreDUpzpQ/uH8vnxmwDOseMWBkemV6Wu3UFway8M4HT0tCertRR
3vG0axZCLnVgc7qBQalBuLiXuvj4CC8//uATuk9pYbi1vKEia4R42vjyWV3QAb1O
ZPdD3j+B8OW0rVu5KCFYEVeRxmyaTJNWuz3TVi4Pbyd7ETFTgds0QFm2UTFTi2bY
/ykjn5tV72pj/n0y4+wgZCUMRTz0fstYELr4CSzD2YTmvrlq72tu/ZuJB6pohk1K
4f4h2iHG0+kpUJURDMIo6ZkIK/mgmnFKbyplhW4GN61pcVcLylWthOU+cejuOTbO
wlkGY/Maa7pfPWkaKN4iGIvkdcqjQdUjWvQuMkooreHVn0L/ERjmnJOj22TMDknQ
TL7O3rcYuNPIujMe6Ql7ZUDOQbhPBwz3xoDFTAyYcjHJk29+SczZ/k7ytvNOj9iW
95xCoi5RcHEEr4oiqyrcHWrP+waJ3J3ckjcFem7FmLD7+vvSbI/2t1b/SRE2VetT
bVvncKH7HkFBya9HwWEv8OmQRwQI3uRV3FnRDxcRoJ8BRksTtR1DiK0e4miKS6yF
N6WLHwL/wSFPL88m3tF102NkWrZAHnkWyIPzteC3Byy8hBsfVoW36/PrjJPTeBoT
D0yPMpU/hyYuiLpWuvGP+ROnknCeF0h80CI9pGipEjSA01MGWYr+1aQ42XjD0czq
jqv9T3hYTwh6d2nvLwhiglmv0YMWtfICYrMCe7DA29WqElfjvuR3yUqEQqig3yEv
TO8Q62cyWBTlmIwemYqYzKk1yY4b45ONBqldHslRSFwkf1aHWC7GilXsAUMOEUrH
3LxxnM4A1U5ymNRcvjCZ/NBE4L4d5YOzMSzZZKfqEa53AnqNY6/PM8DA8cLNZgBA
OkZ6RrZ7iegY6RkQnfGVJGkRfu2MdpLoNb0yGe+AeQsxqKRNRoI0UccWv4ZQ452C
ktbiufM+pMMdxIgvQuzDhApwfCYbv/IPeWD1GDyxjG1PDp9Qnv5qPosQZl12U31R
JR3mQ/KA+3adzDfdrnjV/B6YTiFwhE/wPHLa05rczslmu50mpIzfPQtHqXP2qY7x
FrVtsuzLBhULTvz0nLNxuFysBI4tTEoidBiHyTHrkHrCj1rY7JZq4iZCb75B8pTt
JZBhUI16NK0CPBXVIWVLkBAoqoeyUawbRqu5fuRnRSHy6NnYlRlIPOC6owmCXhYy
7gkODkIyZVtcvUNvi3GXKNspuOjZ9BKmkr73oUK+SOd6kmnzI0KmSrhvPZzZsHbX
v6Gj+9OJJdRwoViT177RJ2JEbpWd0Sz/4daOkVFfGl0LD8XOa/aQl07VeV/ScLnP
/P2AQb6bGLf+iNJIvq74mUhRQIi1onGNNFZtrpm799+DDUYzrrB66ij7TUETw7Cv
2HrJZiHsQSL360zHE8JbNlYzoi81RLWO02nDrHE3Nez5kfaAtXeJ7Ibgym6Rvash
gwplX4mPbFScKDyoIHnYjFdhArY8/TxOFX/1i6gG0SEpFJp42EQiHqWWqVIN8AMX
LdBjeV7eLDhK8pp27o+H+tjYyIyP+rZn2rsVv9BGJE6eSIBve0jl3wBpc/kea7tq
mYCT6BwEpDDFormnklkfEnRpp9zYRp0kXgP5IZAJMdPViKO7Cl6SopglsmtLV0z0
2vBJXYE0ELth7byGtpXyLxQ1U2b7Nhpsae+DYqiCLTpGaIjOEtCmdzpyfAffHQhe
tanhn82m/DOLsRHoXsggUteB0xKjJerrS8f6ix1tvSLR6uRTix9LvVy1NH8hquV8
Nx9w4Z+3RYlUXfBfBoyih1BQPwfUOCGZlXEwEF0TY6/QB1zSXtQkvoNxnb2mN9mK
L7FudLng+H/pl8FG4SG2aOu8KJtkQzHsLLivUTg9Vfi9TFjpP0b+/X07Se1HUhzf
M8TPY7sndA3JIaUgei0pDsQ6s6xZS7ipa8mzdItoS+oSjfggHhXHpvXcqs9r0OXq
BOKXQI9x59yAY/liI86hhGbdSswvB1YITm5RLJAnoWVYGD3MapeJuB66OsHIuubS
t++HiuFYYZ4L2/Cmy2ou3EyhtAJW9W9gAgveN3wpKRY2k9eu2ZY/rW/fckMTfHa2
1VRD7o3oUna0qy6of3chP1XJw+hKXoK8M9BusruXsTVZn27GZWrJNnjB7wISF6qD
MJY1p/IHvzBTKufNi+5Lz4v9rroHHj3DhqnWH1bl2p6u7qMKpTphZiEufO2U2Cb5
LAdyzxKD5krApju8JA9yenadYzzYGX0hcd4Vu9mHFyzKH78Jxr6q5kUej9Bx++JH
F+agSP6NC0OuhbFIZEwrF1JG0laTqYFEa5XxjMs/K7NWNVqVGJ5VbMzYrKkhv9gq
h2nKfIZ8BDkUoGC5kTx5UrRdQ7DDTR1kraJi0Ztf2r5R/LzaJT6M7s2HCgGw+Eam
D5KB5Diez2tYc7eQZvMDtSNwhtv5NJ0o45VRONsU23u8EC7t10TFldB0C3INuoO0
4BIwG2kZRT+Oga5216OKkkWK/yloIS3VHcn9cjQEjFvz0LvDuIDwTSbQhKPyv07X
rFiD5yHXbecvjblSyqVdEofddJz/M9pMlwsGPkctzvIX5nUfZKBsyDwqcpAycXNF
Di4l5xqFGKEIE1VsBbmbmAyMXgN5kdU30nLYu6WFIQnqxacGl7bdIyr9N3hSeeXw
l953X6EbsUzy1PF6f+VhKLdyNkB+2OSUo2yKcFsYdPq1X5c3GSbuEX2bT9V3kyw8
/Z5S9ocXjF2gJXz5xxIHryaBOxprr0sbYXODgX9IQKeti0ZkB+1tHY+qvFPRyIL/
1W5vlGW7jo2bu3YSk7BuLGTQQDS3yqEsZYx6i/lsIyR2E6cEcUqTrBXf+7Otv84e
ZB2xVXSRn2SY36N8asMhjViPVPwlIpib0N8WAwO4ZiOozGjaAmnqo3Dj6xj4rM/W
GC1m5J45cza7dWBq6/YcTL1R4L1g7TlCBGPysBMRWBNF/5Rm/3yW5nw2JHdciLyU
Hl5jK78bXy9J/m34cfZEuvjRY0kF9m0Ypdvqmtm9uXRlf/sK9o5r2KtIacLcAICF
rVB+8kq2hWkrLhZO1XQ4mj6B6xWf8fqBclrf0ZbNwpbXMBDer41cww+5EFx8aZKD
TOLQYFodZ1LiOAI9ejkX88HzS5KZUn3MzrpKTWuuYsXIfxFxBjcboqYlcyQw9Qyn
1h5J9ycmnCDN1jcujohQR1TrkAwv04w2CSHmQAEOQ9FYF0cBm/fiJvqh/GOova+w
Kh5Hlj7eCZx/gWX1bTV8nhrHSmn3+n1fj4jHbfVYIWKZCAqXoawHqqVb7UKdfLau
4tzEJDdjuIBWVbxURjGuoI4E4WV4aZGWlJzDC++zppoIdySY291CY02U/bFyxe3m
PvWrQIfWiQu/tLYTQ6uk3kWIOZjUIBpvy8g0Bk3I6JqBtLFPkOgIWm/7ONqN0cHw
qquxbYhdoY6VCgdr7XxqiPiVBq4VxfN4osLj7Kjd60TNUSZjh1iwHr5QN8eSr/eC
rxi6qjTSNrE37X9P9opsblVI6ExShJPQiYpnRP46dEdVqluQzcf0yTneBINzotgG
r9FVd1BtRmfQW6FxoZ/BIo/up2GqmP7Ij9t6ypkgEe68V/yhrROoitbuzcJSyBxA
m/xWxqleEgWrCK+6csOOgi3M60d8B1Mma1ahsXH4gbE15lC4FcjUPfAitmHYGOx2
UC8dcKT8nr+Kp3T2bdLgvr3xRahORyZuYHaVIxgzyLhCkDbvoFY3QDEBOv2owEgP
mjlfQwH6fth79Er1FFVCCg0qKnDw8u+aHYXQ3Q1gUWF4PPmlUU277EJX+H9qPuB7
oCSh8nnlp2hdTR1hYy+d+Z/PuO9YysOa+KBDdQPpt+RZ52iOosrvJRKrcYA5nvoi
jtW9/vRBuh4ttPkpuFXmmpzCR138EzT2AlSgBgcsElkPOQ5OinAYQ+8G65Cvx9nc
FbpPET8jf+FNaqI27I3hqSsfg0iaH1O5Cx1Om3hglCQqe8hoZNdyUq5mAeDi714q
WyFgmvuzLFqYRDbvgNIVRZTF2mLotz6UwjWVwaKj92/x5Nq67vRUvb4TPilSCdFa
L7o3W7jhiNGqLUG8s04Mp7CJP8h3WP5OIOlteEq8szsVI/nLHXM/M0rVsu+zG217
8k+sDQu9s4WvLPbxKqMb6km6GIC6ONl7e+MqwgozoDaoEeTyNqMcS5Uab6tapSLO
Nuw+R0XPSkLlM7BTI/3GUouwD+Y9pndMVmNOr3gwZPukdT8e/GHWQczCiOOujSzw
rjA7DO0LHAVzFDz9GlZ87M+aMRiMa24zFIDGxo4pHqj7DDHEsP1yAFbuJ2Niu75i
h15XEZOoJ7C48fD/ELypqAxGeZl8vK+dnve8ecKonUxOvrXG5ASIVLI5alXXyx6r
4EMKW3RO0090x26w4hLyM8lhUYPCcsV5m9DfVTqtDdVp0q0/wo+0nd/nfuUOGwhJ
jPG1TQ3gv6uwmJ8nQWIKmitIZ87DywGGSaWNTh4/QWxODCaYIjuAGEytdBdvQFn1
c3HiNBrSfq8Dj2qeZxHxiop9yjiav4NJMKSNsyWG48NzNBt6Urm2AC7ayyjfEOHk
CCo2RiA6lx+pVBkbaoGm+1VaKInoPs23e1LZUA7JtGnQMKVsqtogQvc/elpavGPo
RxX8412Az4HS8XzOwTOuwfAAMr45N7iE6e0RbtMMB3cZqpxbtHeytkFPxY0dzne3
kUGBzbpDNktqDasaTQyVH8CXrTEr0+fRuZSVYYUEemSGAdDDZLMvPkZwDwbXxxCc
tOsOtK9Qo2OIuzgEqpWcaKqCWGDFtu5kOkpefvfycV5C5sdKZqDocR4yHs0pQNcN
zIAfU0t8g8e173nrSOQwU5IiDWILd9rnAzXTHw+h/ZlBAX4T0aDAgQPMcccSmzPX
nC1B/9F0f8NKU1kn/hwKvbN3qjZN9Umhbrkx6CSS5zYifakIdtWhoWpKBsDBTPHv
+wAi916M1fstTqqICeLZgF1ullSzeVYqdhAag5YpfF5EhNyRVskq5JgLyQ9V3GKy
xMQoAvyCWhAjVzfTzzyQl9jykmlfhkh5Zxkv5qizph5LQoIMO2TBbCuHFMgLoI5x
+SaSKMSsTaxEwE3q5F6S31w7tAcwgEHgmgEj82L4POfTt5G1yzl7BVt7lRJpDvLc
Cy9QLOX/pPlupcuHBYF2WFF6+3CcYaMl3+1Zn84S5/R9L8yMIaZnQtufTImDzuDx
YmDlogZrzdCe+ekYIcQc7Y7sI0ZzWADzTsbwhDoTxE5orgqr+yLpgokOHFBPH05j
41b0imjyXtojP74TCLydgUDyjtWZ+ZIb7kN2g/t/UNa4/mMNs3Ya2vO7d5e5Aiwi
9krBmUZ49g30OvB9Hb/l19srbAnct6NGDuHcXhUe6AtLoLlC4LuacAkfxmMt8zPP
Ue73CfFdoDwhIazyzowfJ79BYcwNSqKsViPMGUd1eVBc9DbmBHoNsZ5g/MJX2mlb
Bka7cCr0YrOVg21AdXOj9g3ZCDPCd+J6iTGV3WZbMNa86C9RtoLvsHNaNXn4OgX0
vY447Mrht2/zgzBjqJuqDMvYZdb1SeQu6+J2FrCOCn4Sw3XIVm0SivTH7O/2IhXl
5YzNl/9ezaNhpNx11++lcn9kk77cLsK9sRyQohbsD+IFjJlHI0knJT/eBI8Ugba+
1AyG1FTkEg2ZTKbkb1JMHpAK1vHDy68fIgi+cWX5UGki3UIVOKxdvAQU5xV55lsG
860HwSLjKp8vXYTiLzHUJxewSf6jY1lBI1SfmqpfD/zODlau+gepLvwCVIbrf6Bk
2fRzfMzWoLw2QywnQiPPIRdGDIMwRk78Kk0Wwxtgw7qDUOk2GJprch6FoOg6MJlA
KDuTONmPwSF18wN3UkqCoSpfiTZlYyjJUlKVQW+Rps1CzSourKjKbp2mZVy+fCxt
GtC1EGvcpOPFZ9XE6Q3/mphVLztjCpRcdYYuabhmdRFEMTGWWVrto5juFKswDnVM
/Z1aPGM6FvwhkzFtaL3ZH+srXYZHBDW0mFyo8mDfs1BRjKQ3LNAE4Tj7yqBI2tuL
onRMe2HEhINaoj6eVEndCwmayxQa3wmZUhDoROgTHFLEYMsufkarzziY0xo0j1Sv
g67YFfee+3j4jf2m4sCuQZl9xltpUpYBbT4U79R/8OnWtHmN4DimucgahE2ID580
7Tp1Q6nl9ihaMOtNZtTg3H487xnj15BmxWt7/wG0yQzLKAgR8YSJiQyrvATLyPLd
lvsUaYsJWfeRuD8CNyINiRVOWfXd2oUABiryBWEVdrUDmJJJzpUXKXs5UO86cfGm
UlDoU7MqGhpVF+K65uhakmAahQrkjaDbY3e7IiizQccfnz4HhyfQF8LrtaEY4IsX
ElHXhPo38D4Ys5RW4NFKm0MaMkQJzbGRbeMctFWzGa+2+01iE661blu8S1hX6YvU
54IKJLj6g+4XOQk9M0DvTzrp/9ycnAfTaLGz98zsGdUKTFsg2pcv+voiQdjWtypL
uvt0sQF7Xem0ETObQvFSH8WKrELa+Q+BBjmvuRe1W/xfWjn2ImWvhiVOZ2BCavz/
tw6A2pmZnCR0KjQ08Lc0CAyG3YrapWasFjttjxTQFOYvh1vxbgkxiJSG7XsV+HDi
OyvYmlSfSJU4K2jOqV7U8/ink9GKO+0oJHY7kepm/ZwaV2PhfJP2SYEVxcKewHp1
Yw67XMBO7Vy8eC1QBMjU7cBb99CmUDMqBm5keQk/s55Y32l0kMKd644J6vrjVVZM
4hUpxdd6KMSgsYZfaZ2oOVJZ3Odwu70efCkLzW25sALkv+tEvDhn8v9tQ9NTVFCX
Yh4wCXFgnong6PY5JffhxDhy1N00LiS3TzuDn28rz/W9aCnuF8qJd7EmfnDASn0V
HWtQvN2Ys5DArzl8siJUkbdbo851kxYhvhQ0w1gK6aX6ETmJ/bn9CDRfYMHqHd6Y
oIlA0RU5+IALW8K37b/dcSYEdtN0ftNXc3J2b5Co97NAX+FOYXHmm5/FzfX/oEPF
HM8WnSAvj1l2HLPC20zZvAl760HB27VvSUvVD+hUN+Dil3hoNt6AhxwWNyA6j2Hb
iJ5C2aWUH7M/eLcZBSUEf+0+0d3bNQJKa/dboS5JVyacsoIuGCrKmNBjAJwONckE
nhrNCP9BN3em/LyfLJlEFcT7QIlnzLaZ+TLmwfOF48RC6s8KSzRNJ1+xlmxLc4Bp
eOGq9mZGok3oBSFqaW8cqdLUqcwqm6k5x83NJu56IPQQ+pnDmR9ghDvFlYdQy0Sj
4VeXzQP0NRm61Ptia7WkUuTmMRCN4rkzdEyyW3rjQDav3vufSibQcvrc711DGxXB
1RyMv9iHZXSoubCu+FZt+0SSv5ZtzTOYSDW81SzLtt8CU+Cq1ysa4FO5PcG0UPiQ
vNFqifAvNBfr+i/4WCpjdxlTAA6y0jXKG0Yqq1x3KdAOq9NrIhPVjMW1XssTdCdG
tVCPVp/0ihmhJBAmb2tgta9MSiOJsVyESdmuj5IFXoLNz+1m96eBNKrallknf69E
yUWClj9ubbTQYg1WVNFaq+RNt7/vALtHGSeWNkEdiNemq/kz6cCWYBL+1smnTVuo
V/T1sbHBsOM3L1Z9piPPRJwjlhB+3H4XQiuQMMFdrWuDQdQofrTGbFvFlLo4lXpl
IzHPBushiG2PWUNKgQrz6Jk9Ku1Wm1VosOTiNray/3JVbRyKRUODUB1sz/GoFfL2
9/MHZzB/y5OclfHQthb6R9b2O07NvvBNhqIfueByGethnrbYZwGySu0LkQgd/Z3h
ho/JDHGz01dQh1LMlyTcOmleHES5rxJhgTRauAgOvJjjsnCDGbTgtKSSPtTx9+W6
/LU9QtmkeeBB5gJEsoX7fB/JVMXr2GkcODZwalAVWuRZXT0BdORSpDW4s4bx/Bgg
CdHT/vDbSd57ZdYvtlWlgZ8fbYRukeBGJNfg+C9phzB9wV5WPAAfitBMhZjDFFGY
2LscDQJJMCxZlUDBExrZ1OHNIhJQo0LxJo2ifYSiYry9SSVXK7SEgIgZT8/jC4I2
F83G0mUwFfjmAYaRIBPrpVadtbnOwcb4qdphLIJV3C84TDkQYdB5Sq4wYx95QTIC
slS5l+bzUWFdp6jCZ94m+GXAV77nCRjo0o4Xnc4zSOCy7f0M5Ka99q2QTeUAh/8m
VuooeohZVmD5FbnJK2qU+QF8wvnMVC+X36Wy591wygkGTSHZZL/ZzW0l+zgm0UNH
TMyo5732QAqo0CjWMEmHCzn56KkAZew1MoNy2vKSbOmQpIWxuNjO2wfKmQP5UDBv
YjOoUf2qrn5v8E+sIYroLdTIAViTbn8/RtJokJZSitnhVpJqW9kbq4ZTJLZKkor5
PPk1ZqzX4GRQbde8v/pdCXQx/NyTcY7a7h2P3bitaB9nHDLTF30evka5+VxGDTiN
Kj9UeUlPyJIl9a1nfW2Yr0ZODOOrOXH3JWbXREq8teR5S0pe+8sI/vuOY56/lROh
OGvCb8TiSXEgcY0MrerwXZE/8tN+XrZ7yFLDXLPf5JYH4Red3mYArfXmj8A2DU4C
39otv9UzU6E+bjSUbn9AaSj9ap+ZzDMWHunIJaI9xQzwpPdDfI4ur94klnc/rDC5
kx1FSJraJ4tqchJ97jqDh/L/896VirKhT1kKxpn031KKcmOm+/yqasdcAJyRskYb
u+iAuMkRPuU5KMcBlUJrsaBo+2f5MUlCiKXwqRlobV44eH1UkwsnlMFBDRmv4qye
ccabE2MzCRXyqh9SMLTJbeC2lOhfe827EaF4rtb/iDlSCG+1Wo8BrXUUf3Yuzymu
0iBXNTKIP1Z8KRtC5mhnzYILyuoSS9NsnEa6Ngch9zPxzl0a7GQEC6spFUI4jAVc
gT+UcbpCYcpGYg3skydFZdx4hhlcSNcclFTDgg6X+TOq23P7XsiHDZkaEHuiap18
La0ai18xMhK6ONC7iWDKfD9z/2ZQa6UXFLIZZY30TtkJKH8onNl00zdSA3HAKlpI
q3lYh6LudG4MFzF+326T3RA0r3de4j4kBjWwMyeYvX01z9QD3ffpAUspGM4ZLc7T
RdRKdpyuL8bR87lYaaP2m47nmU4OdESG8kT1NLDakFHpxWNwaK1naTilxPal28y8
3isLNdr3tdxVPsmpAZr/gQD3+MlCfQ/iX/jk5b1kx7zEGgM6Di8WijFtpDEF2sOr
0rWI8oVc5EV+7oSSdeRpwdvR84WPCkl6/Yuzg0kNMFCQZt0HcrExfyFwTSj3VCJY
syeLB5UKtipZ0+Aw7hjgk2DGiBF5/OGQGjcgAhp7qtSIKFQ4E5k2rhdaMKjlGrdz
uPnAfKZgEAmfD/V0OtjbiWrmJXCRV8RAEAR+dIkcApEwNhYeIRGrQaes7negYC+s
FV850TaGV8JQiaWbM95SevUkfWIqEJP6E9/BK6+CUIsBcxoM/RPlI0NngE8XbqDd
MyA5AHtPXTJU8ir2joEC//lYB9weNNQ+lx4eiHcTrm0d6Z8Y+MFiXcEPezkzFw2f
MxIbkK+q4o3xiUqqw5LTekadCQ7Z7jHsKr0hl/7OHRI7T6ZuIIrYfghdXGzG52Tc
ndvNBh6uY9/A69u1Tzfi4Zoa4pbJQnufJRb4llvmMunSxVooyj+uqjqcaly6PklW
B04hL4CaoCavtPuQ2lhb3CT02zu6DAjSjA/QG3jn1ZiuvZD00OVvT/iAzQ42BIhK
BpCeoScFYdqK1Y4onIeY2lUFc3c5ubICtlgm1Bz/71MVOnkEdWOmIDIKrAlo7ljc
opXNGS0lL7x3JDK80yPI8yov2Pto85QEY8oBZbeBg5/wkYCGuRtNbo3lpo/ONfMj
BKtNW0IbD/y/UPVSAlb4aMcWTufnTSzlay8ZKFdFg5eHuK1uI10KcdepHuvYuerS
XFaRScXPJ85xTlwd8B5zDsFMJwphifDJA7g5tWOVDIwpFFFEdBGBAWK09LurFP37
N9VnEqEBdfCd1Ot0inu7dUAxvlXbfBIcStQBKJ+sUESjpxmSg63WZY3TjTBr6lcu
7zVZ3uCCjifDQf0sktuZGacF5LEQYXXsyzbc2TWJj7jzr0L3Aswg8whwm9ldPmZh
JednA9IolKugbVFSbhNGlHAiDtQEbXBYpWPN9tk8N25Uql7FWWmJ8oZyyKYD7gK2
rdGPltL0dqx4re+KRBXZ96lJ6Ez8BtjDUQjChTxw3dwR5NL23geOCcjIA+CJOPnc
r0rVjAEXpKjpcb7K98U4aPEOF3qtf8A/q9uDbugVkl63VaDEQQvUQJT3lq7ej8qd
EUNhQ0R1aCcgH3BCrChEgb//AZe+QksQCWED5fNxZ0EauF88Dg4eJ6SQzrAVezLt
quEtQzJ0I1kiQZuGx2ajWdrQrgFALtBfDkmRPDThL5LTYIpPTFnrHNjJGKFRO6bT
geZUC0CPGoaCUEG/nbcHYr2s87oC7vxQ3EU0X79EGuxPHi9UDJY1Er5LQAIs3KhL
GBVs9w+Texs1uhQzb1W4Pw0leBJr6QQbiEZdAo3HDBUDNK0eCLGMzd5iKcFVvdAs
m9oVdEbFZZ79R8OYbgt6rAjTuJ9UFKNJGEKVxPPv6MQUIrxSrHJmkTfl2jBAEtX/
eYgmIc9aM3qdnQvvoU8gUX9rTAn0A80jt+Pmv4J4KClvxFTDLTiyYx/VSRKCisAZ
6gMTlWpS643jR1HWn47E7myPQX0BapIjO2xUI4Fmp/CwuS6sd+z5PTHN/n/TyPTV
gfLRmqWPq9a1j7gZK6GYVcKr+T321dbmwroOik5Oc9ZIbboUsGibJh40KqtoUiGN
wyA+R8k8zJ+YXcvIUQBvHgCchuexe9ROT07FhwghSEk5el7ER2F6tFCsVaBUCMbc
rJ5DRmg6jaoJfqVqkizIunrNa2nBLavJ8cBwBDoXO9UEuGCBzFvwxZy20TWQWRDP
D5VcT1uS663qxePTyuKduCx0bLWxLsaBt+zI/CKe/Fgc8HhWAHrAusgaQjt3XokO
lp5niZdOQM0t++IP2g+tO/Jf6x1nLL/xXerHDWjIN2g/wBtBsubzB4o/ysOT5Kh4
ob+I76eh7ZK/2hazESMs2v8/97fk1teaa9gbBagdLV6k+P0eFVpXf7Pfp11mYrUL
rYXVT5m2oft6jNU0C7s3UPHfNNbVjtJ8I5MU/PSM3GR55NXfNuNtGIfJEeZ2Q0VG
hZGNnDc0rJ6Ogtk83rh/ZbzwFzPNuQeB3HRNnBeb2mLUT5nxU3cOnY6lObm+pnZi
27fyBVVvh+tIPN8QJ6uxJCFerzGDkkmiyIhco6pIxRASZTHXgC5dWNfiMCPho/f/
NO54NKXHKU3+X+qUBY3bAplz/SY5DndE0GcQPe0xt2cSeMTyZaEU5h81/D0SLgSC
vHsJo7CQppCKRlu2V+fjNXnHWO3jp17fZtEmP/khdgJDZn6xFbDzZklTekCLO7L/
SiFJigSOQM/zqdXM7sTccJBlHsiGqHLebuP65U5jQX6QPsfyBrvx3ipdMQvtzM3L
/DjtvKEbiHqgb7xA2pZRfuo0Y8acO0AZwwLFURq87nlE0Sf8wAd2w67q35rRQULC
2AVarHiJpQ1/69zSdDxiCDnTHv6+/uV4OAu6xx6bP+I3xaxYwQ3m6MBf4F+I/bKX
EGGSpk9qY2Es9AzEsoYDe3zGez3N5tyIz9IWFhDTIN/lAQQ/fP3k6eaWGgbDLKMU
nwIWGi5pEtYwoEqRzoRH6c6gF9WCsaD5rKaKo8oymBSguDXJwdo8tEeoOLl5Q9Gu
1sBkZzbE4P4Sc/1fZf+wZTVP5hLXgNronmH3gPClUuoAomY8WOP44GKry4UtuXJo
zJuDwUURPr+IQl7LoVHQ2BLWuo3S3/4/wzqhgU/tDiC4rLfj+dgGD9CtRC7abKSy
kQFj8h4h+JC0sPipi5ffIgMrCvLUWJXpivpkKebzf80Ih3zdFdQQfqAjjbe4qFhu
ZjA6D3z/iqXT7ghUXTfVcn0L5Hln6CVhVTj/gVhqikBj0qm6i9ZijA5HBXeU8R9+
8xk781gv1eGIPPepvl2oV0+xOpg07cfMrF4djOcQ2pp5iodZFaRXspnVHlXKELTP
VbNzeaYSlII7aezDwyU9y4jbpBkhuQwkggovTnT64RTKGZYayv3yovxa3USZv6I+
LNNiV8VRZbpTeXcLjoeHcjZq2QQke56RzoQza9+A2RLMixPPUn+vFY9iYQh70zgQ
NuBg/yGsaK9VbUHwLDjDxPMc+kFKlaeCPrihAR/7GvVkJUlG63biKRYe/onzGlD+
7y/HYXZlAifcYTZ2DrrBivmUkSRaj1+P65p0Pp3ejhRucgXTAWT5J/iEZRLBdhAB
kY7YgGxH1iy8tcmE8bcpCNe/zOgLYDzzHXAwKTBCv1+VnExX51MVx9tr2IsspsFK
GWN0L60NBrr/BbBHqDfSiHDhAJGWrg8ffpnMvVW5bdfjsvyl/h8qIoy12rUh6EKd
GjbNSADOcUWv4NgNsVOpbZ3UzxrtPaZcmZOnXj+m0OMxGP0m16NRO8BtkgpowKsT
4pelJoAjjeW9xKGDddNxAJAeZs6V0nryGgvHm6dunQmfTDH/02jCx6X6J7pu0Oua
7yezuj8pIvMGCEU0wygSqerCInKWKfDq5WrvZh8v595yomiqLhfk7IAQbHFpYOQV
tX3FvKLmmOcEDw/ecyi2rGWgJg+6BWZcNv5WPNeLlkhwgYLgTZP37hKc5HMepYl7
9bVjzMAb029UKBw7nG1X3FzpkcuRQKrNKvsGBPRkv2Ct625QlxJrC/1vT86HEZio
C85CMqCp3BVVJnJu7FEbx1IXSTxdnssEJKwQY7MTVW1J8OU7rSFVUqKuZ7DwBoXP
19ziKkcw0eVXuBwh00RZfnv0RsbnHtK6Ig+lFACIMQ0ObBd9heJ3z+3dbzU9khYG
adoaBI1j49k4bWlanTu/7cbha3Rk6By2VOEz6FkudvPgOtgOJnfQN5MK1gWGRBxU
QC/kFQTQMXyoOSlwgF1UmaXT11ibrcZcun2ZCtKiED7kzY+QRuB0O8jUnA7mkDiY
xJ4lC/P7NT9AaQ7RGEMkp8lfSfLgb30oGNplEd8xfFDduLU8qNC/HR+gZs7CxNTf
qAAtI9bCEuA9qIegfI0L/QqYS50b1Xm7/KntzkP/qm+q3C7LjFCQx5V54TkOHDy6
Bt90LRlSZ3/8071vmJJXLO9Oq8/G9NZjHO9h+1tV/YUE5PuHSlrdSjkORI7PU40T
J7/R+hgYF4PaZGALAQBJtzWCT04/Akch2G4agtmhURYzowVq3Wcc3HPLTINFcEf7
bnl8A0eBMUwszjpmgCj2crFFAN7hk4KhV61pUbqrvb/M9Dp/BpqzvcKVCG/zi4V2
LPmWClngtWDT8Iba+JeR3UJ46aljKkbSpPzCTuNJOB4DOwpgwHKN/ctAtZMngj6/
vlQ+so/z4A+GN0JzIOHg/rOwwwu0hFOunnmffkRXspbzRzBGVscxtJQiyu2So5TB
KPbljgjQFGN6MRAUH7Ml5Lo1LOWVH6tkkoEW/bIVlkB5Z4rzjXRxByP6u145YpTu
TnyqCccquxpk59Gpzo+jBqGdOIbheTFOjL0v162raejcXhI9pYnkQv1PtHy7P3Gz
7R0Uam7gmVNAGLX7x57ywdYTSCO8x7XfdIVxLyHIZp/2rq3aIFE+cwMgCeWlglpN
BvNyFroBi211IjFobYiRzgrE0h+pIeeNhcbmm2JHXMtHO7ImVVFqDUGywM23uPXB
OjdI6CakNCZE87OLAModQfsoUK+/cw8LJ6j8q1eeb9ZGe9DZ04cZAM+njTxcSJpR
DYWSZ/J0huw/U1W8KOXUL3VJYimIKWZeWioFSlikINwISGnxSR+S5fZB7XI3Emi3
GaIh71uSYkpZFLrHz5ATCZiz7mIDhD0dtTRSPYU2Xn2cxo9Ir8dbjov7SAfAaSMC
sl9wxiOng7wn8nMraqdlThkrbMJzST9wvTJ0xcnEdH7QIPCtrf6Pceh0xzvxIIZE
5sBxb2adjKUq31/HKZnyxt+8+rS+J4JOqmuhXdFZbXvJgLUF9jx6ZhHk1R4iNF0Q
qlpSPT/Yl92nuUCNY4TAVPQze1CYtj7+c0aRn5gNncgq3hNjlrrfASzBD+6CKhZ6
83twtG4J5N2Z+iOuCBkvNDrPZTt36bZfd+aaVBRpIkkFKyB32Be/T2X7dU91f0NU
gz8rXQOGyZf6JG0A9NLqT2Ssv/Ou+c5f2ZmMGMPTz+913xW9fo0PDHG1lTg5tvnE
QHZmPyfClv6lmejj4J+I8Q7SUiJPwIUqM2OcZDhRmbFTn0xi98+30BeE7OvQ6i1C
cVJ2Iq/UqnR8+0CY/5vdM+DnS2jg83G+gBTbAUBRGWCyTZYl3OkPPYiL0y7KNvnt
viPfe1C21COYIaL1A9e+n926SESAVn4dw83IkUknLiSxPKYH43wHa5Iuax6MFNi8
zdwAuZg+5NyqCxizUmv2Ij0aCfNu7GBp0W4VD4g6QvM4uwnedoWzFykoVOOEn/pm
zH+3Tr3aKiEk/c/Bb1zoH0WrIISpWgfPWLVw/5QR7z1GlfazH5cATAm1IZzTjAyA
FMh87deO33fqqbJxPXIdZ8HWyDvObJI4fHqmF9d57RCJPmLoSEijIRDrZhG0AtPV
Fyz/xajI5rBz+cGNG33snah4V/2o97tTqELwOcIX7cbxWtPcb/jDuQACwByZLR1R
rdOfpOy3NN1FerP2vUh+gw//cliD21sodiKGDZgseovUGNW3zEN/4JvEKblbaZNI
yT9ZFdlANTr/zsCeWYkovqxHCyXZvfwDY3eAaeZ9UzbbDoWYoa+yhGFtForFlikX
VTu5pJfvSVyMc20IfMo93onGXgeRyLr1BbOBXv83GTmN+qEK6K1zHgHAiwK2xcOV
UOV2jHPGxUREuUSSAiQ40zxv73KPpfBWbDmlDNZDpryuqseQeugEDQBIHSpzqUXK
McHf6//0iJ0ZTTiHAy7McguHJVCCAMwimTy3eJAkGe8vS2j5jUpsJSMtVW6MmhZ4
Y0PeRsuEwvGflswXx0kGd4AQ5LJq+diXIDKntkmFDEWEY22oy9O3qvQOzFj1MIgO
H9CaUpxqMu8Oaom0GsYvGA9eWrAGnQeCbD/DN1QbL9B4AKzGusHL7SOA35fQmY1b
lmKH8eW+watFU19jWiUgvH1H/hLK5JdXBO03ooK1nNURmAVIkvhEEONqOvFn0xTL
mTEQ+E8fjaWQFYVU0QXQ6Fg3RaN5wez4ME9tOEJT22mSo5QWCTmdDoCvY9ukfnva
Fv9sPL+zTOoEMwfVjVynZSuNPpgg7CH+CbLLD4KpTya2zWSTcZ7KGu1vZ5K9Je8h
nioXK6z4TyF6pVq/pl4a4ix86SeSXs9Vwibv2CUrBdd41QHxdEwsn9fwapkMjyZU
MTyJEiDUwbVB9gelG6+DrNNv7tzjNlizJn+BfUdqxEoVU7GEcWlKta7jQVilN6+D
WuajgqSftt8ubXnsugf05ijzpBrboq/5LXDv8yKg5d61t4jZqhO/HA0EOVkbMYE1
T7dunvJmRVggVTQjlGid06YJ8TzRUToBlozlnqWLquZ6NXOxOWv4BlxMZeqOIt9x
CXg9LCJf/3CX8QQgDja7d171Vm+DNjdN0sqP4nrhBODRLXJrSY9z0iRQVqnFlP6h
wrN6zvkSJT7t1I8Ug354IGOQR326SYr7LX0VljE9sQYxz1QcqbhkWZ2MK843g5r/
UbYkUGGvubHh5I7NjKfBiGfkamsWIxOvKv0AVP9Pp0UDafAwQRi08wyFTKOZHgA4
i6LzjKDHS2jhtqA3ykoptitzPQaVsHfgJmTGti8OB5/Qlenz5XYJMWFBef26gEof
K3b2BUHGhrmI2SOy+VFxkUY/zfTe6KgQG+jw82zeOxjMgMPNqPZP/W/2F4VSazxu
gf4YBtO7gopClnx5VO6+Z/8PTklns/K2YWLJY8zouFAJ8uDwnLfH7IV/MwRt2Diu
d3OKp8s2I9IJC2g2Nt8+YgviZiwqxZy0LRBzkGgUAXsIo5Eektst1Huf5U7jW6pD
1YkiEPcIwjNA3zIPtvD5Z5E/X44QsNm9snKOEKCNhmbzboA/1MECBkVSEo3Q4rGW
c8jC5o7LZatBkWefeuFwE3WQHsoYZk70M5+dxf0ayqQRiJhFgWMjuqaoPErB8X/H
zYeVqnziRhGZx04pM/UvneUV6e7rSWZqNWI+ESXDutfdC6w4cB4XPg2trxFP56uZ
Q4qeLl11VK4fkC67s5Lz0VchWRENfXIDVwvo9O/pkfBr+P7AJKk5mFQUhy3k3KTd
ydJ/aV4t3IJCFCI8Gp17yZLWo0Cek4Sqa9vEneSrfh6MN6xObk96lYN0P/dn77fZ
YadyIvSYP6r+FyZxIIXABQYR5TKXY6wVngL3XhL3mV9BILSMgtm18Dy53v1I5HEz
StYpOE4Ibl3YnpRREszjLLktAnaxi0j02MuAFn9t9+WzlEhqoWLkvcQMxOfnRtQJ
H/DX/QXQNNzi+LHQTKAjsPbJ/yePKM0HDG2YtLFokBCVPayB7bwpGlvnHk5GAes+
C7/X+JuHp5KOJAEEYSWsHFVPSfKhAanq7U8KZqd0mFIm3Hs5rccdCxnmexmPcuQm
E6Nw8MSQ204Vjw9ovaPKYdzMKrEANlZfKr9M9rg36udSCROJzEUIv4u/WFC5TGoy
NxDXsN4RB6Ab/A5QnS64ErJrIhEzpHQUMNsCyH/+vhDNysQdv5+gkMYJPQW5BF74
dOZQvBwNVVU1XNymxW5BSe0BegsuQHOZCUVklZYIIGCy7gUftz7R4P61s87Kdmla
NNpR7C8jACwxcN0IB0bnFXrdVfpX2O3EjrBlfohZLLfBV4R+U9k2YLlhZLc9RBoL
BXpXETWzImjdqfeIbAxZuJ/m2ma+B+Pb8MvHEkqGMvRid40KwazPU7KNBvy1Jkbk
uoSMJ6OlLCro3V1JevlqKeK5gABThudoNmSHVUkW9jCm6vsy/InTfRenpqHGp4L5
PEew+a4Q7JO5V0+8Rrxtqhl1Zvzpmwdw4jQTUq/B1rMvCodUUrTOYIOHRsyZYNwn
DPULLAsf5h2w3d4pdcyFnzFglV9AyKrjVHrzX+UNIVc1qupHYIvI7SHC9aIdtQcC
kvh3KT0p2eaBizqjXIUMbLVAF5WGTdeHGkJiKKevbSG4KWHfpIY2zXF6QbAGAR0A
XMWGt1P3taQ8mt8S0CrnEEqlTDEx1Qlu1oN01PONnrLgBszEfdRVW5/r+sq33hfv
UrYAYGD+3Q+/psiOnp64YHQQfoeZauzW6vAOpIIbJCnaD/45n9tlqmYlSNJcBW5o
KspO6NPIOd6+agSXcnatnPJNNazXQAZlHPbbwxQP+LTWvYf9/14N22CEQjKcowX+
cBcgwx9SEaiMUzLpRCkF3lLNnDYJJmR9AzLt99ow4Lrss3SbzIlIsj+kDFgdWN/u
zshjbthPGlfbReLIs3zHPgUmmSnklrSrmxJA2TAo4gmkbUg+YflAWD7eUTnAvoBD
yQfXO3nhhZxR//bEUJAqsRxmJfHldB4Js57DsbSSbZxaOdi+TziQDXOhuABgltJa
/yXWgu0vcYmlRDmGt0iNZy0nDAlVMJTprTJQfAbDrqxPgXhuHY41VmYDa0Kn7Ljf
+g9fYV1mHYPgQeF/EqOYedtaBW7ws/Rw+dH+6/U04RiGCYRB/GLAa3P4Fo1YsaRu
nB0W103WUUuG0ZbHbjztoTd7z3NxxZL4tQCuGJdajikhS7r7y9mDm9ghgAkeRLbO
Sf0LmlUERwr6v7KWopWHjIGgVFhdFXYtzynkzAkZgEdE7GOle1ZRbZnQKIRET64C
SHH5rpnSf3QkrT2OMTwYRMb5QOT/yiE5x3ZMOiJVNk0+3Hs6Dqpm8yELR6PHN6Qu
66yK+jdesNFJa4FtUvIIIMm1UO8g7ALsCkxpuJhCcJ2VnRLlkXLdwwgx9iUC0VzS
QsVwNYGyT2LKSoWRpedcKhD6GIZm2pFNZsSe/ZF2hW52SzpGNZv/DigyJ2GdRlgp
3jKfWO4mpleK+BOaCeERV+/Cxgk5yY0IIXkrM1CtTT4xgghN7VX7kVaP41HfyCbg
6BHA3FIbv9sF6fFefTz0v/ecRf7SG49z+CrEp4YWempAv3Iot8E74v+6lePs+JiQ
TlvimCmCNs/TAw4v5HEktq6vxPvT9RfqfEST09hB1LGhJZyq6rMcFHoLwwRuNTxr
5kX9wmfNkmb5Io+A+LTtPVH086DNUFOPMZpW/pKScJi1YHGeRkcjafLUGEdVVQsh
2hQZIBChbVBga1LxXlXasewO4GTKcRZg59RjOXrxm0BzSCRz4hHIg9JF5TeAbnhL
8vGEpBj8+YpqyY8upqpBlcRkURjkCorH9QqA0Z/Q9aSunt8qD3/LfVHbDlJggNtT
416sxDbPq+IQ9/9fXct3BpGW9Nl4MwS6R63E72zdhQ++jW71pU970Ru3/8EtKk5b
P4ljiHzCGilGGutv3v2okocFTUO56sx+OJwc/8fQAmfXqMN38Dmnrmz9LarF3nO0
bs9T6HnWmyLDwsHIv7cauKp8De1WLLt2TVnYSFy2yJBEXb7m3iuxBAcMz+JMDPuw
UMO50B4xODkVYeBVKyqMpOhSWyG7nLDtH/6Jv7YrBRy1hgDNQVI4VjwUS/Fax96/
z8GFkvURgU0Vn7QGItsL27eTD+2K4oSZChNLmstHXxz2KhQ+wwx9XK/0BIFyJg/u
bpA08594PFwyAb2+eyac9U4KKlcLLx0q6lHQ/u53k8I+SfzwzesqDB+iSf13rvGx
xBBXsWizCLcysJuFUhcHZH8+7jjVcmjBvZJJnD7Y2C8F+kv6ejEXZcmgXxl5juJe
GA1BRQx0MPAankXGardinTeIhlz5/efNn0MA60Pv67Yvf8e0aUjfx+ohJgqhdKOJ
HCauTwZv8mxTSccFXYjmyW2uFkAh4IgTl/WgsC7aMMbsncq+ocJfWVZ9Fx0afTCe
1pTLyxUxSAdKJicXMTgp6MozooQno3l/2gl7L5iQCA1jeo9EbVEFYz0OZ/1qkdow
UIFF76AS0H3i89F7EV/coftR4NLrOHFs9RMIPCQGmYLH/GqbG15jFW695LGJOpLO
BFTGxBq/Ao1Il7//BtMbqz4rK2bz4xMskq8yNAGAeK8BYLDWbYyuHp2CAXmw3o+n
jIOL29vpSnT352jXyPXDOpeRJO2I0clR8JKlEVgOFlVYTYDKulsxu0WmkYSCYe15
EjQ2Cj2qlH/0RcOsLLQAeMT9VSBZhu3+JhP2JM1BPkkpj+QQqxOzWJF3jC+Tcko5
jTWkWB2hrroNLvka9uRcHinZnyUYFcPrv7WFulNJ4qOu2rrOu0XS/1FskQbzR5ji
EHVw8pD+KOMCvM98jx9qYbeBzNBFMU2IYLnnqx1cP+EdTZgqYYZvxWcu/7TlQtaK
5vL2m6lWp91xOOeU3sDnk1JzqkXQX6jCs0wrV/OpbfDefPLkhBxH31c0+vjf+W8Z
sNRY+/qSYHHU9rfaIaH59OSV+Be1z+6tzYb9icDJBE1puQagiagGQ7WR0GS1Yvb8
9z07Z7wIj/VahdQCYlzkLws7Admscdp+qbHS0ZVqJbFXPWhIK6NjEybY03Q76nX+
eqRTeT5qeNV8TsYlOP8+TDoQjW2zCKn1J/4rP6DHeTvE7DWeKarATcYiho2kA/nH
PtGubHVLccAMwEVn8Vj5Y+DMVSiAcAHbW/XJYfkZXFnDU9ltucRcC8JMXwCajT+T
zO2U5Lj0/yO5ISVDuSNRP/RHblTIvOuO1Jan+xX35YOq+Z19OKVVbi8Da5r0CS/0
1dqWB9rbGdhpSSBYDHUmTHxFV0YkzEDklGLSUT4FLRhHrBrwSnjqACz0Ygohlqhp
dA3bfXj+MWjVwJPkHqjDW8A7LTxS4ZNFfxH4xgcgoFrsmU2lX5jrPfiZFLXK/AHQ
lX+Ho+q4MqU3CiSs8BLxcX/dJYlgVdLLkx2g9GAive6tlk8zvYBVNVELeRBCWbjb
BFNGiy4c9CiMk3/MJpRTAaSnqT6qVI7yoRfUvnztYxb0TA50ZSUjogxPgv4aO+AN
NsXvagV4PuxKPEg/ztikRbmi/+CwZKXayD7sQnl37qLT7jRnWwK1BJ9RY3GWYdd6
OqSIhYpESSKxWlGDCV8Fx8Gx1E6tCEYmZo8B46u65NtrEvK9vYIU/nvYltvqGtpe
D6oHLZNOpr2nMKQFzwGYoci0STgjH+lIHAdMDMYQyJXcyuTjfTEwZ3Td24dWAqrO
luTNI5OEPqIc4h6a1Wu7famosaj8YeKDR8DMmzhclthNLABNNWrvCTdF4WFV9wm6
GjOWGU2VtuPSj2SHRBGN4NjQV+rRxq+GOqyIbg75YtdKhARqbwwCCMOn3ONYfHsM
BQ5QOzu5AGkiiwLDzVdCwVIs6SFBlKFN5FaeBZ3hLuEg+ekmsh87X53ArgihhDQU
qAbdqC968n4/L4Xgw3TuGXYJ+Ck7xKjGb0JW+GUNKgxd2a3SQpxlxW6f7lKZfOC5
0bJk8RjYVSvQPXCDsrLXhoi6uQv6eaIsn1otrvuYD9UK3sH0op5Mh6zHE6pArwHz
AGAm0KSAXyzbw++fkfuekk+tmeF+Qi+CDvJGJYZlLhN+OgNgcPjdOHfM5g0tnHjP
aZHZBtkPg/15DEs29g5M5wqQb8Qu4/LtGPPmb6rmZdCjFaWFBJvP1CAphWq8VG5h
SgucKiXhKdDpWqSoywiJBzBVww7ZJi9hQ7QQjlL4EBPnxnNRvHmQcpPC/uGw2CoE
GBNc0BEyCTcm3ht0cotCmFPMGc8rTcXrwPvc5JMs6VuAdgr3I58yRoXbWb5i4At7
WqYmjSHyTi94RFd0K1jw649iDg/AOP9El4p9yRKrjC82qU/zRKAmk1CdKLd6OPNH
AwPmOZkB0gxgCEN7SmEeBGG7PY0G9Mk/CNMQ6V6OKfzpGAGEtOiQL2V4gz/JDxi8
AVhlmAL0LcGVE35zogs4jduRIWwtnpOdq4o8OlxwBM9XV1IDiEewAuYa4/6m7LB0
QpLVEsjMJG/U9mcoDha7TSUQCU5vIynHeSt+ObrPGsbJP2lVYrv6Rvu7ZPxioG1y
SYdYPCqiaSojhuwkx0qMUeyxtKMh2hvku1DB1xH6dyfMfTTAnT2QDTzDS9OKkbMT
GJhT+Vroe/hEyBHkrN4xhxTp6XfIls/gpETMW6YK7D+kltXQhyBMQzVXv2vgwI0J
VmEjeljgwSQXO14Y5PUJofLo4j+5Ct4jw0wbxLTPs9Y6TLhDkjNfhtgLWiL6sSS+
AkloRI4Cg6E4D/xhK4IrZKW9dY8lwI75hdiWwYQt3OQpDhmOToaKl0s5EZS5Wcn1
SEVUHJmfp95KYfbJIssms3l2QxDqHHVOFdwJ8XLNr6kelIedDnipjzkhpIKvZ7sG
lGt4qKsB4g/hOveKPaQUttshm4qGhXHuhy9Wx2+gOxyDWgsMuimeX2sCiU2WwxbE
2os2K9bvCQocSbRFKp1WV1A8zbmQWvX3ssYUDG6eb6rt58UJixo0gcyAgTooVCFO
aM991YV2dmj3/pWhbo3ziEDbStDuDartD27y2oftrGRqWEKkCw3C+XTrbAwtBs4c
qzwo0eVQwcH8G1zk/MrK2wHAKN5gQCC7FdgtFbKo1xmWKSUp3CNnLQpPatmixLg/
1oJ8M8graTyYvWWqzfPd894v3J5+yjq09OFScRRoP0z/nBDgx07ra6QMXFGGYXBf
7ouwav+ejWzfykWgC6AB00O9bS9lbePXascVF6Il/mjQz9QbE/gMW7FvyTH6U76y
zuZYLQhc181ydmkSRbv+t74ARxx8jWLLuCSRKNpaKNX4Rj6JqcMlvE2XT8J59UcH
oZsJSi/PBgIqTti5X2bXoF9j7zqbp38Og+YdvoCuKQuRMEsg/XzRi2WdG0RkHVoy
L63zdfSNhstXEH2Yv2T3rXL/Q3lus7OCzXdeRbpamyYkQsskU+77gd9EdP8D57t2
2G8NgNW37c5rVSHDci4CiNrby6ujaMVRDo3kChVN17thZzjkVf0hOpp0UOdnJeBm
Kp1tp/hxcZK+6QUNpwTQZQz6yMv76k0Pi1BteFunugCV3nfsiArKh7NkLCZ9x6Q2
oJDUbkUX3nzbOtTORiMFJvF1S88QpvwUvHFWONFc0OvZg0F9BjYK1CqQbEyReVDK
Ds54NLWq5YfAsEstT+4XxNlZDcQ6c9M73sv+nxm+ztgfviEPX6D6BM41be+jcVAy
atOb9ElCu52HnhOyALYGl76Eit4tY/wGtjTB2R+TkrQNN6xqJf2WUCRf4FIj+MSA
7GEafQ80SpYClUFGm4oMU8O1v8f+NTJ+cDqtnTb2jkvoksn7Me42oeINK8sCZZdi
8E1FaLlCNskMw591HS5/xwo205zlHOIosIwnGBgbsRwTXLMXI5IyZSKy5oc2OUgi
sDUQjhFk3rohypRPm88c72ogIYoqhqz2gvpm9Tv6h3FXC+BsDI/rPZaaeCaYT/kG
CIHZhHupA4JufrnRtJQMtDYZZoH0VF2YX8beDpx1XKwzYEdWPWShzmJ1AD2svuws
vPeExRYMc3ge78Plo2j0GEv4xDh890Q+zqWoAC6Kptz1fNmZIwwMW50YeKHEH3EA
P9iJf91J0g9Kws1EPrh6GHzhn8WlSm8ZRZ88JFJBK8g9auOuyn9WfLecXReDf8Sx
Z4NkbWhhteQGs/KwTLxGtkkHr8jt+uAgV4OkNQqI9Oi8qmVV1e34ZNN2WoEhkr5x
lw9roxCgqn0a5SxK19uppYwjknDMlIOu2eDjP0EZE1QwPdvHxPAf1TUwu+IN/Dtq
VNRroBPQuQWj0BfgCrMbuPreDOluCOEylZFXR/bEl831F+U+zruXJNl7HQbg2sPd
CjHrcYS1ObYVIQDCOzmEGD2d6LVHl7/nRScYwDR8VHg5EiWmD4Spla6BjrFlwwA4
Rw/IfMsJdueVu1laM5dJ3SQgnj1JKGoUrH671qem7oqj0qPYkm71//stGBos/7Fd
ZCAB4aEjE3TFRbly9XI/L5lqxRBnUD97J/qJMYBZ2Xl936w1/+89BzQpkZDo3p5d
kDwMhtpSdXTNRuRaPaCPQFeM0mu2G8gw9FwAMnlq4d0SPlO9eeYWgQrJk27evnab
XHyg6IsfiVwKzyFGNyhaZP0TRgEV6yJG/j+V6ZJcKDg7wVMzAHvqU/zkN8lARbkI
4Sz62JUVUYZLDUqMRZXzeE+BvoGKQijRB7w1k7WCyKsHhUTMqx+oHvRl0ZYcJBmE
5eHdCDqxYxPDFJj5F5gHH2BXEag/Tdfbkze4SpsnNerzR1d8EzMdRhIzOQPzuQwY
Uvp+vKoWM6g7nyd8WvHYCrnwm5E6dE41pbwIzvyklugf4AemoGIPL6muLMtIdAP/
qR/Rj4V6yfbr3Wr7Vj6Nsqa8Wy7kdYHXooOVrOnMvxgyMLIIojCmyJj0FDJsGyYs
Kwmfick7BPGT3/wEBo9Hcx2wzDgECcr3tub2gFjJcfMQz0vMXOJKuXVdP9AVYyT7
bJ42bGG8dcU5xX8gchHVXz7cGp3KjKV7W402HB07e2PvZZIl2NoKOWnDNe3BPaEX
B71EsDrNb6SOlkjxHsZs9+MYkKaXnsIL7hCqBc10SmUePK0UyN8R7sjERiOsFn//
p0NlypHXHPAGyyHUqEH2MAFqx25aOJLsAgSv+8XNdwy/q4qJ6vF4MrF9DEefnkHp
XINis+P77/90c96mzCHBYhPXddlZR/YxF8FFaWfu9g16sSml2nzZ+LdnimDRU6lB
r43qs23ma52FqJB3c+ZZxg8rU4U+MZwXp8HdwQoIfpZK2GIEuepDD7u7v1JCUlWM
58Fa3lqllGxStZ1QyYQabkkHG8/ObpJZUFbgxNWsivektMB7HjROQMQSrwBlVbe/
YyYa1yVscw6OjN53EYJkZwa392XXsifI/gEEHFg6jNYm+vqtYzJdNTj0b+iaXJzg
sKo0XN5R5jLdpm+eTocRtCYxKyVZ5Y478SV6+UIjVyey4kw8yeyxuCmVUg/m3V61
4POE8c+4kg2PjOZavmLqMUtd/Zj5VHMDuIdwOZvW1psb0d3bpdAaSmjAB/g/uWIJ
PtXzWDyMKC49kRHVag0lehAMlYrFt5da4l5Tk+WUA+fxBRMab0MBhS0yGwnUy3eb
3UCnTS/otqdcocdiHDqei67znQEutwqP1pI3YEm2drJMgYkCrHba6FIQ0MgzDsWD
3Q2ZWiOf9fXIMvkSbNbDhXUhLQsAPEndCxIOJeKUzBKIueMOloNnKVmiE3iy99Ev
ARMwWUV3cJCA/mBxhZdu7NZGpA5DiHavrFs4aS76RkkOzH1AWVF1DRfUoBdYpMB8
hzIwP58oeyEZpEyVEVmIVkd3ZeBUBfrhOpZlZ18YD1tyr0e81d9LolTP8pvkRy96
RLgBsCzjzHDg44GnmivStK+MDec/0qtsMF6LdValhLY+tLj9S30Ahzq0b0XnWVvU
YuTRI0VvVWgGLsI9AsADRZstlRz/hBUb2HvXsZhSyOsvG8BodJi/QMPtqnyIMAdu
4WjzRDXAjvo539LVehAP6dtC4glm4K+yLm8TGg/6eZ1pJ2H+1oBjcwH/Dj7mCn3c
aIyAgyC5b7HyOgC5VWxQWK9hdIwu4Te0DmSt88bKhaoEwPRIJg5+XeuOuvimf1hC
FC/BBRLc0tglRXpKZOMDFNU30RZqasx8Lqv7nxiOHwDuyJJ0rnE/7XyFzfi1dz+c
h2lr3M3enAGFW2RLWRfN7vgs0p2Vd6zQlpCOUNOZJzscmwiT3EMjjOr38VJgatZh
UM2azZJeS9xe9TcJKT/1oxnuyKNIZjLYmHJHBS/8mP9PWgK5z/ULZJdkZiMJs5nA
l1c9qLkbcSWGAiKF+PcJJX/vJAetiR68DYt5+vYX6GF9nVIrAol0opAj3nnedkn6
QV3hticGegbj1pKr628AMPO81TezKzprLK/kDwi5A+NqLMQs7X0wtlTsXJq6IJz1
QaxC5bO8GAjwKy5vH4zzF0PhBb2gR5FtcPy2Nzx8QW4IfaFlYbaavwvvzg4Zgu5q
jUO9fZQjFhfuICKAlLWMh0lwtpku8K1beawFKjxcPGxRosvZQTlPw+bAu0ndp+66
zfx2ZmK/VnpNSlGKMLvc2ZHoGLLPJTWRYeYZX5Z3qfnjAlq0xS3uH3YS1sp/eMDM
S3phcYw+fYjRK57MfQ8Lstj93JENK7p81PkU8NKFOdz9EtmeZNET5uWGEdBy1hne
eRBwWWUMvn9fjKUjTdAF9zac7VHax4pClMyKEzaWxKpqWEqAzNg3YRUJXtc2RpXa
EIlXI6BdvFYPCckixHHaxJoGXmV0mYpUXtz7lQc9rPCEFPCKzFlIfHkUeovH8qvg
sPBKSMcM5e9xUvQ7x6jPEf43lvcIxJvfausyaLTE+KHsbRyt/GtY7gi95Ro17nkV
opB7ruMCPM/HIT+FohCpK7o8I7iekzf8M7Pz92KqeY9Tj8MDQ1Bdw8dw+eX7zyjX
4i6lRGKqaiz2FPVc+7FvN4JWIfPGjakGgLSZdNGsmexzLmojko7UoHVcyzMEXjLX
5MBNLELZrYVOR/eEazo6I/fp6qMuj2lVauTFBmPFNwznzJe90soKbXDdNqGYkJc4
UPFkrCCUqwvDNtCvfLMtpp65fhubbNIz1ljb3GLsdoW1bh7r+/0XLdKosshSmcBf
83k9LT57V90z/+npM4fR9XtlcRu04H7YqML/cVvF/C1tuALj34Tf7nfoPPyFJI2x
JgZVHblmO/pDYH2V+lyKOuhKQIGpWrn/WbbISUFPAxRGhC5XNSo0W6Karg1aMqS8
sJzhE2JL4e80MdYEXUKzCMsjMd9DHrdRE4JoIbuaQ336A5ww6FEAdPIazeX9cDiT
ChNCrvwIwdOja8uJIrft0lzo6enQNfm5Ve6E1oT8FHGmcWFRZLlL/2CI15+32yIJ
kFI8+hXfnEtwUF79jRmlJE6InYXAZJJSyZzeZfiaXiPl75uTmvsTfDNaPM5MKs9K
mcb+kYDOZqtBs24hmnLb/EWKiHa4AqdcwBsgqo1kvFc++J1fUWD8fE20d4S0JEI0
rLQ9I88+SeywH9M94qlExOANjJ+5xP4f/P/DehybrW3QMou30CZoGauqvm634sDw
esTNSyBII1nnzKdi5NB+baEYxXEklIxTiK/bFUvEqzrQV7ftr3oQYUfJnqB48IEC
FeTmdP12mIDPXFCQVREG2pfJrMx10lE500Ovcl0Hzvt5iDHFgW31EHrIRj62iOrq
YjBSYnzk7BdFLlR7dalnWCRJNaGFxEV6HdTNUqm/WVOCpBri4kuDclR3YFhAHpnP
GyMSt9A6bP69ZNXPahOvkjVdDbXJrV2/OFOB1VknLsEY/KI+x42+onoiSpuH8BlJ
DoupJAE1PHD9uvm9m4CSsHplx5VMh78+3ZEmv/N+EaIQ0LtvIuuc6jOvcOJWqc3o
6M0rP+x1FlcGfcULwxBQfEnZg+fxrDUM+UCYBptYpwN8kppIafydKoyB/hACYCBZ
z8VgUALB2jPJBSMn0HMW4hR8o8s+YEhB0/vbUcEJ+OCaa4x9z3z6gEoZZ4J0PMtX
9zxQqTUBnewPVBgwybDrHcKh70+EHv0RTLUdJtaebqU7AI3rs1651zDicthDHE/Z
UGfVuIeDMYPZIzbWNrj7LdbyYePrF3nLVQahwe5WtCKxPYDGOPloLxgQdaKF2IcH
IKU2U2vDNks/pbeGdnLnI5wAqxzlVVoFgddm6/8h06nAvNGaPrvwo8ULV+79SVI+
EIq/bH+7yFrMheeBCSc/L4cHXtTYLo2RzqyeJqNBVSyxPS0Uajg23btPrlWTPx4A
gcUBXqK3ibpCRt/H36Fx5HgPmd9/Ft3ujW0MUOrM3bhF5NKCyPQTiAgYvu3JCZS6
UGDuTR1S26Z6R4dnHMb162tZT1WcYtqH5g3RW7qNS6MQYHQ5w5yrPOQgKq/1PfaO
ky+cHOz75ujRvPacHHEfijETrpw2vt/tXdVLIP9LcoGZUgi0PYc2dFYjc5Qs9gNZ
jX469CRbPfPGCb9nSC1wLm3Mwh64TLp63sq00fiHRq7721mEsaVC6ruuDoPC1YUZ
QKAxqW1443ypzPUwgHhrh+m1V5D0ZFXozvRPNuCo4B+JMK2fa7dSBY4NsIelv5dr
3HEFfqQKvMp0j4BdezFI0x9/f8nQKoiuESqI3wAK4OjA46j0J3VfISTjzoTl6rq6
2WW3uyk7T5hhIbp5UzctpO4BnDONmsLEVzHlatniNrsFt2BAZceo00RJ5owGuT4G
pIho5ANjMOLeza1Ugt0sgahznFdLmkNN0U0P1Q4Pg9ssnVgJkimrZGBgO6/m6WE2
Q9gV9ntXJO1ypWbQMHcroKuz83LqFNewVOI8ixzYDFnM+ElQE3gZ5S6GPg4LmfP0
zYu507mxXgxtG9GKog2MTSxfcKWe9zlkaDKQ9L2/qQqsBzCrWTbwSF7qF5Lm5Ri4
zx5fmA29MQ1Es+WV0bh+S+jaSlsYzqTGPhtPXYWYpBFj7SAtFnlk4OQhAzjIWAac
uIH/XQ7upPkS3MPWtggR/SgIELcBe7kql3UZqv77NVpPCODXmEbL+7a22/zWusI4
+Gn4T6zGjMwzvnSLtjvS6Bis1FLKvAZwyDY5n9/D/H7xBFO7S+7EsTUinylto+FV
xjmE9mZG5YLky0JbnOK60N/Hb5Xcvymm+u0M9GmjQUOX2sgpL9CzOlKVYFhpNteU
R3PzPs0MyD/+v17Qw4t4UYMjrXujIFphPYUF77q123i/B6FQyP3dkgf8xmTWAc4V
rUXC9WXeCnJk5nv1NL5+SalGXqF6+oM6vZgpqctpsH6Ze6+U3sWNQc8EODJjhluf
CT+jgJm6wO4mjLsW6AhKjRRZAahGVvBe3PFO8D7Zq7tVk8sV76oiDaUXTaeAySeY
2Eu1m2GGGX11lma4aZ8IUr0zk2ihVwJV4eU6ebUB/6NzvX5PI8RKCyeI6Fruvwmc
FRUqqHNsJSPjEC0Ue0sJSGFGD4lh0quoq+xVKpvV2Bx2+J7N1BEGYTZ5mX+FaoHo
Ex7PSNebesrNG4VyqKX0721x1/MwtLLtmiAALYXg8wDdeAg+xeP2ZwCA9EO9H8uZ
WBDZmJEVUeE942vf+Gztjm6UBdpXRgfy9VS5ClJ347H0iyhlNzRRK0di0KEdC+ob
cfIBhmEYBanPvI3luRAd+M0+qMFL2xN2LP9MwBkPGUuHjm2yFxFhzzhniOKRxAlz
jqPhINLAFmPonGikXThcdBbIcPaeadP9S+p5NNlwFL7q48hikwERDoFdBV2HBsFT
ugQiQTlh3EttqthEC9QgEogtsqk4QPRMn9pilsm4ob1MePWc6OSg7cDilWWYYI+M
5qTPu1UVBTYVbTpNvmJs4itYxiw6yl+RkNkpfPQ08mlZYlueiDEpIlXQtNfquXJj
7Ya/bPqTxOOc+NRf6WjikedoD4j0PNC7pIRJJThNHS4F6TEzWEIRbI5c7F8A8j4l
XWumo5DczPm2iCVwrDERd8pO0mwmFp5ECcNUovIuu5Z5OwwlZWUGymbnegn1xcc+
mRkAO841cH3jHjop/bSDU8UbNcPrP+JTJd2OSF4Edm3kjtMuWRsmTMbZWXCfdLpk
YGzPRpIvo9hYHQbnvjlqH5m5/2mny3fq2CKJyoE+seFyd5riPLSNSVeGCgAEknSH
y7WdvdCzmiMGCKKpEgkcT96F3gGPicEmJ2fixbKm8iDWFg3ob2EGrXzhSke71XhT
/LQVPmd9vmYP/VGJPreU5erlFe8Oy85Tuubtk52YCKsaTlHHXnN/tXn2d4amAbtF
Idmd+lTcBBgCRfhHsCwz1Lrjzv3T8m1umYGXicJSwWPbC2z9LD4wEe7ESbiYeYzs
rAJHX0gtTCUeVOykmmlZOFlPZngpBTwTftFXlsCfBFaoUfWvZQHJH0L9vgsmqgvi
X4qnsiTTyFJvCYhAYIj+f3UOCyDE9UKXYI0ql1De1zZrNWRlcHS8LQKfTL8XGTxl
dAgFChV0y+exqLtUoWPTog5803Bi/SyiwnWAkXH2w0V5FMyxYeYF3TG8OBbrjuoY
168BaJbz3LCo1UltKXCcTcYUsbfELX3xtG6yoB2Bp4aU5sH/g4Bj9BieTksAMYv+
91h15Udl5LcIj44LloGxu4pbSuzsagEEMLXoMOlijkOxXI5semzyujvyn9zMTAUP
hRNEQQ1ve9DzWDY2T1UbVYDz7AHv0CLPO9bstHZjf994IJQAJL0MIXf6qUHmjBCX
vNrzSvGcS2DFCCarQ3BHeW6OQbI7UKqq4JtDTnqAs7wbd9gXj1fy4HSSKFCx1OP+
pSwv8UB8J3sXBD1bR9GLn5fV7Mv0gxZU/v/CP6ZJJ6e49Rs/EeJQORf4yLGTArgY
wNZvpFfDoZ/AQo2QAJqQrrX+aYqqXE4cHAxGz5VUU55sUTalxZ5ur5cw9Ekn1C9T
XEQYa/ycOwGyBYWDAnlW2OCt0vbP5gb5cNxkxRC8wpjWSV3apwVVdZRZ78/nfphS
kJWEktLTQqUribhs0OJmngD1i7c8KHegZt5rxgN1JnKtlymJ1nXwjvrT6d7NKvIX
2lEHI5YHPjdT9G+dcQbhs+EYz11cQBoZrSvDmlnF3acEkqy81oFZSZ/c/n0Wg6kU
G9TTgdaGwf6zF40zE3bm0ggf9SwaBeAaQ5l2cxdIUNZIFtKoRJYMrEU0LoON7Fry
bZ54SXUgxRImM6eK2zQF5oIMDQ4D79x0Hnn8Laz50G4TCczXm9L/jrpWIO62C1g2
kmHVOIE/7kUnNLsc9Vya+nLwKfGvpIaSWwr+KvvW7N4SFvjea4p7KsEZlHr4Gbrk
sVt1q9Csowxoz0Wu6bZdkBcjygHHqehjF7c9yb7gdztkO1iPIUkVD5SIByme+eFF
yEn5juPfRX0rDteylreu5D4jAgb257BS0TylKKSJQ4sVKAbRnkk8h3BjmsmKAQGH
3fOCPzU3FJdy1QVkUcD6wOlevi6RszsEPbj9k0iM33IPiMaQImGJURAzf2Y8ogqJ
h2f4gHCXkwWEOQvE0eV9NGj1YXumoaC+S+IcjEkoC4ygi3vSocqZxJpKAOL5RXLd
LXkIp2I5Hi51VOVpJaG1YKqYsaX185MZKiRMo94syA/RBjMYM1R6Y9nTwUhReA5d
g1L8ZVzY2ib0/+Gx3hrGeRuRHF0epTN6FN6AzccnY8Yvju2R0kANaZ3c/0C0yYPO
CBgD+r/bLsS/XVKMrU4kMiOJLs5/ROgYIK95gSI6ai8s53PrDCkF5qCO68KdsCha
/h5IgZMTxrS/LgBvbS5BHknTjXBFQJs/K5dJWrK4c1MSKQshbVqqA3rt5XfLYXjO
zeviz+1uFeWkiD4/g70A53yExt1nN53jxuiMJ4NrZ+ttuEHg+lc9Oj1wAlLKvigW
RyVW4vK2DYoZBHmLc9jtpFnrkynxuMBQU72nzuOso9r86h24EiFqYS79I4T+C0zN
2p4atOMXRlcwGjjl2mXLst8JT77C+To1+JjfoQGQg7HmtAwuyVgTziaZTzvFgr+z
PJBUIeSD+HbmYglaGw/ArYcnCbHOdTL1SOCWpLpEYJziMZf1tEL5G4hMagjj8HSE
gaJIEP7i08DeE16XRusISYH+tFFIt/vOhFclTMF2uqoZJiurcDc2thvBaOq0wFY+
sBED1TLV6IPiJhGjH82c0RN4gT7tscCwrKdwFUyS8TU2e5yBID0LeSstXXwUlXts
Wi1pakaWMy2tZ22NMv7HsGzguBQWlQxUcMK3wjzN/XlwKtnhfbJtSp4TAnWIcg71
JbjNVClTxI99w6CAOX9qyTmAR71jl+STs9JFfw5tVeJNEBFZ3kd/3i3XXR1yFUZm
EIEAbu4Wj9DjE67Rbj9fUVqmWPkeq4479XXlcivay93Xn4vl2qSa7zVxUyS2yBNJ
w6cshxnMSkME0rvLk/4FQAH5AG9UksOAS53N0TItcZTsjEroVieVMPDeIKU03cGq
jiBLNMf9R1yWWbDWHi005ahIZM6RwrSfRrdEEO1K87BNtO2Qae94mtnEK0Jba6tu
FuSh0oiiABmGSmv4goPZ91180Yg0eipau/XsZMGcpUsb3Ur2mlX7zrTAuxXbkQ+p
GX8jjPQb7zHpi9AZbaehUVKUM3NcFjBZ6WztCWklI7xYOpqjdpaDnVHgvtpPUcFr
qtxP3CPS8Ot794qn+yzW9wPyuHG5xKAVn5Hmnb15Ev8ugWpYRgZPOy2ew3HBYe7a
TS+sC0jhz9OGZvjdXbO8/09T9uhhqG/gJIXpjAUltENDSjCXPhfTyWxOAT0rweIU
F1yBcnu+UJ+iqTyL7rYindfUv/LtS04jiEHIu0rA+L4O3xsEJFVat8bdrC8MIZAg
y+97ffZTtYLiddqGZN9us0nVy340q/OWgasFMqRWsG+44QCMURJEm6OpM+WNBsys
3etlANnzDphMx9mLIQPrdD/c3GuWxIcESn4rlw9Rqi5grG8r+iXBLW+eUhEwg14W
g+9tY5dq+hahcPehdZ3Nim8Z8aogpoHEluCIJPR2EO/xzSJ8Qoesp/B2Nb8ZLESN
B9i0FGVsziw8mHVKwVD93v7dtqaVxr8f9AvPYwURQz7jSPWYty1hqB41PqYsstAs
BS8stMupLb6Xr+wbim/GduL3OlSnfRLDULW6FGXaJRx2YiIt5A77ZDp6gNlFWUaX
EIMgTFZNmO8GCnfQADhK4TwwwELEUt21/t7xYz+qtY3SeFBf79pCuMKM2acMiERi
40FCHJQoRsfbxQscUgdUOCqvofvtvF6imygEmhhB2B6v1duepwydBFDacjBFZiPX
T5IBVfP7FfWER2T0uPCCdra3R7xJ4GYKTQbiB8pj6sUvaqIDAtnmEIUPvdT3fcQP
2Z6Bv6I/evzVmXUxYUvbJmuIb3L6SkKaRAtRE4c6FxPoI/m/1Nmfb9uu4BJPIivM
UD/gNXvY53LnYIg5VnL+EvqZnoveC8QBlTMzmjJ2JDFLDVEUT4gooOLN67UUu6tz
aDpmnnudKxh92IlKxWbyv+ypr+nEIZZYQ+AX2Wlbuy/vy3eHn7ViZMobHQCP2Ef1
yhCn31lz3Hsf4jtycd+M2XR6vHQuyNQ3B63h5WLvzq+Cjd8Pg/yya8k2pTsMJMfK
UiysEeSwzxgPmkXVZSlx7SThi3sCjJfHw+wirwEnGsaHH3FeV0ti0enr3kQb05mA
0AEDdXx71ALzc9EZYp/1LGFRzvq5Br4qeFgYwhJQJY5zkOOXtPmzko8YXVK0ZvHH
7T3xNwyG71TEGnvqidpCHbjGpE0/XEntcDmBRfEhUm5NPktVMdDWCxGUGLFffk35
xE6D1ZNFYum1AY2AZ8yqjl7wgFl8LaRp4i1f7Q2dm+OgJJEOd6VTjUMgPZp0MgtK
KV1ExaYQ4aMk5cEU3nTdTPd1dubNFc+O5nYFPdIVUFCPfV6RuzXmQjaDujpn5SZq
W1WtTZ7Y4ZrWC9ovOv+ubAZ27P9rvrzHxu3V/ngo9dI6UZNJjhyfYIrCXpM3viA8
sdtjg3mT5KCmeTgwMq11Tm1CK4c5c6CNt3ncGrlm8VSTV84U8BpOAYDrNTgXuOJY
E8/tv0U632a/rs/UAAqD2jmDpyPM+UvDwnXmjBTQAyX7aHqkkg5b+41jvk+0Snwi
LbA61jdD9pJ7hZt3y3HucNB1Gt6y7zVttSrwhoRtT2mt9cDIyxkLCqhsQl+cBgmM
3hZjOOMMgGMag/1sdZHq8GmC1yxA9+zLcVQPSUYa9+vzJPF1WIV21vhJBhSE9LO2
qM0TRaGSfugMmuSAmLiBr3ISO4GhShBrRcLbzRfBoFxx8n8wjJxopBXUpL1Urbrl
Ha1e2Y+uYBpqYKzzjFeNaYl/lpdJ6sIoo0KQ6nlY3GFl4zHdTqYj/Vd9wTeipuMk
RRFwaKaOsriNicm/9WayGOH2xjfjiaURrXee8HdRElSM6ULrhxdr4R552OoW9+Ry
EysHBT+x3OPcWn1jEMfLvaf/+I9Qb4pBG1nxiMnykfsyGZSueSta2BmdS44yp96Q
E6nuGlT1PrSiNynhIKwcjiEGkuRlyacyGQdbyPrQUC5cUqGiwL4MbjaETyAuRZAW
YsHSXUcynj08LgK00ZM1S147REg6IAKhjAqcbFzPW1tApxzKyRKbI2eu6F1d5Zd1
2JoGxIqEpeMzmanUDUJeGyrCOuyE7DBu2hWfE4H08UIJiwk5S1XOZYQkKO2B38Z/
AyMYM8NBFljSX34BsgEQiTBF5GdXkxc+4oYH5Nj7uvS1esLBnyb9zO7Kn1pt3l9M
JA7hIHCmVXxG05cj7nBEh5jhwkiji+PFpFoPiZWDn1gmwFLWewvYGWjvfSD00FsC
ySO3wkAGcPWDGhJOmlQjcRlf6H6uFSwL3ERZAzD9rKpXFtNHWd+2HAJb7V0vOBc+
GZ/C+5HkJ1qL8M2Qza/uwmeMkBPssqGKx9c7g3BM4RWSKn87lsTeQk+gaYxER5eJ
h64nh+RHut6yAYV6Ixa+2E30hTrwfo4+m3/iaGsIscqET8bF+sNjjB7t5s+jjtzk
xBRGkfDneRDFKTYU39NLjxpDBNW5mxFT3lmbUqJPv2YnznEpAyvPxw0iNCMGQRGP
Kw4TvAXG2IL3NfRPxPJoo8A0rGiRzwNpWGlpk9cBj38mHtkyQyBXX0G8k7E664r1
6B5feUCLccYUGuJmc/1lm5sWsWjdgOud+Nf9PXpehby6Xv0q45tlXKRKJ7ZvvjM2
dZ7XTFFV+0GiwpyzmxSBYpOuMxMs8U6gOB46n8K+mP5NpfzYSLInSFEi9zhnYuPv
DU/caHSK8p+HvXUvVJ8Wj4S/jmLUM41xVQ//RaBCfoju+yw34t1EZTXsVUGNDxF0
peov6GgkEYd0IgVB48kE7BZ1DxfwA9hAh0WQoLIsTxIuGgQd0dkZyxf9DDl3vHmz
YsdpNlcJecGnzFbfWQIftX7gR4XISsSepFmULEXDkRGAs0xUMlVzky6uW1HPExWl
ggvkCqqZw+GLKuXs/qF0QLEelvBWiGoHsLqXQxNEvSRQ5JsBPi4KZyOO3r5cCvMJ
ydiF57YtcU+Vq8NtAPMBiYsUtGwHICnu1g9iI64/v+yUMXEiFk69zdWrPptOhaAl
tuCrNzVJCj29d1KTYr16md7ettqVEn2YeM63LBjn9OGpFlDLh+aNjNjxpHgebXro
P59bkVs2Je61tc5ZaEGgNJx5rt3pZ1jQvH8vhgwWd6NgLTkXO4kUYSoSqVbFPEB6
2iYMd8gdNqafdmdeLsgAhOHbJ+f9INQgCmLo4deTuR8Uusv+VqXDRJODAkvg47zu
9Q+eTfiK+2wFWmJ3lyZQtDZqHkNLhdPyg7SudWOW3Cb+smwBZC30Amxf6jby9mLs
qHunC3UrOKLWxfUKwqxmSqaceOHnzQv+7VwVC6CrvqLxGLi9YTSGMZmn8ubBLpYF
26fcSUEPtzYaYO3/XOqSu4lygmDguNdMl/kSPfYis4DLgqd+V5yKVq2A3iywMfig
yzg2ey4K2ZH6WmxQ5M+18gpIziNjWIctGHTw+GTO4E+6KeyuWpeDbwvKF4D5Irfu
7LvQ+BA5zZPmNK3ojqUlYctsZSTgOWBrqB4L1X3feIzTUywWwYS+6hQalLBpfC6a
KOHM7qSn8v0kUFmm6cp+rea0PuDbviwMOsvtgfuSIA0mSlTQs7Ltp3cztXWTS2HL
VdYxzx0O5vKz+w710WWUlHuAZRSlceuhCh+mCH8ASIYBTyujVpj6Sc9cYl3eAEwT
EnlvJhs+TNb59eHBI1GPpdzarzLkYfWEF56R3yqR7hXu1kgJ/8iKH+r0HnKYeRd7
HuZVIA3Bmndz8UMdKtqvqeygI+ixFXU4/HA4118ECxVK9YJWFLFTNiiNdApnu1f3
gdlqCHEAHE0GBg0J+WRnzjbzGq/Kw2n80qFcVlE1u0YBBpifupRWJaRNbU27Mz4D
xAS37IIn8ftGS3XjAgVpVPHOgvo2XBJ8nhj4MIi/cfQyVehacMdZOhMGhwN/4Kp4
sgiFWNg1r7yFAwkhvNIj5E6IThSV/Ea9Krq4g8IlmCXrKGGT4EosXLXTMbeoo5eq
pp9HkPil95Px7M4ZyxAN7l4dGRmb+iV6lYlx71lZGBJayKxJoVyfyS3ukWJZyHMQ
1HGybkY7hcEUEOt+N3dry9l8rqwd0089AkBkUidjwx/JUm4foBeeSTUg5CQCmViq
IAblmJ0Eyz/CgkxdiqRu8sNliVfkzaemqgc8dXlOl33e+ae2I7qRl/Ol9+JTPR+8
9CsAdzNhNp1c9bsb//ogAQgUzfCmaz6ncDWRpJZ971GXx9h5yTzfvBkKOHI4nXUt
XQcYJKYgq28qUN7sLoVj8ZRdmFzh8U2ODY8F/PkOUThXVnQpJzlo59AYu7lqYKNk
G8uOqDNsT2JUWlvaXki2RINlqzBYvV/1pL/sctLEIC1osS9n9SOkua4JOSpXnEbr
ajl/WdZBS3fuZc1VzrFdEWZ9qQ+l0GiDAMd+y4JWtByHT+tiJCXbEe86yJpVZDwv
3La1gDhWXw9vTTAvgQVz3Q6ERJTR/Q+U5oIXIUMLgWOi8FtuCe+EZnrgR2Bkj33S
uaqn9h+u4MrOZMCdRGhtUTgNAgU23XQ070IkRzo8x1yg4iwj9gP8jMp+38swc9xq
frWWST5k4zOfvYOzd4L0chT3FTxxF20cWi+5US3SFklXlMvm12dUsQREIwuug7XN
q2h65w6dPDQc8U5u26dkQYFdldvM81yii/cacvWgw3oorOLM98RIr90vi8vPc6b4
3aMSYlry4PGJivCTZ3yjQwDv1M4OpWrSHGbAYcITDWtqMb+jKhQBfPREFkbj0y3m
qQeRaDtaTHT8JcAxpCkb0O4tu3sZql8D64HVefIKM1e7s1POUJshxWN/85a2KnSP
IBGLGpNMWkD/SAVq7YgNlM5hElodTtzpY+Nbt56X7IWTU8p+qSFA272SGw134pdg
h0TyODZgpXYfwT1ipi9dGgSF5eWbjcaGWoIBsEwVRSS7zBuArNlfQXyCJ2HWi79I
RaS5bKDJRj1CypGuvDAWwF8dQyhNXfuuTIMl7sxX29lKSCE77BmcJbPOYjzfhTxe
7X/3Nyl0m590bVvLAG35Icmc7DuyFUNrW+CBvqA9Ck0dMVngY3qcRoWIElzrGX6R
cUYJZK+poCfORXvYzhWowV0/X5XRJdKF9C4fB6/sv+Gn36qjSnJC+mumHml2xeFX
3jPs+ZaR7a9S1eGP7Gyohc8vVN8asSBoASft6zl72Rj1l8bZpwEc4d3tbzmIifOz
KYJwbbkHT9UuvI/F2e58myoH9MDpXC2+ApbHWxGKEEgiBOf972eTv+AJkAkIGUPY
8FAgbJmRwV4eM/pjyjr1isWQjLgaDjzxtVf2UBtfFtEBa8em09ilmVcVwbfNT9M8
EsNXyuXofynuepnbuFNXo9jQyV6zsn7HKPpWK+9dUfQzyfs5a728rYMuiHeBtHWP
xm9uVs9+oXm5+NK4aWee9reCO7oifmO8s2vwnwxQ0ZLYqknfyOcEbNpylschrasB
PZHicuU+CBDGUtEPQ2Z9v/M7Co7J0lBPhKfRyYiObU6XKaHtOrQDhVDyON9EB4KB
nMXmaGc2c+V98YnGi84joVb5n/+zovyT3XUraKHjITRPzwdPC+1+qWWCpVTGfbzo
fCduoMvuoFPRc8UWyvz0XO4w88F2KmPhDAjdCB9iZ0MIG6+lC69nFhr9f9iLS9n5
VnmzEKY7zcFP9yT2jVQJTsBs5pKzAFhvNUX9HPUJXitzYAMjJaosiHPUixV0NLGP
ALtChEeft2fMZvHS6P0jcjd2cOnCjzLsZ/0seSUVySPLo0ncAGBr+TtY7ZB2gdEC
U82pDpHlvPcLuejKoId+4aEWDLzZ0osQ4rY8r3HVf+QhGPpl610MF0Sn731hipx1
HLf/vBopPATX/o/9TpJP+DC/mNKUAtNBd+po/QEFo8LGHPAXyq2vXVz2qy+s2Jao
KJ5s359qSpcVw1cUEsIUoVdXAZqieaw7IuZkTG+y9yUTWpGh2zOBcAOxFSS6bk6x
BKXK3uQSYyWsmRfi0MJHlj8QU9CjZOknRp+CTHPB5Q3yo3rEiwTw6V/IyBzAqBJK
LLG3+qETAvp7aZm/3ZUdcyu6oMLmNMp8vi+dRM6twaLjPQfOuOsmF6oxooqRRJ7u
DEBPL/bH1VO17hjYM+u9KKYxKE0yCdd/0VXG7iZP0zHk5VY1VSByXjBXtkpvrASo
Um9SoR2hpF6YV0Nh4/lqtgjDcyeUG/F4iUg99qKv3S4GdRrvKz/btUChEao8f3FQ
O5hE3b9AXU3NSTbAQImBsxMuWwxvTUXkWSMx61e5MMdGEEzc/50hunHrar65jeNv
ni9CYy9M0CRLhBSMm+AEYfeSTwcTbYKYVP+6+ZJ1T4FEGp/jyuqxBy863BKT8KlT
PkcZNjE4y1hmdGfEiVzjvrt/MwcbEMpukp2TmsHfuOnafyrprZCtEVEHDLMH14QX
G2dRyRIAWxFTDD0EeZWhfP6iaeQfPeIkvPe/0rjk1VNfW0KFmJSbfgXEVt0Zys2B
Pq3TPMnF5EAuipdi3ZlGL410XgQ+nR1xeinOsFywsF8Q6fviYzOO2Qx6ond9XTyG
PWq3d/ULv/Pot+Af4WREG4t/eQ8CaoVIsiMGjAVUoW/JhhidrOnVAg+K5i0jyDhu
JgBx0TrsTKw2iYXSecbyuVyOxCu7yNqCDe3niuFSCaog3IwKD85BNLYUoKop0Vyf
Zg/g5IF0Cu9JlbA2GZ+8qP1pi+Fw6CV0YXopfwOyvwzkLW+XfvEiNPROtaLFEK75
wL6eCa7dA2wFltcXnbvU8ioGbxA12bzZfM7lzxzEyPXqelg+RnFjBTLLXOVJOViz
luzprwM+ugQmDLkOcaicqFiFGpOvF9nFNbSFxb3Is5WNLtQYYRn9e3A8/GZIuQEA
LCV8bL5rKrit+W+YDbDxBgFw4yFlDkYrfWmCHUUrG+yTTs/4dMHhHDGrQ9QrLnK4
aLHN6lPdlBekiez42CIiRYMrDue+ye06vdJmA9QgxOejAl04uAp1JOscexgrN8us
EVK0w8iHalxbMQSYxps3o1IDjIouOYQDVcsVTzIODlw8MhLnXc1S0jmHRd0WaHCx
TNb2TgpSUuKn66X+LfEygt2APqJdZ+Z2GjwpiKFGTtCiAPFgDhXSVEelTbLFHRr2
kxOQtIlpNdRQ3VcF2TYBIELypICCv0ZLFw9PuW2pGWxdAqblxWjDghjh1eNinFhc
AoEzJYVVBQJnUF6esEfRcBHltfZKBzdqd4VqHo3vm9kD6/nnTUol2XCON173XtCm
9UvAU+9GvbuyMz/eZ68JkNLELcA3SP8vZupLR7cApdDmbhrVXT7rv1LenmX7Mhlf
Xc3KeDt7oEAuLVcREEr0RMl5iQmiNqvlGmGq9cLPnda61yQWiKl6NN5p3zdmL9pS
UALSVMLCyyN0d1ba17m86GDx4jpDLi9msNrCqGUrwD7bDV/FCxdnb2z9NeOpjfRw
8wzWPhK/e6/soObP8RzacwPsro/9kx6RRU+u75T+l3La93wonzQm94FHyp0+C+jq
NnGGsWlfJ1Qh7WmVWCCjEp1ynp5Ze+DV3ynO9l9pRWAQhOqwvL/+qZ/yuUuxyOoN
OfUOLdHqYioMVmsadN9xkLUVeWS+W30OlTkAVprq4adyB0ki9QGOGvbEDKqEE319
A7sD8ot4j3/Im8XdsBTyrlljPE0tRzXtiGYyW1RfGqnmVBvbmR1mSAtmgfdCegFg
xehA6m9GQBwS8rgu5rySfJ4Kmef5KNWFn/gkwyH0+2AfAFppQLn03VlFBCmi/7Um
Y62NOIH0G+j8J/4uecxXlOAhsVN4AqG/xqLZDAvunYkb47+DG6HjfAxe+yeXigTj
bNyTJ150eYPVVFqAGt8CAg+QFo30eQdVemwy+WmIjZQC3Rcl9oQhpGKcYfjsda9O
iEav5xv+pECJS5aHB8q99FT+s5yAMqzmcZu8Yt0Nne5L8ZD2zWWokFhQ0YAu+GPS
ndh3rIcJc59EQm1oS+PBVtCXQQuO8Mkn7EbYevAqjNzz03qoK7bz8TnZO1UW310O
MtJCYq/IrfOB8sXaZEkJVGtW5Y4aI2tQ7edNt6c3TTLKXzH/NN82E9H2ZIX4R87A
MX/yd1GusFKyywe1F1RVFquEEqx7XaE+co3pK6jLaCmudRpiNmviZLkHDICX/KfX
dwfPCabVlIC6bnO1kM53kRVR6YVcuw7hYGF/EJQHvw/jgw0a+IoefVAAdK/d4W//
GsjTMaajypq9J6Q0pBRYTJNKoni1d9rHtHd21FcVMDbDCna/i+IKnxKANsFcudrb
ovqblDJv214hGss9MbqAFaIDdXxpUABBogZhdKVjd272DUhAAJhluwwCVeXsYs3z
BlZq+rEFvsP3a+uRonARFygUCgyR7npssdPvNJdozt67gu8pGDktBIAYnJtTaY16
iy3eyAyAUE9duhTqty+wxYVM/pe/2UK96kgBhamUAJxTsLGv+fXfpfQZpiasKea6
V/n1ynKQ5L0jB97afodXmn9QFioKKEo99QgzDV7hHBhCIC3zq1AxMFTcxxMwwqPW
6TGpsxs/g5L7orYij3fRg5OojSju4LDl5Llp6KXusDw=
`pragma protect end_protected
