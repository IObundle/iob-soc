// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N+1NDb1Hg1rWet1QVYMkSymSEZ+qZOvaKXtW3UiA+jF9VSuIBy41hZSoyhg7wvVw
GaPJLz+iqCI72z+IVN48LZlCLwhl0jzJAYASNegqjU9RS259D2K57ayQrafGR5FI
6N/4kwcAZp+bseGNzM6/TTfvhdWG2pVJyXmYOazXHX4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32400)
NNtVL+LjXf+h9IPpIpQHUtu1wyVgLEscwPPrQT65G2sQo90HTVj0VN+6OR/pc56P
gv9p3FTZxUPXG9HCy+W55Zmvy0SC1ms11GsZndwDcwf9jwJwaXibunJ5DIyfA6Yr
3hzHaXyJ9/9zT4YckF/qr6n8GP4JNJwVAtjPwb+y1hyaCIxrv4G5xKJvg7iVm/rV
t7Og0Wi7cbBUF1dVd7RbdSiyypDjyEnGbkn1NsuFuNYQTHZ46QxtaFVepiSwZAjk
cFZm/1N0hKdyULy5l91ummcMvNrKv+kKUOI3p7l7sYPni06qSjQtiYV7Q6QKIOsl
RHcgWbkiCJr8fHkfXsZcTt+SM9VQRy70cwg0N4POG2quXYYMD0r6nHWxProezUw2
ElrF8eUeNPZz5sBLxEyAXaCSd7oYnBkfM95zKdDvoTUHSbTWtPdGuCvA38Mx8bWl
WGsaBXGfGqhMouOUNSTYuDhoooI1+Od5YqABqj30Yvla4lrzSltzivpFiSLCWYIN
Sbpe6DH08djwLC/f+D1B6MYmEY4LSxkPRbvkH7+88SRa2qPnJae/9EZbo9A++gCu
XB1vWbC2LQazt6XLjLJJwpyjAeuWjKqm7DvcmAJj/aKCj0x/VJIVxYVCPDuYetRB
z/Tv0ZZEz2ufc+b1lAA5DAvO4OPLfHlJvjLwRsSGkNReLVtP526X0lpSaK1Eyvg8
AHxXCz5PYB2Q2glkOj+5FnzKL6wvbHu7aTK3MwkgGOEAegu70JLSXJ9cLR0J7H3s
oE5u3t+aSiE9Wwqapuo9qzkc7GySUqb8fPUa6LOnqP3YC3RrwKzSB6a0hn0u1Wzl
4HGI3KPCSlDq+H0AvPujKUMCvGhep6JFFhL9dAKqOOIucg+FzcMRgyTm0OELP7CK
kcHFz2WLNzNFz6a5se8nRxi8obAZQRZNbxFgxcPMBtY0n19i9P5rUqEIzRfDg9m8
pvW6KRbSpWsxqHTQ4QHAstuUkeRtPsffE0claAs7oSVgDVvFT75v9TSRxK/UnLZb
XybWqrMbZqpPSkuiCB9GjDxgaJyKdhnzfBTUbpLyUpPcr0aF6wQyVMlFUSodEcE6
ucGpbqwSqZfHgqAt0JH3GDBFDalZtdx+YgERyXxnK7yXLjZnFPm2N9UII+uUXuXZ
RbuVmDKmf4a3EDBfPo2euBZuRnQus+EBMZOPfAgUf9L6n8jJqYHQA+XCTcGaow7s
wvm2HYCfNd2qgSIxHAkRQt9wFDQCKWTndEe17ytmPU8o9F6qsFfiQoTFyMEcSdFW
D7oxvi62L8wQCKqP0gxy8QOaDHeECenZE1flRxJMz62W7BhKbXtp9HPKyyscRSvc
I5B5AwBxtfuJFrD/n+oCA6Cz0I4fVnIeSN+errHFdtL4Z2CKzKa5G/haTZbDP7FM
8sro1hTBBv9Il75PxPsx6i2hRXs/aQYx1OrKQNQ0nNFP9yXjJfE/hvSly5yoABGX
JEx+7uAoG5wBJSdprC4W5etFx+GfP9geHlyMh5n2NZVsdn0fw8B1JNiu2JA8AkrR
qClkSNkeGJlj4rBvJEgLBvctkzoHmApf6UH1PK/r3uqU+pTssmRm0I37IEnctKFP
SLLw3IiuK/6HrySLhBAkLGItC18MngqMF6bT96VjSvHewZoJ5mEYmflGRO+1+9u3
QIdG2cBUMnkM5tUKdje8ac3RaxcYYLW7hAfg0CatasWlvn29aVUgDfnqBSyH/SNG
/MZLNu9gSvL5zjgoYRRzU2KzswAXkoeYGlPVm9Ajfn4uo4Qmyv9b3ZLcMBQVXPyz
gMj2ipzNUIm5nXW5mINpVmUKGIsYD95C2S3Fx91s8r4eHl5GrcyxKlLPeD91pvrB
gOT+Rj5IjGmUm1KUEtl/N+rdsqciYE2dD1FoslDUc4Q2JZEoasoPLtShjtwtDENr
dJreJ1ICdPmXLEsbkJkhqADavg9lNi6SFxYlcMb9hNstky1BxnPwoib5XiIqrT7n
lZeV2FRlohfZwT7DZ+WlmEfg7GkkjGJfS08iIAKoEltCUqs+hE7WnFqLmBNdFs5s
SqSuF5iVcRZUq68w2d4lmbQFjHwWVI1scMK2sgxcO7+B+KyPW/VzZAr8LJzH0+bT
2WNE1xe5T7ce6dQg5fY29XEnu0qM/XaOTHyRN54ftWTFMbMrYUTz1qZv+q/pA7E4
Jr0DjOTh0aOA7MCIaE4fF/wuHf567zY6UXqtadvLEfHlfvoXf+IShtcwyx8Dm0TZ
9Ez0ag6LO4hn64gDYXc9ze/RoGK+hYLAjGzbFxDxBA3gwZfez1cCqx2vWC38ClK9
VSJCZ8ooC4H/6UbmKXAtoMpMoGs5Veiux4qA9Fy4wIUBpIVeK5Ys3l6G70+MhEwk
gj9a65TvaZpTTXrVJzC6E7mOSpUuz3+CejgIuLEnsHgG+syM3SqdXuQ1e/LsZ7Ow
rqQPkRxFRshs7iACxHurk8P+dvJcs/+GqpKyX4n4HZOmWUOShRcUhbA4IlqoFshX
6UbR6jmfOj5uowxa6b+wrcnYGnCu7j6AbKb2Nv1K+0QzA18O+5onNdB//AcOYoJm
h7luhORnyezxSqt07jX4+/Neve7//5zI0+v8nKv6ourI26Q9dA1WhfwSGH5itaci
TjrtJgPw5qlKQv3VxoP1+lDZHRlb1dRox4sS8IcQaY+x+VSB1ZJEP+4sFwtggSnE
zXK9mMeW+qRab+JV2W7tClVYdbJaaPLizfyebdh5Gi+kdm3QZTQs+8BmP+4HNkLp
k8VLFV0fwHLCGmXpgYxHdPstmZIJkncFOqrnWAr1T4eTMrQA0TXFPSPd7EbRM4cp
K70DI/3D9MreBN3Mrk7UibxUCC5SmWS3xkOWOTy4qZ9a/SW7uW6igKokSxfeHf8U
85O5os3MxE8COD7GRBigH3PVpGmJ7e/MyMiZMfjtBoBLCHpM1ZbZx+38wZNKT2h0
I+ZqB6oKzVss9jdAvknoKe6d/ObH5K3ihuUa6FHnZHM9fvFjR0sXcmkHY0bCOEPv
O8rwX0vpP7XrhXnoFZRg3N1VVwuKEKZ4yz/NLrL3lPTRmxVbLdnfW37f3a2Ek4ug
8NgU6p4S5oA6NY4Edosn1tVOm+zEyFAsBgLrM5IoxITujSV9m3PpA/x3AYNwnY+F
r001g8joGPr8FEUo73g52Y0f18GHvMnliKefcD/ThOjsGNGbqVBImOmHn9c5VlWh
B/eCai9ou+oQbVDPH8UjHsZ0Bt008SLdseXPLRwN5bxKVaS7pcgM3/GYSkrkyY9C
xbaYA/E96bddZ4wqHT3zENhdZ03guS5eLhgf0RdWQxqO5zttSAfwUegrxhbyrGvc
4J6VZZIOKxiSd87f3D85Du5i8T5wqiwAaHuK7RzLW4xCfmkYhx1jJDp4o5yG9ikW
eOVsRe8p773aP4W5NXVLPgk4CMdmPAdFk1PD7be2F4YrPMeqynbpQi7bCurFNvBy
SD+M4mASYtGk4m7wtQUrjVZhVCmqBnzZX87FHqmE9JLAW2rgI6Z6uCRAIiVUL7hG
SCERJ++4qrlNW+CzzelX18AKMEiZF2I+KNL1/NMlYRLXihalKePOvimUX8BFdezS
zYAzd/MavGE6NwfEiyimg4cH0XB4hdRJSFP3SfQvhKTPtMS5Jaz58cUiWGjNR934
L9UTFaUABfHJaWDG9UgljSr8bWklqeMbbdmBGy856KI+9E1FJAA3Sq/GTyLuzGel
o+Eaqf3huAujmVUja8N841AsTi984KowyApTsGjvUeuioaJ/w2yvKxCwd9Uy356e
fU9nqTP7xZOKKf8PgMFXCnBsLUy/6JgcV4PfB2MG8n+iHzWGpLJwPrBFtCR9LdHQ
cqPCkJFJRBWgOruXvhF3zLqSjcHHNVV6tRZC3LHvfME3ql1E+156PeW3K36j9uWM
UKVBiqRcYG9IOgUgza3MJv77rS9kUvUbX07yHsfkRtV8Erxd8yNtKn7hZCBPRmWE
153H+2d8hVoGpHTWkUv8RebbdzmbeW957z78v5prVgbqzSiyC7Im3sTnwNJ+u6V/
lGbgF2Hz7WFNQ4SI3Jogwxfo8/K/ZpmvZJWAFS2/j9NMAIdKlIdpqzAplSBj2bAW
xocQ3A8Dda0QHQ9+AcyKKnfaLYeUL0f+POKOHByDui1mcoF/1FyICbSQVyc5DGtu
uY3M/7ilfFXORIHOad1b8FVJL6eT2xqz2iS4YZIb3vTmf54tlnnZvkb7oPeP2ox9
rh9FgHqMuTkDv3OnWt4oB96v8jCXO0xuyLZBtta0wNn1N+KrbdchU1izb9INA8hg
WerhotkRAscWww9Ej2GAwv3RLumDG1AOdfQFdkTwj8Ib12lMOnUe3Z5JJnWMkJli
SAntxsbhigPMXbxWI4yCFZgkngNcwrfKwdQJXRA+kmasmnDN8f24xc9NAiuj6ErA
torhbzn9mtcU8f8degIGaoXvgGpw9q1oNKsYeRYI8z6lGyPnLTve9LWCd1XhvhUR
yywgM8O5ZHs/9eVhIiJBjNDhQupYRZE3G6mcgIXx+LwwCsjTTIICn+H9Mh1RGBNE
HtLykF5oNsmMpdzV1+GvsYdqNuzSDx8ELE/SgUAs3gvwdf7uwknu3/nvxgywuxD5
T1bn2YZe9eSh9xkhnpP48rJGad3V4GMIoG0q3CGGUPHVgQsp5Ke957n8QcYDp8K0
sCKWVY0PZeorsg1A1ycidRfzOuL0NBy1vuuf/FDPi1dRLnG63IrIbu51tgaOMaVi
cErGF75XuAVR7m4Ca53UhNDZODF3JNkx6VxHYELxBLyLSwlHNhJL7HlpGIOiUUnZ
JEcT6SZiTxO8jM7AyBaHHZ2cr6muXrz0ur84NL0psGApO/JUxu+koz7JkYFQkj9f
QBpHVsMAv+SUUwvV+C3hJ1ZdZMaK2XNR5ExevOdb9N9fuZQwhLQbrYJa3hXe+dDP
lH3oIJ1r0Dpbn5SOePceG2DGI6XOJeF0zZDngg0YpfnWu/GN7pWlywi2J7exWxKy
fun7POVwG8GJg3qIojHkf1A5EP0j7YUSdPliNwRRah4uYJywzsmnpY84bkii3pT5
H/gGaIFrRvq2x+lJ7sQ2fNldCCLbk9ypdapKak+3lNeUmFnpfz2hFrQ+5ACkJmQL
BZJ4Bn1t8SPz5Qix7RMmROC+BSTjKVkn2KJfFH6j1RYzMAAYoUoJqULZuJ47T1QH
32LjCtJcehLg9u6TFVlqktxg57nS40yvb/IiEDrMDKI9ejaVHXOMWh1dg73RA7G7
kyvQRmHIN7CkflmQJO2DSS/hV6kEW6vmVCMCRrKKFkSsU7odBB4QBBzAYdGZTtdF
+qnn9Gl0FO5itUXv+gef3sbDvV0zEi7QlYJGVeyLLaC7Grcp2FZh5bco0RvsbReO
SVBLEJZ9MRAGrHQOHvZJz6oZu8oV91prxry8U7VK/Gs29IOTFrc4G6mgVs8939Ag
tlPNnT/J4oXjy9QJuEmLspA7mcIj1VAKkEONd7xzmQOR24ps57awl4UaTHFQCw/9
iEa5UPWeHZDubSl6io9Ty+9vPo9jJeoPizAChhgLaG2snByKu0kMFcPLZJFnOlWP
Y+lSVWYtozp75/XJVOXvRbN3RB5zC3bhFPWYUvxBlSefx/NzxlfWMvDPvqcpGcmL
+Sj0rQxbPh984oMxa3TbIG3dv3c+o1wkKna4vYD5hH3+So/UMvHCO1dpArVEtO3z
Gad4XHWWJrq98QMwFbxdno3PyR+SULV5d9Blv6HCaj9y5KjtIuCRMxfs8GvYG6l8
KpwFSjlQweUxCuoaINQgcPKDBWpWoO3wVryKgBehIzBEk04hPIPUrTWX/Qgv/Szo
XaZpLjHhKZst44aMYmr9UrDo4IILxTT9XwkYnqrQ91hx/U0eFOBW8vveObLTKauG
7R+bJ6fEEfNBJQmV+a80gkVfiLErMgqzCaT+TtUQeb59lJW8MV7Mbxp4UsBKGr0U
eZrxudphQY7FxqCsNzZNFewbowLyGHQYzvAflVsn5aatqSjcxKUm7Ed340eo/kRj
L9bCoFUwqV0kGLkFf0JALhvw60Oswy9LFSSUBXtL8vOiuedxZ+RglGvd2KAojl14
EMGPJIQbPHzuRjSdP8Rx+SLTt3QbVxv5GmwxQIFQrbQSdPTFscAs5K6MmkFw88tB
aPCjaxecExIgrI7pK6QIlvFz7vDpr+sfUBIoPF17wgPNJThj8fMBPxFxH3ctmoqT
GdrBvWqRwD9XbQ1ouqhZXMAWfCc8Q1y7unTs+aglX54KhfWuBPLkVEEbTslywqhG
Q1/ussvU3bIDcpxT8pGc4+tLMMzQnBxrFHgQRb9S/xJlmpYgN++dOGZswEae6yqL
TzBLuozjN7bQzwB7ikhV6PsP5rXRnxvSRer0YpfdHefm+4tqKuGi4X9nirKKbzgA
1tR47SltcK4Dnp9kmJXL137g00hppzeAtrSSZb73PSrX/rupuD5UlBnxiKF2phd0
OKgaEwUbynJD80cSqHXSfQjBgp0HkLBtg1RloqmoENpzCHeRp158q7qooia5ciTm
a93Z4NvBrN5IuaPHH75JbENoc0Z1+8LNgEIGuPs3wO4AtW1Vr4sfRiWUPb5yXcHX
GRW5Npr1Am5uGsvCDGvL2wTlesiCzyUC8a7Gort5j7VxWuDR8+Oxt2nZU5KUEax6
GG+CCYbBDZvjmgeBiAKspGzFq6G04pNMLgjtxVyvyGtaJvcT07kCPdJcsZPzvzyl
cntaDcLEhgZMwsUn0T/yISzZFJagaN6RO67LCyjUq7MmXTSneSZavlq3MYpUJ8LS
C60jeuoKPhMYhD0AbfXQJ5uB8qGjqiW7bj686RBIy9Sbxl7wJDwnf4Xs5dzKJX4Q
jnEpiYHOAdgDnZEr6xG5PuTv0gZ/n1VrR8ADnx+hy56YBwnivqN+qb/cwBBXqEEo
JQ7jN21iM95gqYcvxdiuGYxmcR/+TgrCYTQHxkWwKXWPOjTdp3AF1Ux+VipOtFos
OFTYqqT7ST8AZCnpc5e/n32L63n5laxBzwMro7EChnqjoM/Tk738WkS0dfrWDwtr
2kTYWhlMXc6qs8mR7feVs8rCyhEYHrEfgznhbxDybphDkmoRGpskn7Z/XHiSJmx8
U3wxEDXyIy7/g+0TClSvxGzsX3M0Fl8tbRD7eV8bMLysIxccAYMnU/pLrIABC537
853/rpuZZKW3WlA+jq+iCEUWo1iAtDbPzbli5TY/foCGCkuS0MecMMQW7I4bDNYU
Koo79vUW7Ibga+66UY4/qjxhdO4Yah7BNpdMMlU3vc+xFH7nkFcEy0v8aik4uh6k
2mgkmaRqyewGfQgbmL6799Dzq6ZHfL5gLRULZnavi51zUXAzmbLr/NDZuzmbFSzn
sN5Q9vIt/Rv4Umi8ppgcqSDpoGQx0AEf4psmWi7VCLmHLStMvw8nWOt5drjJQJ4f
ePBsOcxeHvnonMNfc822lmDxTgTX42uagbKlCM137TMCjGaRVeadYB22rvP3PfGk
uZQlInD7uGYGuqetbXnGg1WlnwSjKRmCT7L/sFlZY0vKKULfT8HJTiIGt0rhtcmw
reMkhsYJXhsF0NkGsgg8F/rAqoqaFlcu58JvFpclfj1T9TjyEIQDpR2O58ZUzYcy
lJ6akR7kuf7yJF4+01KEl1NOKyHBFRwZZoRq1OrwqKKznsRUky2dzTRHbyqhijBl
Md8KnNm3c39j+OVvy8N/tXH+LWc7KjUzXTrUdta8U1dITc6/A6tZovdykJ7SjvA/
xBi+9nO1P0bRLqYCciOh2evwWiVS2vgeKAQB32LrgeWejcJ9FlsZbpPQshCGzod7
gmR+l8gtK1FavRsiW4JEgeDvg82nvSPZLmFxCEBd0shzWZy9IclbLZgzD1NQdK1A
FibSifsvdXYylQO5Mbql4kX/fAGfjpF4Tyt+D6PsB+lspDqOV+/3CqXM99TCIw7E
VMrrrU0Xhli0+yevLCFJnl/v7QJofGTjCUDjdoJ+T5TQzFXO8GTwFhotUjAhizK1
y9qaTeQ9Qud3DrFgHo+cCef57o+T2dI5gNllzjvECV3HiJgbY7OpYZ2xPVROorXY
qSL1zoVI6CcDy+kDsUAz3HLDpMAEpo4G/f2Maqq8+X7FQg18DvbeJZedBcY1Rdh/
giyP6ms3fR811m1aXh1S328r5hJFjrStRofHpfSO2Wf9HvzjTjJDhTH+tU75fNKf
iriBByG1e6IG/nZx9A09BHFwXkAuJMi/Ge4eSCaA3zBfiF4v4o8G5NPNrlnsr3dW
3rIUYJsplxehlCcPPqeWIu+Qcx00XDhqHw9PBkVddZfwGH/giuRSOn9Cf0o9pyCT
tRmiJeuZFt+oza3gwy9LkhwrIjzahzo0YkeEeR/2GAtjcF9JD9TBTY+ptJ5OKlsT
rS+hHpTVJgyjMqgxWY9Bgyvjx3aF6wi9xqSb+fQuNOSpW3tItd6bU6OA70SPjaZ5
ZGvvnIUUvSaNbcu4bk1uib6IXkwLmnz5BS+V7APZkdM19BqY358KaD9DMnoyWqMJ
WhDS2/S7tvMXiPbgFICcecORrpB2YLwM1bYO2/sO+jrITimNt7s/KEIwOzANFbpH
hg195aRGW9+M+r2yf9TvW/FsM2OUARabj8URsLgQ0oAcoD3bZsIABTm7Y3FUQpeI
OX2lTX9bwSlXLAxyBkGGgTAZzSFCEnl8AubCVIBHYxKgJ+oUJ3adqs0fB5SO3jsh
QkPj9rYhyCL7qtvvd8KKVoc9syg8W0KcVBj8NNvbekswG0ahI1oX05IAZ4TjEtWp
ft56i9UR0qlCAm7j4ZYDyIVHMr2qpd+IvJBnDnNmakID50Cw2w17SnG8vvTmGqCG
bt2ODk5XjZDjZGfM+7SWizj6vgywgrg3zXFYYbC143+vtUmZDjlpXnMFnbYVBUSi
fyaPATLfczyqt4wTKlMWIqtf4y+IHm9J42+19akNG0BC9O968UqNQzFmOR0umCpg
JjLwTEDbrZ7azob5+zm9r8r1xxIpST7n4rmtfVL4iFjP306Z9Op90f8HC+oj/5Vw
DejWGWEA2fMDs3pvdKB3PiSfqgxtAZs5Ddx/sYCzlLqEpnstpJcb0E8TBh/9ygxT
r5thggD+wYWrUAyQl+fHl70iIOQJz9djw9W4sNiMcWpzzI6Qel+3AipiU/GGa5uy
T1WXqNs/MJHTS8HOM9xkvkmifO93i3qXs77wc1aPIOS7quk7V9Vp+RzrF1pHUpPr
R6Q6pmI/chm4M7gW8xgaVEuqUtyANS06ZZflYuocruY5dxVl+m44MOqkP3zHGYNe
8bbXrw/+5cZGP/YHlkx0BzfPRMOXtYiG867jwTMM8VX0qopVOa5p2Cu9tr/vGAf8
MRFxyNPtnBKLGlBxpm0aZMVhMU3YvuQ4Em/xS+pepeyEoVuLv/yLRdoCDZBe5DD7
7+uGSAnKtq+DjpRVmJDqunCu96PJnn1oCxM6FFBk/jfYcUhd5H8x8Po3rQHTqAOn
GaTCS9/gkZdoUxzABgXme2NwAXbsnoZUWHIgclR2k/4rYX/NlEj9U1ItqzylALwr
4+wxK+UIXOCLkyOQYixBE9IwTO7PkiMauUD3ycIOYQEmBvYPMXD6ahibz4p9FKPd
Ipd/4RJ42TBQqJyelZk6m+KC4Ao+0hD++wkmc+jQ88mQmGPnM/TptNsn+0Sx78Y+
87p9pvSTvNvwNRQxO8iT1Apa/cusvTJz7qZ/kZNKE7nkKFUNzg84O+D2OU2r6jGA
Vt76D4Zcb0HoYlZM1CiHG4NMiL1PODv4FvZHlXP+w1KVg9D90ciPSG0TWaTgiVAp
igE1o5GZ3uhLLB1iwaWA5tWjQW5APl1O6AOOqxOCfjiOURDeKmVJatd+EBERyVgq
mQEhzCO3a1Ei6qmZmi5+2Ql3gfgOjlIvtQb/ViPGqEkTQUetNRBU5bbsX4/zsfrv
wLB1C9rksToAGkvUB8AN7YGF3YvjnhzNg/8fzqENBFNq5WGajyyzdMhp9fDoRlRz
BzGHrkMwD0WEIlOr4u6pL585aaUiDK2PVVu372oNpmxhX/Z16t/Or6IwxS8tj2Ud
7zwRFnEeSeibfVnSuiVv/qB+ctpzkyXTZRBtRCcMHxvXFz86C3+3nMtdxIefTXtS
3dL6AEFzT5izJCfpgHuWYxgSMDWvKHlrqo3ajPOLtgRD3uCEuw6Ife7mYW5NZ2s0
g+0DCeci0Pk/TlOT2YS2KMT89VVaF/ur/DCCU7hKd1qnBu51wJr6u0s3ZsDnXO1H
TwlqlKR1q0AxUBzgOYA4nWlY94HyZW9PSymGtyeEJrV3KD5541XGI8n3YNAe5Kg9
NgEDdEPri2ohdQsYicP/v4No55FT6uBiLOJfXQhurcSOxugt2XGTsZluoLUz8jyC
QIDNJoEUU+Cn7ZGXBQgeTgxcGQxoDfvQKtDZK02FeLuvpuMOeUsUzNs75diFyv9e
7ExI+vaxvht50G84oP6mRNmL8Fd7ZPml+MqGmxmxYJTojxt3r5mAGZomdhK2LgtT
93zHx8T6d9C08kjw9oIPUla/y7pCKdZw7uEbQQZPT0wWE42inweUqGvOB3O6evxI
8/0aKLFmWfkK04+V1wRf8rdguGr66vABxAp7ViP7DJlXV0mY0nr7ASEXG3Cvj/gI
YzzSARf2KdyUf5gZOsmlrx0+lMv9i3QPG6IcSIMgmm6FkXmVVRQoqpt/T1t3PBpu
WY5I834YV5QKlpjVJh2n/Set9SqEiZcXdZ6yZcLgUtHTotvRwbLqEI9rbtrGNUET
jWH4kC0Wdljc6XT63csUd9DlbPzWzyR2NVaZspAMrXLwHBo5teBSZpUEPc+ntIHv
dDkVI0f3OEy1RuZNWl63RWbv19ThkrNDyFjBB9GfdibqhnArLMr/uTfA+qW9GmNS
S12SBG44BfsRu0Urs5Aeyd/MwpWNjUn5TfyRSgIow8o/Z+LH7Lf14R68bAHjJDi1
ZImGyUTXPYV1vjhSKyrU3tnqQL0WUrJYgeaxg1J4RAw22YU+ENyrSIuJTCdAOnwj
rlmyDZOwAym3m+hBuji9d9J64y0bzs5DZloj7ppmVz191RfMuawVqrzzKOcq0mpY
1eP91Uxt2hKDW4jt9iatLNnWaBpeb/5GUzeKJQhlaijOG3UAplyeTJ0e8ljVZANh
wVVfFi93TFigAGoiuVknphP99PT48AWnJ44aCGdJ1ZFwxFii7ZSM95JVV+mEtMig
ZZ9ulPWkvR3MTjnbcoHU+oFOPH7XL9wB/ppQkuTfn32SQ0UqGCsqk3E+4T++ZVSb
1oDd9EUZte5mKJ9QZOrvZGw2rre5onhLNHMoJUWLkobyEXI2w/OO2HHi6BTOQDxv
S1hf1A+StoqwxDFnUYVl1031116zSadJ+1os1vS4sppqjSNB+eqyjSBigLqbUVzw
RLH2FTMv6hdYxWLNf+zdJK7YM+QTVUhUy0Mzgvw79H1pRvkqk3EkEHmSDi1hSlg+
cc2gUOSGiNWbTdEQqRYRWeiAtNQiXCD1nP1yBXJSmyreBmGnO5nT+qLiRCaKut6K
bsShZbpJlwrstjXy9qMCn65E9aO45ckwNSBheyYmovHkqSPcs8dE4V54USIycoqr
TeC9M/laZmjGifPWRGhBrqpTueW+AS8a5Qry1OwzDojrvfYqno1BrZ4Gr0KU5/Yb
i8SGmCVheIndYRb6ebZUbuGYD+D15pmRLh+FYRYghAeXewJc6mvKFcfKjoII18Px
zJXfhIhcZRBb2jKQKORL/Ex1eHzWSmnFaERqzNV0Wmm21fmS0p2lnYxtP4zcjHtK
v5MPUrd5kKjILFVIwOU5pSvQ4y/ArhkXxYMXpcsMC7MTDNJyldX7CFWdWf4aR1M8
LbR8u+xuR1tRCT8QVtt4Xzif9tXsutVjcpMyWMVQVGnwn3i7m0mgB6ht/nDanBc9
Ja6Q0SXUxRWJW+9kjvWF87kzVL+MYupuJnRxk6zImykqihxrcvXP/3/g8gd65e0+
qnsmnHBAb2KGci6nJ9QXSvGBFlKFkBCT+nXCIuwYKPlFLHluLSQbX9FhkbtWyKzv
CwXCyxEduZRaNaixsXKEKN28aHvuAEo5QIRKmu9TLYjcoKWAtofAQA9Uks6j6XJs
Yy62e9G2VFw+mmu16k1ZsyMI23vdXMlFwUsnd1oCHh3ejKYZpemdDdWdTv6d1pQ/
2hW+htSCDo7XwBaQ1rVizGigHFL5xXQ1BBG3vyWqN/Kmk6NvwrhlNhkIySB+/F3N
KiMLTFm/ykGbFqWLQww2/GOQ7Jdx7kQJiAXB7FTM9XI00tyI17CuESNsKnIPfoAs
YEDID2xhbMWpg6xIKoueRVVnUxZ1ekvVj0CDqL5Zqpax0owJrhmtYqWjWlu9EyYc
iVRHXq7pQZ8bCM+oOUO6VknGnmFG1ljS1rfk6htfWqHOKO3qYAO2dgs8HjLnQ+w3
xSSccrcflAbuJizFXzdIg+uitNOVdQVhLoEsZNshtu3fKvu/EgK1WJKnIBBTkco3
LrghUe7L0OiKi/90Q+XZPTiRoSs1reuqmCDSvb7wp+FAxl/gp7+oAziEkuMg9Hf2
c6ZzG9K96GVZe8vSYL8vGVg2t2nXEsrcwcK4UxLfkn6yWzttXn+GGvbDCOxY5tzM
Os1za06HlwjMBctR3lBEcwDn2M9NR9rFJyHONmD4Eqs9Si3wn+EZXQzpyoHr3mRi
OKW5UXXEpE/OtZlq6B2n+Is/73fiII/ttJMCWBvp68EiAQOsx3vQSF+0ZkSgURTj
f/kMPMwO8Wc/sSBikaVNB/NryoSPrjwR7O7iEqUMwxkVYAgt3XP47aTUw+kWwola
0bT6nZUo9kR/ratO/dhvpUUl8jcEOSFALdJNO1v0uoaqQR/eNd85tVTNiYR9hnn0
92HZ1TFQrHZb5hr9tO2pxN1vdUhvH3TUZ/rL+ccCNXtAkaoTxyA+cV99ULmQDnQW
6/y7xwtOrsnIXS02lPqCqrPXBIBMjiKdk8nb7ezWm3ktqjYBV8xbPfDoi3Rcw1Mm
Nilodg2LkHOijuPuURo9KrPsGHUTAODVEfqZqyv30x48a31jG3gQzQgjowPVwNe6
GX0z+Rkz3UWkKpaWcjkBIk1gaTNuOVgyrXAjms+JRw6Ox/P2+hm+xRdJbjHfEYVG
6/mrl+HNj4qIecP8dE+JwjCakQce4cFxzp9iWXOG560KPSIRaHqW6Uq26o5JkcEp
TRViX4Daz2++Oh+gG/uNV9icsuvO/gG5FsDAOnNciMe5MNe5uaxR7jfxiZpfgw0r
UKaCnBrCQISQ9dNZKCnv1yX18Oz5lrwIYascjXj1fZBa3dNa9FM0QW7Ddh6iveu2
XnrbpBZu6MPCRVOrO5VeI5e90I3q2eEfj2t8m5BH9K4u3xF7YYISQhNCf0ugiRsS
cknzNWpXzwHKpeMpkLG0tUi5rjUGt5TUas9CF+kyfrMr4+4LjW9QBl/LKul3Eo50
BBQx4GdQ4dpCmabhvEos5PpFXNFsZEuX4+lwNaaPldn0bDvPeA+156ILPbzLBer0
ICa+uX5FMfk9eUsWKpC9J6eDrKhCfZT/hoSWfxB4dbVwi9G+a7PRzF8b8+V+0Ji2
AKB7SSx1xobmJXWIFSvHcyzMW7VkQv4Wmx+YWoM6lzY7d379CItBXkycMcTTcrm8
gQDggeSn5TdjsRVGT830NTMSeDEm1qlq5LnHZQUVNTn50m/tUMXOsnEv8rD32+Mt
UL+qh0s0svxsOwa8wwpfNoovHBEdeILSzO4Bo0YMmcNfAhh1tRJO0PPoOkUdr2f5
8ZFRuA8jfwXxVsWcpq+t2ZIOMwtQZmBKR9nuLtgSh8s65huYmpQhm3rgDtp9tqjO
7gVDZ2Bo6mcl5+XIla00n/bObLme3Z3FkufqwcZTauvhvIx5Z4rspQ/RldQOXhz1
yKxopfQq9622plkEtz9+8sob4uHQnfQw7DxeWkMh+uxpObU7M3E5M4h0GJ7oHt1/
uBdzehjtJ22CqvpnXfQdGTAu7LLRZGz1xa+LqaHEYgA0rKqXe9LRZxXNpyBlPMLs
kN6cikMMjIx//sjAVKf80yrgR/2heZHIBqzl8GLbyt/zzwuSADU/WT/Nf7Odc8If
UDAbXfrrnoluxGWSppZkI1aV0BvmIAWC1puf0oZcnnOJMTQswQRBCsi3AUF+ZxFR
lMvNUYlfQ6wJsG+eXYcwy22WG50jHxP5igRl39uVaPZVWDyaLkdiIDKqAiFcjV84
2GRS3TaudksNrKEg8f+1+EgbIkdvwQORJ30HL4ub7Ak4GS/lCzKRC982VR/xWaW3
57lCui4gAdtQJtWOZtL3bJQoP+4ohLezSFup7KiQJ7e0HWjZAcexDgajD5zg88I5
6LAnGb/NhAo3wDg8h98q/ygyylNuj417mNhanjC8bYiyItMGkoEsb8KHi0id0Zt+
hqqm5T+ped8Vlv+KRSG5lRMVQMjjBIBR5tMCvXXL57yAkEVUEpE/v/OvKcC/QsYB
Kr5uS2FddznWq7W9qPQUxquS1jzwR2wCCB6w4QTj+5pA0BumgyhlHMoG8cnD15px
hOvrUDyP0odu5mXlCfxxUJKPhIajA73CSrEm7MMmRJeSKLmT5HC//S1t3g3UxWzB
Dw5DoAkP5256zPKdEHxzp5lc0kdrKUblZUqozn0028+5oH93EOj+mtts6tRxLsME
FNFcspNnZ5wf4NkBjytrSQWkfzGV22hbOx2eTKBAb+V90ez41/UigppX61Dn+ylV
xvrE+TosK+CHKVgdRpt7o0kAV/G9yR6BU7ztEu3hye7u5YPlRyZELZtt5SBfj5ny
6UMHs+U1bsiOz1UmCS+F6dgZpJGia8CVBBeOdkNciH1dJMcorXD/CMCVvdoK2bLi
KMsQg7bVTTxWsw5gccleyx3FDXQy3Ik0epDzPwOAzUWD24eKHcT0IGw71x2x7YoQ
vS0C1mM4xHColomQYdOyEdrtKh7NdWDdyow+JPssyTqPTn+40fSqshXJunW4VxQT
hrfp3Hc8sESBNSA+YS5BzxjQVd9hIFB3CL/C0+wETCbThq595KOj2PWtHUAfd7vJ
m9RvZ4VXws0cROERyYdXHoXD0e2ATSjWLs7ab8MXoGW6Ah6OdIv99GjCihXbzbxN
ahE0Lf18IBjz15rENe14OPJdKwyql0UA3ptOwGGmces+RYUi7/PV/YlkgGih16C2
2JWtXbn/TKNRg+t6UymByGj47P6f76N7uRy/d6TObC++6CjH7UXYJmw89o/XutJK
yOi6nxRd1HrQf8mcrAd5W/0sEe6JoE8hpZ3TnPCtxq+i0Hc1OMUBQX3hZlEtmVqE
kZdPUFTe3bz0s9lvE2uifqxC/wrnIxKHWw56yoboSypuSn6hcE+vcwNsh9wxL92n
UjZYf+R896dgK/rgNtSX+Wi1UGdLZ8f9Mdp6uAkMFwsrHROuWnK95CNbVkA2+vDn
Kocgb0VqUhTEpst6uiJNVBQkxHKyddhUz0TPSCGhXW2KFmU5rULDouRQxhdM7jJX
Ym1yg2KZRUxQfSMh9353hRtF5MCfascc0k1/8MNUKvKzay/x2B3peKrHzcCa+s76
S9WZMwFqyiHVwGqijxIw2+WZdraThzuvP7cRABmj9g75isV5i5Yl26ITI/kG7rVE
+NsOoc33g4qKMSUsVb0Nc4Ub/40lqCkrdLMxSZcomFcvAE3LTh1ZANB5nmBhWFkD
RQiq4k/LHfgavyhgWZ0JUZlvB/lLrEOYFuHcLBGDxrFsWbdd8B6unvxWpLVCOuao
kn4t8eiSb6m6nTgjhS/QYCUXo8X/9J1GUvXjksbsCVEYmfuLmBxFn7WZIb20k3q2
fIjj9qvr5zInNm764f3UYZlp7LEtXbDOlNyV+F1qRfsuT9iG7Yv+zhdHEIoCzc6e
RlPJ0/KyP1ggAfEnaIHcgUt3K13wr1k/G901G6VNJfC6D6mXH/iTrtyTTtLqKQmQ
kkqdxcj9Yk0DudvIHCN7tCqGzaJ/A/Ta3DjnzGi9QOkVTodPXlXUxuPHbiPwitD5
1Ju6bb/uQQTMXbJCMXwJJiQq5HeQYmMcuT6KCDmv/7ROEisxjq50Kz5CZSyP3Bxf
sa89FqYYOkzGGinMHIqudaKVrm5i94B+1DNt8JX9feJouAGf9gbxH22cZnDfj2ou
oOeSfL5pYdpaSDT+UUuu9wySKQKf+5R+/NXCU7QMheRY/gLbmJNn/ws3CPbLmaKI
lY5v15BgAeYimAhKk7SvCLsU1IXX8Gf65z/sc3EbM+ts8G62udAfREn6Z+LZeFSu
qMOHGsmHlwtgV4IkbioXkBOUFMi6djKQzpTk6d0mhZlZWzdnH6NvzrdaiK3ctqif
OnwGUxG5GcmAbLPSKWjJxlIqTLczVRl1CKZH2ApgoWjbDWapox2PAi+8/953q/Wi
b7LqLs20H+/v+fGK8wPEPCj2MTUY8Z6kOReMg+xQpx3oUbKg1EOqTRfmNwV69nZh
iV2EE7Y+H8AxLsK1PnEhJ4BkT55MqfPoqOT53Qkmb8TVe2Xg7wI5sXlfhnJCj8zp
MQ7X8v92SnLtTffW/1X+kLLCav6dB5WF2NZgPtc9Spt6dl4OPdlfB5LQOxfyYwj+
VsieQIENPU1x5a4ly6zLH627oMNGv5riWxzu1j53SAt/Ugtoo4vesMWzEFcSMNm5
ObqbV8l+ZzHOkBaUWXNbaT6l9rqmOjelNmKrzpHax47zjauKkeUSCNjlflgLwPx2
VYtEw50nsYYrkrM9YfuVxHpSOwNJW5EcOao9hpecfGWkfigI0so7zDCigHOAqxsv
81c3ydC5E2mnazqxMYL2PsK18ZL9bboj/3C+ofCeDJPqOPlsuZAv4InbfMAUp4Hc
BrqrtyvByEnq0NvQOUmtWBzvq1XqLaH4wXpoHNcH7HOORGWE80xvoSQhNzs1Mqra
J7VTe77zw8KKBH0E326UiPtV4ro/lz6sqVNpLTeFKBCaE/onVNh9hF9cquiWkXmg
c9poXo7YQJIQHh+8LDFYdrS6ZXXoLgeDiEDb3zKGQ3+26OmaDH+Ftxf9bEJAA6/P
5+hsgAEEMlEZZChLmO6IBHoOlqgfYcn0mh/i5IzCIZrGSPeLMsMk6OIEclMifdvQ
BH6ADumGOMl8Cs1QL4gRoyNN0uxCz835rXxrBolu9jm+Bmz7SS8rY3CFSnMxKyPg
+JCuXrxkb+Hoc7T11cOgHH0HMNdivgq7TM/jV03UWAUUyMOEZnVB5vmXtw7QueSu
b+ogZ1XvDaSzJr8Yg7NjS9iHnRvwmOu6WC2qffke5KJz8SLvI4TBkX7PAlD3WSjL
OjdB8rUgU0f+IHB0lj5AcliGdVG/6Kwkbz4QD8Vh488isfDhs8fcu36pi3udZUBS
ZemGnvkkw5eMkvku8XPYTmmuaYxSl5Dl2O9Q2YQYEdjuQ04SIugmDbpOt/kaJoEt
8xZ6pWSV2QZ+NMovxDCLMSRpUmn/gZN+irCXo7y7xfmP07hzwqagN89PwoWV3yhm
QalFqs/9rFz+yB16jMYUJbOMlKnfvD01AnK9mQ+B4iC8x8U0UNv9RJwDJWCeRZcY
XBukInc4Rn50MU5adfFTZ+w57bbdXblPFCK4ROxcDSaYEh3uYJssqhE9/ImVwIqY
u9FkpTacIA3N05ITaaHxQy/Jnf8NyumnGXtM1qpGcAt8miii/bfhdcfH2j+1E+77
luvZW95eewBKBzwIJkmGLDl7uShn1DRB7D3vZonCMIjZuNhgNY0Y1MMMTgi9Wwcf
lHoGv7k2hvt+nPimO1UL2HzmH+4N5RTPr1CDkQ3qQ6OhpmYyWT/2bFm2VjLBEsQN
mE14PEE0fRenLHBe5l/OMFcpZPan4zSIaqs/JAf9TXweE4NvG+v8Ij+9VM4b3Ffa
qw9z/kDLIkgRaJfYXfo7CeRLEWvVsPQTOhoVqcvOT9b5yiVw5UuTUzqJ7/fqaEZS
E9CfVXn/pMXVVSS1ha2z7Av+o836t7k0G9XDh60Y/c+1hoS6Df7npPHdbRbPmeYY
L0/pavTOmQULa3RUc8OgzOChtOAFr4kzzK55baG4rBUcWNbUAleEZGp5up9tMqUc
cv2fLR0msPrsJ4JqW0WoaibbbsyW4zHhU7lltZfIRKPFVvFMdJ3D8folPumMnVC5
nTqHhhHHYzGGUpv0Yb+nqOdRZoFUPnJUj+pM0LJ21AJgM0tMlpHHkZEwx3BJk0WM
bqE6WBvMv7/gcmQcRavNRyJLKJENA6JN9ZVVxJ3Te1I+CZqVSga2GuHDUrai8Z8K
624HRq+LE6Mo2qubmuLQQQoWytstwzAU40UuuwwMl5G2X9VtK8Vac3zBPWDuVxSK
cOe5B26pSguzKbxdwNrXUfNtt+yOgZxAm1mMiIqAHVqCDCIHQZG86Ujt2Ufz1gjz
0O4NfupUi3yfq14LyUVZdYjzBGf849DoVCFFHnjpwcP06AQl3D1j9sHUNEeWCLrM
tT3Red9PEQSjIYZnfH2RZ3+MvVDqQ2KnTxpI/2crxetMc2F72KdebfolquM5XA+u
X6BLruPjsHC9q7xDo2kBiRv/WDV4idcLXHAYlpLPV7n5zJuXLPgcjMiRVMmv1rsr
C1dDFWKMEcE3QvOzD/lENXA0/3aNQIbpnRLncGH0k3bZaxZnkLaiSVROpMdJErsG
WwKylkH26Fg1vyqhHyCj56rYIgW4okNqQ5xo7c+mPBHewH8CsePlXEQMW0Nx8ojh
WAmHA4j16nrvPUu4unzgLmrVgHRWtQGfG/TUMoKdUPcZk0W448XNqrMPkP16EVxP
yIz/7OfpgThe8oUZqDdON3wzJ+siGGFO8zjg3Nwd8e7NVA4XD036WjZ+7zPl3kCp
oT6m6lwt/lznlaE9n/FJuHLT5sQPmRSJfJd+HZBVHs9eViZwxpKXYI+r+szCzvmr
BkHzbmkkbl+kMdT7WIjMUpU4u21PGkmMYFvgfsmeRRfgZLPvg07DMBFSlwVbULzr
TtPJc1w62pKeWhyBKqoKCb6m+hnw+3Vv/iLI8by/wuYODrTds8JvwY5AWtarFRAE
AAfmKhGIxPaFRQIwzrIccihxuW/NyzM7/9UygkK8nJUaxVENRKGmwtbAYbzg/dSY
QFB3pAdRv9i7uitYcD+KMzG1ajt1G8VjWTvHCoN8sBwJE8ACG1eULLKEIywiwLLN
1WXiRIvSbpBus6uZlJCQcHIxTs7EnTUlyujJ7UvvKQ/JF41tu6mdZwpBNemjkZq/
mYA0H5EBTqGxNzABTG8oCZjpHHYChhvIbpfuuXVS/KIqdDnR1uLfL2pz364/7kXN
ACg1s87QY+I+0vrWaOfoXuxzhf3zCaw6lgqYSLQpOENvgNOfQdQ1kj6b0RFBHsCL
qHYt3TGgj9kI2ao8rbDE7DJFO/Ep7i1Tw40FOlWY5unjns406XPCT38rbO2odSU7
rpEKp23V0y6EGETpoBUfeDt/xnYIo4IHRAmz4j5SiDnO+YdSjSJqamwbBJn/cG83
BqGXRlt4ySfF/mkUzUNGouAQPFx6FPrXlu/mWBjx7+u8s24aLd8eBkpQo66KXxVa
nw859pDsAEtKr1wjkpU4Stg2XA6oMixnakuD/69NS2vcGlI+UkOuhmVaN2NA/A22
CplE+mSwfPQgNfJaq4k9BUYxa32GG+pEk85kcv3/4gPN7ALuUFVO9o0itJ72FCWN
nBtZ1hwd/QRMY7T5jpgthfXSlnir4I8yRmXSq88zfmwi6zeU+BXRf0jSMgDW4Be6
0JIbeJR/LgV7IIgWlT0LPXlMDc50PVENHpYuRQIvCLuzhv/RY+JH8o1k8DMaXjuG
uq6y+/D72znziMxp/TyifR5t9xBnPLJxJwwx+9QQUtYX+6AlQglZXVEkBa3313qC
FUv+xLEjVWLmwUCSYW7QwF71D84HM8kjPa1wOcGRtQM2ji8DjJjtWbJNM0rPyhMv
J1NkYcBwx5w+zVE+ng3x2DVozGIxFXEaXewHCXoRK5XHcJOU8oUk5G22AbS6HkvN
4fmSFZYigGrTVsLphalhU1AhXameSRoB1fMsIbcmgvU6OIDgRjNAA8nT0f26LLg6
7SrlNPx4dkJJ78OnrmbqRmXxKuxbpzpmkq6AzslfGTfvkbmeD0Jd7fLg8PT6e23F
JqmmicGtVV8BcmxhzCZfkD2hhfoEt8yMvzyJ9VshTjheuudtoiQGEoq7fMyrMkfR
2c247RmurngVqlsgxT5BY8aKq2bYV3sxBdSZ1A7ugaAxBV7AnxuL+duKmARm4t+W
8czDCGFikjEB0rV3gtqgI7HHKa/1xGJ+Uhzta0PzN/2hp47VfxG7yeoma8n/bRcm
gcWFQ1WFo5/5QGyB9TVN4hrOyD5Eeu71paFETRx123H2X/PcPtclGEOT7HkOnSjZ
KBoKogstteP4tkLdpJFHJs6FA+0DTXDbJu4qbdIIxgf8IHZ12RZao64hAO0VRW9e
LrLn0QPGAKmgfD0PsYN8IMUecO/OGzqZRmyFS12Qqt2W4+Xnvczy4Z0H8eXSSo/9
HciK0J7wshSH3ZeFIJt9JKpX5yhqoIzi+XsmWKixTfxa7w5CifD5EogOcbVBf4eT
osWJ97uNRYyFzdoLzlnq6br7fMnHtXpMox34j5AiDR2QloWkj1MdhAmYnkHmFAPG
M08IJsAC9eTugaufaaMAn0L9sAp52MOAkybXWjYEjPvB4Y49OCLo3X5U/YYy6Qag
JwJEls+LcCRFcMDQCsNfcVXKdGSxdd99tDfcYkH3X4xiCFetSBjNKkOFRR9Ua+Io
hVQFPpxk6VyFngqMsSqnrC1QktsyfH+O+YhtVzZAyaCfQzJbmeVfnmbCM2w9r+oM
WpeDjGBs187nnk4EZyhIkE/nI09uMZWGrfc3zhiAAjaeluzfWvry2RJusmyD06Th
wUrdT/53w+svxP7p+nGxg4f4a3iOrtWtvmkNq/W/bv/Ht3E2nsu0mWiKG6ZVl8js
e/XHAg/QmBhkl+yzIS2CVA9OE7NC9N7Jc4dbduZkL65mENjYeUcr9BvA5TW/Vivg
MQU9VIYLI1ncO0bH4l7hqO+N26FZysljj/Ltv57w90XVxlD8y41YXVpa9ZT+pRSd
Jb5WokWopCR8k3HJZovx/CIVS8sgxEi6dhutIsaYuRbbZSlWFVLIXzoZqSB3C4ww
qhMlr4tRjaMoQciJgjzgCRbPuMExK5d3dFPtsGUYCIJEEmXMhDfHxS7ZdY3E9+pP
qw+lyC2+dNolwO+8a6NXCFEemeCba92NeVxtKJTyneUordTHONndeQKvW0k2cYbu
Iu+5Ishuy6fa1nUqJJnwwHyi097Ix9zASV0Lk/VERQzmw/G4UT0pWj67mn5qtUaA
TzFRt0rodQ83aLZCgXsKqTHIDyvPvIWzn0+HQIR5R35MpoBiRC0DKxtoARiwEsmi
fX3oKWqmiNSR8HJrAekAfk9S+rl3IMKV7e6rdvo1mRNNtaUdilXxZ5EAMGy0RpbB
ufBIpL/f1kbXt40xpi5oOmF2B1uBdsLRUW2TIts+uEZxUMSGzxQOvb1TxkK/P7hR
luxPnx2HKTkbW8qUdukk69pgxpKY3h6BsBXbG1b7GPz9vwZKPGpFZDreKiCGeKqx
DmgW6HHhSyqCdQJS39nlYtFsAZRNp6Bv3CSbSqta8EPf4RInVIDhv7TwNpIGkW63
GyQXf/dqpqTFEU6+O4M04odKfAtAwaBRTxcSG10yQ3SPfdKlz51RzKF0Y7V9QzsD
5M6x9xxPnNQ5tkKLml/Gbrk18tiBgBGLBgtAl0I5TlSYGKyTbcerNIqaJrylq7zc
fQkJwbLrzjBtO4hgw1JS4H3ijdEzRdSVVdCWhtSaVx684t1uzhRMgrhusCyOrGmJ
h5Jif0j7XjIzWmmeBT7KIDNHnXjjSQpACCDqJv77C7bAVbzHkk+gmzCL1gaTA9Q8
NYXx4zuJ8wlJjp0kh9Og+38eV03EFZPeIHB2TrzoAt2YN60P0/3U4e6VJHZlQOJK
8UPkJovaDxc5i1DTqDJgDSjWhTVYMnV6OsTOuEBTpWkRjwt73QrnuFbSHRNkOp1p
Vl8CsxVTtb5Umv6AYN7tEU/3LZwTnaAnYt6FMcDZfrd8nWUJ6eQuiRKtxVJ9nq45
DJzCCuZKxo/3rFGEGPFJXPTSRfaLhWt+WUjJETjvZwEpghfm2v0lB6bmoUjyyDbL
oRFRcawAysxOJRla6YMdhQLutbkSqUXUPR6SXpmrTuqKh3/8Z7LiALvBsARfJ/wH
w41KQjh03uKIfEg/iTE+dMW60A1/QeRzrsQcyuor3H8lEWWH32GAEhluQI4xHYEt
ClwsFH6qj9hsHdRL+uKq+LuOJIewvP/2Ssexnmuw4KbV/ZJefd1Ifo7J9y9izmr/
iAikaaG2W6tmNZSX+qc3aKjBSo5Ccpp/Hu8Zn4Swa/4xtNlPDZKddBZSOZgcoUtB
CINbF2mQQ2k/QMSEUzB4oVt+AzdcAOMR39DQ+Wq8Tc+QRl1IMF7694pJcqS0UaTB
qMnn8UZtQsLn9ZIulTsRZ7hB3MmaOiDtc/gTyeO067K36vUxhc7qFFP19O0zAO2Y
wKypqg3K2P8a8iUdslNuHD0f7mp6oFCqZ/o89Vq4bE38P6H9NU18injSIM5Ep5gq
SaoG2WP5c/+JGd8PuF+TYpVZzeFKNJ9R473FA/XMyTresSFKfGSenKI5AHBlh4Ll
zPrKN5I0iFJ8dnyrlci17/XZczQj4Raf8amC0AvEMFGYtUUDdfNBAsOtHrdlTcuA
WpayDFPP6xKWEWmBFU8ABCT8JFJ8yMDyFXtcYpbQJ4p65XbZMDhw2Jz6XULZGZjw
n3dMTcNTNGgY9+ZYoWa3wT/4tSDUmlV+ZaPLS4ohEBC0ya62LdBxSCIpyM//+QLX
QdJMgOYrO41RzAfJDADIhRNUxLcpGKsUHeomcllPlbzTjR6ytJKIKig3ixhRnEt0
eP2BKKsznUDIsJX7L9B8wy+yJz/aj+cuFNp3cyfz9xY2nr8Z2udZz2X8b5un2H2/
a8gyakeITc+1tdLSajVOUpRcXrwOu+Q4M/lGu+3ihmw8UAbFiL6zYJJszy9tpOJ9
r2u0t8oyfIHmv9e+GoJo3uR6/+Iy1tE2LU+guzDdCq2I7t78Il3crmQzGGIlfLpN
K3f37df1+A3C6bhdhUHu+S3spbIl9FMjuGiltbQ7Ph/HYRY1+pTBT37A9qc5FJ9B
+qagrcwwQwWTaJLLGfx74upMUDxDROx/JGhZvnxmd/U7NSK5ROrOLl6ErBCvb0iW
r57mK7osB42hKbN6hi9j7BS6ApiPs1R/ZYQBk/MA3bq/w24n2XdZzu/zRS16n6nN
Q9OkWBRbFcLBoiO49rHI5h4XKykmtwdCJeNHwWlxLEphxDAd+zLXki8MLz3VOmdx
YG02lpcOgzUgLQXqzsGqI9+6LU6SZOK8RuHdxOWYSpHuQh7jdychsoTOFVcUAG2u
FH0+h+h5V5u8y7npgB5v9Z2A02AtBa3DfWWxPolLhRA9w0Dk1rlp0J3UdeieDhkw
pxFbbYyoUjGoyyAJT60RWqDyme6S2cfccAAaPMaEdNHnayqA1oz93bA5JFXnS3TP
tePbWl8VOyFytYVkWLR35Iy46hKBPenBdPuGsi3tDWVXdHjQdKMp4CQEYN7XvKxA
eZyYwyHaF8zxEbdaYvM9yuKb14DVErZgrkWTOZFOrbWvKpbjIlxZMOi08iu8JsD4
JnhpDwP01fUkZU83vjXPx2Yf6ycTZbDh3zCFKOezl7oXWOq9tjDo7TZWIipGShji
X6oNhxdjYdq6J7LSw2WrF6AI3DduvKnujh6Q/p1XsEGbGgdedZwk/aEAS7rzh9uR
AgWBPRkWv3E9XOnqOXsZVbtfJQdjbsccUbG3ybwGoXmBQ+5VUrb/gFjP4RP1w4kj
+dudpX+fpAsZWPPnMHlG1EO+ttQ98PJY9Bd7teFF0SkRMePMTq5MlvTzJksojGyt
NupJ8JYT2XzY/GRFE30/ebOCvkJ2Gvs/RL0sKfNVFM4AcjuhRRNto/yZYUkyYGLJ
1emPdWWwokMi8CGy/SjoN6yOlTN8hgbLu0F56pIaOXp2vbN15o3JrfFlzzNnxO4N
1rqRr9Ydj/qmLMlWXcfd/NseAiyWYtkoJg6mMmDP8/FyyYN7rUOaoCbhs+5/rnb8
OJsMDwixAxikhlIahheNYOj79mVPNiSNuW/B3ciWwHfFa8QAIQRLw87nFJBZX6WX
laUh7M/a+ATcmUuUvZSIbmSJLb+8c/3E3pSkcS06LXrbvpqzVbpf6/++pAfRu0fl
P45qoR8d5Tz53oS51l6gJ7G8gOrh6IpNUpaIs3jUVtMA4LPRH4Wj4RoEO92pkmT8
1WqdCkJx07P5lwUSpfeHaPWXYBPSaLZOXNkTZMKVg7Bl76xwvnHF1Yi192H1RTMo
+XTfaE3wiOzN7n2W3ULPcU3uKB9zFvhMUDobZ3lllO66Jw0g43jZXgKbEVR4ZrAp
YBu7rUUe72STdejDb6ktbfCbL1wn/tJl+R+Q3oNeggh9mDLK0Xn5Qp3WJw8Zg70G
2fM8g7nsYwfToenPQVXV68mmfhp4shmDOqp11TnD1Nj0Vrx5RvKoll+vsrYlJsTP
Aapv0BoPpnWLbnCxl+K4xGQRRAwb7kHLnXk/074VbnAreu4xlh9d7UF7W+D2WUnU
zhSa3vCQJFzZfNlwf8JjM3UsQu4+535U9wHbwYxeLJAluWFAH1o19mCTmiiDd+HE
jbgYFLGdNSodiVHIvNVBDpGUNK5thLr0SRn49Jt7l0iaDMN4ivIH3YUbp9HIwTab
WAX4nCOLfEdQA93eP5qYtMxWfwGRtvuiyKOHWF8aHpqdEqabZ1ItOqwei5KL80sf
H7tZtd1yrenlv8R0JJ37TXMlr2VB7aLYFletridBBlq8LbI15hIEqsxDjwF5Wa8c
PtTtFJIhtEBnF1Rmg/TG+LcHZyRddbehj3TCO7F9fMi7iFThnkHHf/8pbEAQYHwY
OO4oHr504LBN7wIoQ/tX66z/UpijOOZtZxMdLCUUcZDy1vNt5Nj9Xr6n5E6aApnr
d3+2qLJ/uSbHPYIA1NNeB6P1bD6lLFOWiC/xfwM/Q+OHh2eBmntLjPfYtNCgiXno
dlRK70JIEOTa43mC3ygyzIzMvHvnRtc4jp81JjkP6MH95Fz/WBfJSuSCK+V9On18
O75X69uWDFII8Nj/cI5QQapHSUEPOfTyNxiKIk7cAVmo3cTx72NJ/Hy5CXsK4U0v
zcKxpbuDILFTOKn0lk4bO6Vl1AT5RdRY10eZkPPGNmnr+eWdAYYj3JilVpqWbK26
j8nPdN8ycATc+lZdR91kULuYiXs/GSXS0d7GUuWhb0XWRdyFoDXj0rEAMYwgbTUw
klOd7pEAjNiwVrUyl5Rv5dV9+MosgmP4j7Cxb1HIPfH2EwLQNbRlsCVChd0wKyAk
JOW5K3yZtOohCBqRjnNzLQdO9L6JOiSin/iujOHg8ef07PNkGG/QLVWliXyAkwzi
FPfZDTROVRnP+FGM0kQyBqonXq7vz60bkyBQMfaEKq83B88VqF6hXus4UyJSaWml
0BbSAiI/XnCtM3Jyy2dG1zEbyyljD0VdJ/nKBPXsiisDdcXfKJIA80iDn5Rp+Hho
waAIOVILI5dqbjGJ37pX3BmXVMdM7kEIbUP8zJlTlL4ZvK9LdqSCHKEdnDc9C6I3
7kgXd+pzZgo6j9sGDxC9zELGdthZOBFeDm2vLlll2CoANVHcsWFzpzhqgoH70z33
JwvjpfNgJeMnmWLqJswMq4Rwp70vWB3ttYZf9DyXMnqrO+VmqD7oAOi3+x/BZ3at
za5ELJMH/MGckZTcWZ20uCRLLLM6IpB/qg6HKt/E9PsCnb0MEIXQSavzEHhRG+DS
g0uPL5Z62ZJ1e+N+oe9XUefm2hNiozDYZatsGlhOQFMpRFnLBAKC7/UwBMoAC0Ao
JvzlxcTz9he0JU7ILaBW8KJOJhBRsEOOdTlqVxCWg2QGEGOaZidsSQmiSTJ0c4Pr
QN8nPNiFrj9OR6sB4esZHYPdf74JCKeMMNBts3IDrh9PtXfeN8Ujgimn0WFNIVRk
oHOu7VWV74rJoiUx305EIq0X17VS8kuLcQU7wMDxCr2sf5dE2p7Pwqg+RndVWJ9X
UqrGr5NRTKwwE4XA5I3xJRO/wU0cFS7x5IucwDaPC0Df+II8dzsG78eFicizENAW
F+fXAIIoTUiIEQZVfCSARh8d+gqLDufewg5L5rPue+e7OD3ssQRO3R6qbXkXaFRf
2vmiHJg4FEmBu7I2s2lPOw9h3JLjuYfKNzS7NPcpwpiuwktMK/TCkiaD9K+9SPWW
KAjcwPmGS2pkTyK/7Hs0oNTXkXfPy30+MfJmhuwJSLst6VJqxhjV+dQ+PU2gGghz
CqES/vI6KhMNF3R+x8zrqw2qiyIV8iy6R6q8rDXp9y6+cnM9jyvjKeHvM92gietF
NHNgwP32btPixAhWreCipQ+eI4HywmYmUEKftmSIGVK8Fi9SBS5JtjCutI7SubRP
13PY6w2dMGD0QNfZYwrWMij0F+OLiMOWX+NPM4a51dq/wBVbLU6RFw27JOa5WTOo
s+QVKOV5rfVSBTXyX3cvoNBRHS802VcVS17lfz6DI12lvWzPG6bVw2nHDMtxLQw5
87QPAJUsXBbbGD0dexIgyVXz6CZX6C2F7Rhc96kcsynrRkecojHZygqyYFULK1ux
/OVeU5RibvEy1wHMiQjfSNcYwOZTJcBnyYHnnV7fEPRwnk0piemkuTqwXYRRFoO5
qlMzR3P7fb/XlFtIibsSTKTG8SYK97D9ZcQ88gyESFSwUhOlOoAb2scrsZ2bI/Ib
9euLNBOSV4ng39e4Gyw2caWq0wAutow2T3ovL0kz/3W2W/QmL15h7HIVLRE4kJXd
D8XuN/3Mx3PZy1QotnTahEM9NEMDNMFwn8SEVkMUfSqW0zPME6rFGgOAU6o9BRTs
SH9u3tRBm1s+4QeMVLKUwpwgf7s8ickzdENBImGnjL3NHPjEicvcqGHACDQtpQhW
cRtirDktHuqtp+5GVq48ZPz6EK2/BPEn4ubIqvlGBKy/jMbZNeNARCUbaLOm17qf
QeJug+jN687kQhk+xIKWMQP3vQA0GMosItM28vS+oaJ3IQ0+Acx+eGPggNzdRCmg
Igrr3q43uNiI4VBSO+ZK8BAkuRQO7jbHjJARddJk5V0wSh/Jwoucllp5fMhR+xlr
NFx4gRg5dZA7R+E+UkcEvAIxarisCb47oeKAScbPUzDzpWzw5Lb6sIXdOjlrcqOj
QhjVQEpf1i0lZDPXCh6Sbfr4tmoEX5IL/CdReFHTLhhRbc0MT4bv05d5as0VyIhU
CoSj10EVQe3Lk9Sg+y7JKV7K9o/ZtH3ba2cBSrpwGZQFGS6w3io7Zi3N+n3OOCBY
Nw6H9trvk1UWmw6EC1iR9IiAN7oACoFTJVm5MpNdP/62EsQFqoXmjVHRpGAF7yPm
e2+arNcDE8Yzhu3Yn4oS+wKbyMruh3vypFJaVUAe79m8L10jxwn0rvm0D5fBSsN/
VPJ7duS+XQiQGwmtvcteoywB0+LljlfxW/w8ypxq8ekkfbUVmtQxim0iEtIA6XNm
RjYpHGx51j883YlxNEvsYP2Wh9Bzcxc1jYodWBCaAtErjkyGQoRxpM2HZXejw5+f
mBoOXbwr4rhouD0rnvT7HP6PQ4wlF8GOupa5W6tDO0F4vTpN/024C3dr3Ue9zPRF
Qe/PI+ROCrm0IbZxdqHpXIE8FpLveEbNA8s3F9PDFbutpHCOIvKG7nb0X3k4/Rkd
H/ZUKGdOrtQF2AVPkkAtakt2SM7k6Sz6tdEwIno1hWrn1d3wchWvk5W7VX3oBMeE
B4ihcAK9AdsHxHbS3kcEhzzjVMA1lf454rTIveqJxrmWyp0vfW4ETbOfUZjXFj1e
/MI6Lhz2T9BERaJHitOCvjwa7a6e3Q6qBZdeYq/L356qLtjkO1S7DgeFVkjPuK5+
C1Xx7lFVjDLoa4YDNuTF2/IKvkm4g/RiEZhMG1JjTT7uKgkAfMhX7xomAKHvtZCb
56Hw1kZzqmB6ZfD69WMHPEtI+qodM7iX7NUksdyHQuBhFP54aFmUNik/Hfodzy0R
sCJLS0ZiINVWSQG/fWHOefeTFwfGF7Ch3xKVxvb9rqHg40T7j5MGpFUJdS1yTgLA
TufVgKij1pdHRyk7ZLnSf0vvKfb0EOBk9UVDHOqKs0ogHXs+x1cSsd+Trh/rMQv5
F1OM4edVhpJTkv9/EeOHzgo6r7xjALKaJSePYrZhn/Rh09z3sofZ4GbOpwhXgNSp
sjfmykIpZigfJzmQNYPHaUtXMotBigcHHd4NmJMXWsWMHeDkymyjpxSvT6Ckx5jS
Lth2qMpZKHGrM4m+MXOmiA6BsRAr35hCEdyQWrLETLsJuu0FEz6U22KtOcoeW3fm
J1VcfED2Jrhip1sPFYM1W4CpkTntem31C7t4BiTbgIXpe2RIquvw6xDAAPnf7kUA
hQsd+FG99izLigqKQlZz/LoUNHEpkYvBBxp7Yn1RCaGK5pZ/IRv1QtQVFPBIh5Nn
I/JEkzmfnhp/c3yPQgroVTJ1nkx/WJKlqbXfRWFTTSo1rmewWEFcspQI/EBvbXmE
TfVULB62PwNJJ+r5/F8c0cjHv6ZMC3DEc/wTyLnAQpYgKiZJ3/FMU4NDPctCp/y8
hkwOsZuoqHUWIzdJ2OLundOvS66JLJi/5uYlqrCdCwQPE936vSSmHQj2wXLY/+s8
9yqEQ/46NVIR5xU119tFCJJIvfSsgjGhymQ1En59kl7ni0FrplrjnqI1nzz4Q2z0
LHSzFgrgAxBj/yZFHb90HRbbJOi50RNRiDHNKLVBYgN4m8B29I646YUZNfiUEohF
R1xVXBm96bV1bMywGjmlLy+264sXdyi0qsQXxzmJ8JHffVPUTfbpQh/0RFw9xZaB
Su63znY1w8qbRsnStOavRzXtXhktOXDfc7HjFOJtKT2DoO2oa+lL5rRaFC7AaNfB
MAig4gBLpdod/gVVr3HUHLYZh0vIlZSuLu+bjiSS3QEw+eVmAEmPkjCp+xDhV7z0
VgEMX0QfI6UsDUA0cbBdCO+8Fb7llA4y0iIwFUrOnd4vU0KlqiXbMszAQH670dHN
DHlowf99NDkKtEvk1m3ddMuZo0fMZniQLeDytxcCCB/0acwZxAnz0vybsogLrmxM
vZNQMnct4Je5Wsc6J9LH2dYPK9QUSPasl7ZZi7W5IH3gkLBShB8iTXS2eCphlCAu
wXFfjG5LV/mactWuO1lgWG/rbRs9qWF8vdJNGX5+URc6AhuriEahg9xxXEEm9nvV
s+R+kqh4/iWVrf5EM4zerSuHWIHR5xwgrYiTjk09zTI8ZEaXztyEmy2NH91mrO+/
1fnU1voBPdSDaNQWTuUJ+Q2CLh8x85ShM3H+ajVUWz7VW+vOK7HFba4w814dFEQx
7mC/Ou5ZuMKSb4zynYXgWJKamnwqKp04pVamS6Cv9CCu/U80YXAiaQK6MSSlwZ0/
6PXM80XluBsDpoHlTXoqwKF/7KZN0ddrw/vPONmGlVAMrpF0ucT0P+IWTlhvfZwc
vr9G+kN06MKa90dEPsZmLdxmS8j0oRto4rmH+Nc2W1T2WQ0fnkagcWR7rUwNZMFE
kq2YMZPR0R9TeQwi805K5JW0bV3h4EvFpM2He3IvlOucprlgpoHbeUtFPlrw1a+A
yxaaEyXj3OHzpNY53SGyrXJDWyNirLHClmJPZJNM+8ESIDFiAdTcYMv2ysHxWEWA
yexc22f5OrKRTJhJQvN9+bOzUoDGzbk8xLRPhjfI6otgo+COmR+PvuCtFyISubne
AQL+ZNw26OyEPEYYAAsOtZsEJsoI3+PaUr4A3RHAFXnReOvlP58xM+ohf1lATWiD
Nwp56oqkDKMvxQpdnucfKWDx4zdpMu2RIpkAvcVEjfC9aypBwxr4WWLJLHL7UWB5
9vVUVEelJdJ899LCu/NYnqM5h3xb6nkgUYyjqGnNGccDIhbti4dQrW9d1/k3iR+w
EAXQPXUWlHqsoqRUNy+pjoCcVNvLNK/7W7gVHgQyt+a3ZiMzm0cSY2LVCz7DXj4X
T94+ChXMX2dYgQsQW/vFa+Dk4z8dvGg09goIeWxfiV8/xW587M/MiKGG1BCTks22
ut7pQrN/XGBgl83jZ1PI9q0d/zDYYpaV6f71vbVanxoZgv5Fw4/rhwk2O+rX6Idd
KU/87h5MZLx5K+Ca9OTyusGsxijYG27L0YJDw3EPzs4yvjuJYGkohL5t6cLncI4l
rgrOOxXmrjnbBKHb+1tfYX7vuG7h0WAFwvGPYLcnsyUwDl1GVOqyCUfp0ykuRHA1
M36mPVrdzo9UIJXO4tQjLtfblBOLHSlLWlDLEAy8pX+lu1z3S0QXz7+VkwDORPFN
0/dAG2YGT8gpzd5snwwwou7u/raNCUVHcH++CbJWIOMJD+4coCQcYrfd14N9+owV
mENGZlhKbChibIlCPmcqYfAfRNr1r1F5c+GgOY39OMVpkPU2OX/eEtEC+t6Nj2cq
WIyl5yCqdoR8tgCqhcfU0dwJ2DwXdG+lm5FXwpSHnCBVYGyRqlon54osVVdVL+Yo
LYaILfHTYGohUJkB/mglIQJv57SpP7SwPL44eIrN/Ft+p874+/25wK0+e7zyowoe
2yB6v176QtI8i+bYA7MIry/v0HfQxYtnaSs61A/950J/tJSMpUqPO96dm3yIS1fr
A7w5r/ZHZmU+W8+xA8Asr2xUNCfh+7hkySvuDGle/osydIBMgfAeERsI6wwB1dF1
keqYtCz7S/FkydGF/7YsllGp/2Lcju0hT0rY30x4s44ci2FFBowfxl5KCzKf5Vaf
r0EdDfDdkeEUEOSifT48NmSIljGsaZdNX2Trs/r9GMsHiY8Fycj5VypvkbOA7U8i
07TRqXCfgFlbSUgF2BsaFYqrxouwOa8aNw8G/k4TxSnhnveuSVHu+Y458hg5rTzl
wcTCRwpFGTOqp9VUOQ+nnzG7AOWxYQugFpY6R3gaf/dxB6q6nIcyR+/q0tH/TmBR
bfZz3if2Q/UzmlbckShIrBOC4R4OsdP+SPzvbPW4R7stJy303MCg2PvYS606AvhU
ZxUGflqGZHXsoFvXgO01FJ8B4V6thsblKkuu1VUd0uY3KFnTvrczBvnuuyJ9YB9q
hfKyN7hebpojBQAUy63T4XcnbkmjJBiY5KPrQ9op5Xj04b1ezxkPoDVk0vJNwoOC
G5Vdbw7UWUaF86jZgX05v/8TQoiJPrtDDflUzMl+LcQ6mRUpgsqt+4a2ZHlOs9JO
YFvgR0YNUc2jBNBXgyn/s0UsvIMyPNaopw3svTaScUVEmawq2ysweUejNTuEsxaD
DhUQjfSOjm7LlDHGQuw006PB+QVz9PiPBPAIf3eJypxY74Vge3LG+PrcJi9o13mC
H7Rv1tAa4jZzo16AQiD1dU42s5KD/0mRX6+6rfEz2FMPhKnOPHEOjOgaYs+sKPPA
Yy8PgylrJitkVW7J1KUnWJd1Kivu+XucS7NfVTwApV0zGU+rgIFLiB99S+rn0ERc
p8FH38NozdLIsPKHw/XNsaE1rxw3eyrB63zI/J00IpN50tohS1XoVr7ATebb+YM8
vJ3wIXVkh9ZwltMjwbIeQOSV55KCZyu12+K/TucCiDvsoYpzd7jAVqvk1pUhv2oU
c+lpQQZu+in5if4DyUixdus8fYrgV0f1wia5XtQUkMR+qlJPisq4v/jeq+DP8c0j
xKiQMC+7O9tkAP4wfrmno28adURIfO0auMpdz6Lmf7wUvXd4MGxV7diyWxcio18g
D4H/JJqosIVcBwSNazzp5ljonP6pqUd3QiQUXYl6sJSLC2CiQk3EmyEAfhMkF/Jr
maMs/53BgP3OPwsDbWfBvgsTUkx25+Xe0Gmwe2SOAJ+EQEZ8tIj9nddU3w78eFJy
96haELyvzcsXiQXqrcChitsL5Y1kTwb2Y9pADNKMeN86D2IX5/GEHCMgVF8sItrD
S1Kwn6ngYyOR6K1DALZlxKuWJfoFUCeDyvLYHigXeE59k9f4j1+zGGcVJrA8cX+y
21Pt08mTJjgvI4uSkQ6Ken5bxApZC4v7l+LxX4yUx0nWG7Bb+ggNlGseZYyTVj2g
dwyBvqHPBgi/xsmhCK3qE8qIxUPL32sh5HczAkl9dusTSKMb7K2s0me87blTIkwN
pWDrScLMjaTDC7jlpkpr0RJyPD0o3V3LmHRmo9c5BUUPIdz1zXZqXM2cZHSxGXYU
DA9EoOniWzTupXwh9NmDoKDf4dQPMNMUV8727BCGi/qqdjdv9pxz+Mh9xhr4Vh0Y
H/z4i+PNgTw/HcL1JAyjJvn2Cka81b3Al6HAA+Z1/UaRhz6O9QDELfQ3yzZ30i7D
QcMK6A6PTmcgKoOSUgGd4JIpRe5V5+tbiQZJ9BEU9UgZgyzb1j5GDm/RQr0dbUml
m3kzAztguyQ09haympq1OqGFYYW/wxmO5Fvx5rlWudnUlxcpCOvoMu9zgdzKe5Yr
KY4z4WvHzIt3qVV5AKNLBYfyguLItrIZEtSUy2x1KtvRBIxZU9dOOP2hOqJmR8B/
k6Ujkr6TrVDqVwIRAE5X2ItcPEcbQcWvYUZRG/RZkCiH/qJ6/OpChuQacyxVwnbs
UyrHVJRIUdNb5L47OurHqguq9EueZh7fkyUs/SNaVGgTtvLnZ85wLILSl2rhWTfK
MK3eQ+ZpsQvFW0SFIriH8EW4VJ3MnMXOOy8GAVe2DEnCgxPvohjLeUGCVUU7woGx
x9TzyOoeyjD8wrHM/zM0IoLqvRy9lpzXxrQoLzOIHLnqS9qvOTyDZUWZPOmz1b1U
i65HYXkkf7uYWlFgSSwrEGNAg8KsyQ+0ph/GqcIo+CgJoNUyrMvZzvopvXNK6Ofr
x4b1eHAEIdsu/NP7ooNtQlidfNIWshTXpyQG5pWFwc5ixeWjjQvFjPBjzgsE4Upf
MzIwI2GJH0vEPAqFMAE3Yl09cRS5zd4BTU3OiF+0DofJPia+gbP70yTU+DLu+hk+
bejoh0dXl5S6GKw2kU1lwznDG8EyahPc1+NdtFLb3yN8Wl7wIz0R4MqI9PPP+0Lb
ygblOXBTjL3XEkIy603FlOGg6y3tB7FzizXyzXDF8ZoyWNZTZxXVJjldXIkGPOPx
jzctsKmMJaqkEBPfi5jFAfMREuB0LcC3b9NYvTPSJVtbQPOSP/kOuFxA/PUTdCC8
xx6sKDnK2RGBkVaqnK3KkXzDk4rFNY66xjL0t6Il7XIx3Kc9Fzdr99ZW6KVkEX5t
bJE53zvW4M4jplObtztwPWVdG0XHi/LGJnS/bOFIIjTU2x7mKnIhN49UZKmNcMDC
s20qYyyv7Yf0uDMD0/fnVkcBKiPmspi6O7DcPDsS7kdqjXpo+0/yPuaORSV38K8Z
pxkgfn6rUMztElHhtDnHDXORo/pyKOeDbEiwl0samOxRS/Ah/VfOVGAR9/gdgxMG
fFVHgi58hMiJPfF5yIYQL4eVwmatLxKrYDLhl1SPjYmZI/jZLtB3UBs0SHJtUdjT
oRCTjylbhvdVxJ8r2ns72kwIwRIAE5ZptS+TTHK6hmsRRkIVX1GtYGwlfbIpV93c
yrlsFMukBclNUkFUwXarc8KCeW8crPMgdVX/yQZF0piMBPsD3DIDEOzq6GZ4/ckA
/GLvxjx9mYLGvimftqO0yOXdMOXjGKd0BO8gcKHmovLESu8HS7OfIihbsVsE0MxP
JPniCrx5noUt893UpyR9j27ih1r5wFPfbg73GXtbZaUvmMolUkB72JDj2QhROM8w
s2DQcWuHe/c+p0J84hnDyBgv5df5Tk9+RYhL4EaZ7nnEuCa3LahE2swoD7S2T//q
0QvVYsQZBCi2wms7EPlsG0Bdde//fXlG3U7kk64StMBRt4XEMdIcTsLPvet3sjTL
hWZKmhhhHmd/okkbK1YbXI52RV1Vboo33Z89TvTNQ4sd6a3WcL7JoZ3G5P4hskPv
cqHfaeHb3gf8bk8ywr5fZCJXMkrt2OKdS1upjGYlQzCEfMXDZW8N3Vhc87hyFEus
DpNmP/5uv2b001pX9NXzgfaTfnwKkkaVKutYuIhAec/VukJqw4FatGrKOrn41n1w
SpthaQD0hzNGGbptnYiNgKENHPAqwww0kr7Zr3Ey3AdI3zTYMvDvdse3b4+jr6WY
wCJZ7Fn8ND6rHonxZpLwClfQpMfJAddfnTIIc1GNW+QhC6r6+rEa9y/RxH5nP7FK
wDznKMMyY198zz7myyZNp2me8lh5P02lT5jhvdeEepSX7NOm6DFNXh6PxjjJCrXT
r9xMdo8GAmhnfDM0CEVeqwqKEyrbzaQTV7VlDfJrw8yuoZx7jS4GbY0XEZdwXueo
2/lxHPejwXlkquBCmxyPtiLjzlmDylrHfE3cH5xcfhB8qm1CqKfgVg0Cw4+YWZpS
6h39iJ6IjULsdaXLlBWIE9bbCY5DeRmHworzu1M1cj6FJcWdvcPIFFHblO5KF1Xy
MyjWnekA80EUv+JNKngXpL+V3mRUntUVAT9ODSIbzW4+nDxftMiL+skSI7zSOkJT
UpuQrNqbyUPDbgrzjtVpfb/fReUbPhEjRk0FoXlJ149bjj4+2imsA0vXHmxnlVe6
C04FjmFsDGb/zovOw4XN7wMO+2HEY2t+FQ5F350K43mIMj2KFm/B5jyZVrMkncCF
CfURtiXZJyrUoSrTtn+/UmNM0os7XuW2MGyMgAbcJXISil6NWhaOrjXN396PsvVC
OZqKcrAcpfRAGAmwfCHLCENG7VkpkIBUTd+grdthA7DaJvnOpOqTaMYLUidCO1X+
f69ozDnLMXhh9Zji34p8eaweH3H348ZAInJRQRiBAbKM5KFxtrYOa5cg558WFE3F
15AulcWhDcepv5fStxbOXM2lI3K7x6Z5dXy/ZWe8QR7YFXyBVDK6FakfG99UzFzu
f7rm4XcXc5RjaEHx7NMo8CATsqnA7pnwXwvDFC13W7a969yh2i+81RLEQ3UnFlaB
82e03T/VzOjGTXVGaYroXJGxJzGPoFCrx3123h/+1nxKavRXBpJr/XV0HL4Xzjtf
xes+/DFI9Shi1RqYqVNT/aIEWBw1vKpu2Q71XxOc99yeBXE0YXq0S9IdvhBKP2Qx
Tw5S2pUwTjn6kBPTKEjgy8orqCg96OnuXZgD14M/0uYGpoRgWExzyAZYU3pxiYIa
TnPyQFDTr2wHqy8krQyc1e3U87XUOftEZ4lw5Oz8okXAmVlU3P6SXwGXd8yXM82l
QH5KmlDOLTXdrfVVONwpFhxjQeB2vxGSl8y9fSc0fBfzueYE+5El8rLC/fz/BIYG
GGkz1HrkcOlq1OBbBa7C+5GYeecxgyTr3+t3ax6B6JGanVViddDOeaJSlZGr9pBC
XXngty6U5a5kR4mO0jEnw4wEYpu9uYpS214+d+aDaAtEKANpQXuPUfsyRqPPpRU0
R3jjZhOTxykyze33eMXEUbhfdSSNgqPALfwXhpjUZ3nXDynxITSL4g45qNC98KsL
WsJSmIv3NK6EU1HsXUKX664tkWPmDa4InS3SpKpX7THJ2rLZvD8SD+H1bMAQep/7
SeIwW1Sfn3Cj1ZYT9030grHmJj4G2/EylkjJT6SPJGi2DZzQTG8nIPzucHhIENJe
ysYB99GW3e7zL2PW+hdiVsxIdqoiU4HGeQk4xiSmZB1Cu0xCa5cA5u0UF4gnTXWO
XRCpNETGDacGszfVms3EskwpItVLyeZLyJWSg2gqiucwuPj6yBcyCopev+n9MZ2Z
GdQMlmrA0ZZ/7mcxerTWsa6VmJVSOHmuLZyCtNTfaGeGbmELgRVQ/0hqyFyr2xAF
aXbycCrfSK6XEkGRzj9f7m++3VARffHDlf/FfMZOHmRO456k3SnyHI/CjhGLCIsI
ppeDYPckwjMWmtTrqKRP6eP89nJtVOcuXilajsY5FhBSJQMkaxkQ+v7LeQDsj6ra
QK4mOqFCctixgPTYPRpiCein9DD7WER7cetdBK6LBAVZZAkLAN4dHp2IaimMpmVE
UcCPHANVP/4ymU25C0H+p1hbgapw6ZOl0DIBTqsdxmQo0YLRn3KCbLKAVYhPJK/7
CLaskz8b2F9D87MqO39R515C1efLlPdREpUaXdtm0GOsGi9pANGaoVxDG7G2T7yk
xVHrVOPsU8kwO2xKiOaL5bt29L9h8trlCqxQHMYJ2FKK9hhISetaFznQNx4pB9LK
3JGtxOieys24fW67z3uB6mwcxgGST+IinLyekYXq5Qnf1iiX+Ua+KcFPNiZs9YPb
/A6+VF/sOaTuwGP1aPomkJSDVqFndllanJlzqvG6TmFrNh4i0Av9owr52lFg3Lst
WXxU0bE/gMRq/C96fdsLi74XoDC9a1V9SPT7/R5pu4TERSJ8Q8reANPo3ApwR/dN
IUldFgDcnuCFfz9q81QJJZoEmJq443BK6tHcQ9/sGMcpSCnMwr4Z7CqwAXkhSs+f
zZ2jM3kY8TcXpF/V38CO7bfF0UGoe1hmhLvnviQEJaUF3l5Af1MIn1e3VWx77WcB
INio1M9R1FNMnGVBAFPrAZwKMOqA/dtsVXzPUDKaj126ieZiW9O71cfNoWqSLm9P
tpj47Ku0O5Tn7YUVzU2U0cpyFosdzIg9xIYnDe4wN7NdjMJlfxr3qUPtSX6PCbja
W3HFYCl2xPZplTKYwGDidYfGL9ovaKwKVDO2aKOenThYx2nyk36d/tzdoL3d3Qjb
XIhLGzpkPbSvmUtInjSy3VcZzcdMVR9sSY33cCGjyGXVkcJaShMnWc3v2+oMMrPq
WzEOgqJiJrXMb8K7b1Mj0r4w/AIySlAvhWFiPpNBtLyl1OXRklC8q0jlLeuiDjrJ
JriKIpMCKL5V/NyqUTwQ9Ls9+GScPoxlM5yBs3CVNVHXjxSBw0Fca+HvoLSLPxeX
YrpVKNNULEEPacwtFrsUX7lGZf0uhCeYQzzh1DAeEq86c9TpKdylbb4n7cAj7B2z
tpYrkWimWzGk6hyZs4ElLnIVYZ/vcyNt4mULoCbZfBkeW2ZgUL5qu7XYClULT+zL
aTvnZFypHKtySG4oGFDiUiCz8hQUhADGoc7jcwxkiEp+IqcKj3M0SazdWzldLtXY
z2Myaxdc0pFJSuGkXt7VO29k57Tw72q6vaFGGgnp8cAca0DFeO6BuDeI63de2q7k
K1DPAxNKfulBEHyqzuuGUVc+vwymoLYUzdBU3sEhXdnQK2IQQtPvC1VMnjUz84MV
BphUbBv5nATTJV88ktVSTXMFf7VIvmLyDMJrfWX0Rl2mrnSDxB4U7W275nn+p5FY
GMjystjFd0FcGq+Xnp+p0U1D4qF9LYM1I6SWJ+1A+Fd/lucH2vcET11x4LxNxAo3
nb7qowsQV5Q2wuxQPf9P9s14ZKh+OE+OMu/ekQKx3o/QI6jsyD/8oqXjZ+fjji0y
IaIrUYAE0YyDw2DV1ytZKrrlZAT0zbaeLUnJirtiM1i9LBpnpN9/K1czH+6IAM3F
LPbw0NY0phR7EDlcnKRoGmjy89qx/VxmXQR6dAYICpjyXr7wMg5ujYDzZnf6MVzb
hrKeFY7PvRq3A1lofd7mPutlgsGhNKeYHy+UJN2msRAe6PlMaOKQPSmS+AD4v24h
QqSFpu+FqcHPyqIOGDmItNIqnG2Ch5RnmM8b3rqqZGMgmFlI2pwY6hPjMQZZLaOw
vQVZ/foz/PgwEdYAB5sNjYS8CmOd6NGrRGSpSUvMEX7/wVG+0CMu4QijR45VMGTE
U11B9Ojoi5P1nE5b5PbIvNyp1nJZn3KkOUbU2wZy3jXlBxHyCM/Ccnt1DtXARSGx
HcPU4j+0JRPW3VOXJZVt7rRttqXRjU9KWjUaSE+gVKamBC8ASvNeiiI52TqVFv/9
OYnYO4d99N9rA9lXv+MloK7z6zRTrBqIKfMhavenSKx22nyEYb0ZfaJZigG3CHyg
oKYkJtLgvaGEF4aXDZeHpEJpJ8q3jQ2IL3JPq1C96BHozcEc8UnEgAxo0mEhvzcG
XfCCmw/rrmVI0wmCCgMAYXJ7zhqHhCbG/H0z+w/20GHhgkXKOhN5c3VG0l8q1AtH
EAWt6798Asdr84hlzP/cJxiFXjJGwf+mEyx6oQrkc3aR2tKAVeClQ/wm/xCP6qxf
mgkV1R9OBlVg/H3al9mvH726JjMh3wr7bBIk5kArkqk7/sYZD4/FUoaSqgZf/HMi
I/tCdu9m1XyStxVO9l0T/IIXQK+dRP9lKlaCuMjjHptlM7Itx6sJbavdqZ4B8AzZ
CrxCR7cXVIqZplBbsSQlWgXC9N2P40Mq+JUrfvZdj7zXvCBv5W+xvPxpDTlPblwX
tDTJWB5ss5CBxR7EyU58Qxnk8nZWxJm5J1/OPONVmLoFshpj/KBD87QzvRQh8UbQ
bqdJ1xquV+epkQJUxjJ0DuB3rjdb/0yV/1C1mMID2wYnUowoKj+9B8oAER6pVtjT
e1zq9q2SrsRWFqbSG5LvOpeYvz/mLk5INqdZpmpzbE3oMlR/0GBDPOVEz2RHOi3c
geByb2wkY0A2zL5wHcaXR7FWNBdHkoOZO9wFDEgyFpq1Oed8UE8Tyce+eEZL/C7K
J7h6IXe7yx6JSCxMRxP2ARyqUEZdb4H2ohjNF43XTiO/4tD9j3p0SgF1Rktz3DQF
viwZm2FdvoM/P7u0ppPqoIjkBNO8sCwtQU0D7ipnRlgHihZKTJyxIchPBh1paizo
QXuA6ABSFxTHKteKUnqKL2EoQEbf09JspC93kZ/SHzi7SDv4EUFLeBf/wjbNxKih
QyxUtEs+IvDD8n8dYspNnqkGJqIC/DoFbjvQj8ZoABway1oRrDbwnVEQqOveVi2T
HbqZ2ke/ghcozk03Ix3L1AIxewcIlKtpstesQOPRtahkaetIJ93FkQPy2iVqgBxD
M2zpEbZpxNQHkbW0JQry/BxFfs0va7Yv+IRBroTIPvN75IF+sT8nSouo/KxA2ND+
ltu9pw30ZVU4C6iJze6wNCV4jyVCkJAUSyOiNzE2SqwYjX15odlyujO6bM05v5/c
Pr8seuZ2HGZP5aj1MoEazGQ75wuIn0HA1Jx5W1rfOrIJ5PvH9UtWghcM59p3cv7g
0xfqKj8apW5Fzb5ezaVvvgsJ4UZRAHRja3beVtx9dTxxa270ktjPKdaiqCDuqVrH
d3NbEuK4g3dn7MkZgQeXMX11BBUegBsr3mntwz4qXsDpIRKRBp2l7H+ZZk29AU4u
YIzXATorf6c6tw/Hr0APMfVjCHv+wl24Vij3+XVguxRuuOiJkhPJm7l7xuxmJlsB
PLUwzxyxSg+t/L5h77oas5rizN3apUmZZCU8Qn2jLMlb44b9Cew7lLMVg0nk8RAU
6DyR1jxhICMqYi/OUGvNqyherKQ82x72vR3DKYGCceY2rouaqpOcG/901Bhj9lcW
cjvyZPdUxbr6h+y9X2jeAPXKI9irztK+5Nsau3Tg8xbSsXUPXJLe4Ola7Wuw1NlY
XYAfTSElf7TvVFO3iZpKfHJhMDgjxMRCUvkyHmtLITuUZk3Ku+/BtnyQpZ6siEBC
UkqIUaXqK0CrY5qyZ/89jHJyvVC1knJ7xC/Curp6U9Djb7ZK4Ti3LrFPrSMPK1AQ
R9H3YSkuHi9N4Szf6sjLYKc/x0nz9KTmTWLdRS6aAFWTVMjhEU6LfYRDAnWenlC8
Kmpg/Q+gW+W+nlZLWBeaMm5kjGTto4fm++4y6/B4CiugOD0pfl1q4S1ftf43a9Ot
P7iVY/Sb+2s1xdbkS0NUW0pKY26+wnUq9ja3bRLeJ4sx1BJxmas46LHIDfStV1yI
ixAoTUBML7+z90yYMbfPh/XQV8kDdnVbcXzvnGqr7Xa2qjy+wjpsOYboNQrPzieC
7Cm1vvJGgb/8Zb1bmANHzgaB6EHvf0SwE4FaxhQI+eMmcXboa6CvF8/39SSEjVGB
ynwygJZ+++5aLGCvL5ca5eAMzRWigCd76QCzRZeN2+6+yY6X6yvRg0m8CxVpqIJV
zWwN3OZ61GheD3vvOg9RkYW71IzxqMv9bXcuQy1azhnXiaFXSOwAOejm4OmwnCjA
EetNpW19nu6/qkrGwwLDJkSqvUKlftqsINnk4pDMC7+sdG/nzfTMz3AxBZkzyDd2
MUNJ39euhc5TroAvJsTml2SuU/SZFen0z4S78iZaDR8A99qtkKpjDYFVianZhlAE
/06lsgPv04GzNdHhgZqEwgpv5OOQ6/FVpkUw9ltpPH/RpT1eCukeIHRttplSUeHk
//bY5cfNC+OMl71XJotbrJwxewsMzlXs5chd9+tTv88ZR3vciPD97rw6n4pvzXVl
a7P4EvG6y+uOhfJRfHKVpwDxwdfjEqWy4uHQbUxJKoKuSgjTfiRx3yIod+gqrCkb
FRIzX4yEwsfFZ4tdS+ck55Z4ONCUa7NfprLcgc8vZBcAlCRVHXRpyX4doyDPQE5F
IyBFQFYZsPijEcKv0Wd0uw3fBbWVWjrF47Jxj8QqutB8ZHw0/2ioz+xHaMqe/fwC
WxY7xXWWwKFnITVAvEA57GMjvVCu+1fzSUhzcTQD9N4V5xr6tmowaOWlwiCqQq3J
k8XW9mLjfKkY/39i0RYCvs05b5j6isKR8fc8z8r+zaeELpcEq8Wim5mfS9hUIWFw
kFhRCrJ34kpISbAXjy1Z/k4gjvec7QOgoU08PAsTpxmLN/wruBBQehHgBBN1JTwW
8yjRvouPAnr0OPQ70lEQsHpY4j8+ePJ+5LdWKvPsKcHn919wi0SKje0NXeQGi2jZ
QC2CW8tmXivACfX1uDAwTe4SWyPtVFfOZsqVQfY8OIIrW4CI2rNcjvt0ocOrbxit
5y8bF2C02xzwCUo01JDfoP9nerPGn8brSvMEzGDERW6Iw/8Y5IaPa8sOcvuPmalO
6XuTBYx7aN7J45IP4PFXV+vT132sgE13Jfe3bTRwckSr/cqgRvUJmJGDnDvxkNCD
7DMAFMuJpMAXjkun9EDBSfSWGXq7ji8wUFqcPRc94pPkM6ZbeDlAX+ljTB3XjdRj
48BEEOBRx+ljwDEvUx7xcUDKpo3vObGTD22P9zyMZC0NqjYxkwaqR6cN3X5RXXXN
gSejaBuGZr3OLhQthliCgsccmG5+U9YOuAHdfaHuvWOxuIxD5D9vMGhz7v6cZ/rC
BL4Jd01a6J8PNxWXhTng0LSLHr0GRddW3pGpG5nVUz8CpiyApITde6thLQsMwbr4
sVco1j/r9T95lSx4Zq3fKvADklg+trQafYBfMwBkX/Pr9W1XBi7lBEXj3mKcrrTq
Z5GPnSuxPbVvBACpWEKf+QcjbzdoIA9nVvhU9ZqtsnQWlNjO7tvdUS7esCxMZeqF
rX1KcFUMt6om8oyKbiQeSgQzenIEnF8vTo7GmzVNrbxbdOMPW2n9peevl9aVX1CP
m8dCRK39MhrgT1bPYLg5E408BUEUrfwrOvJUg+BILQj04MSnUGfs2DH31o3j3VaV
1BDBQOEonMXEF6o72yWiV2+7rmbfJzdkzdANDBh1w8SfrV1Ofp5a9/ycm9QPC5FY
o8e38RObBusVI39w8C/fzLZNixXmchi7G1D8xP2SjJKfhjEoYopfI4afpNFgSpMI
d4iNN2pukGQyC9W6224+wTRvmWPXXkE3O9U1i6fxOgaIIKdF4UB8W4hRbN3z2qfD
qQ2GZ6bRjGXaxVMQ9K3fMgY3cM8ARoMeeo7xjK8enpJ6rQeXIJVu76jBn35+N1Qc
xKLECLt0fOvB9cZXiXgWHV6jwz6mSSw24QsRnmamvLejv3s1MDrKm1lERV0NUaCf
QiMAW9A5NOaZ9/7XaqIizrdb54HVYIIx8mhiUBOB2rw4YhZNjqK8WVONQwc6QT9b
mENe/c3iJNdqbNTAqDX7qJY5hWiGUG72sWincOFhOMktsiyqS0I5cn1CshoAJ8jR
BzTyW6/v6+rQ2Fh6QuNLYEg2twljcCvRtvcE2qFa7oidOCzO0VtXviyPnDEiu2kc
KwYKwmx7lrJSIilS8dAG3mn9630cTvQV0/Q9yUogcVW/lXpbsh4H+NVnhPmM46/Q
m9iAf72kmxBbgCQ2eW3wRYggmfgHnux4zrGLdTPB0yz/DRL7HAv4vl9JvLQHcpX+
P5esYY7aFgzEVodXUs51aHrYe25Q0+TKEK/rop2uyYeKa7hR18gij+jndLUq5Njg
BTmpVd2lXX4afcp4WxMzdRexFc6RoPse4Ul2+9t4AYdEnJOIDBUDUBjmJ5DtpZtU
WUR6oM4WgnhsmJ/Y882zaUoXdrfT2M3NTTEklmr/79V0hwQ+Fvy8RujztglIL5m+
K7HFRWC6OSAX0eK9ujJdNYFSd65ALfIPnrxO7OGCGiJzu+Oi2GHN0l67dp5qX9P/
tzGnbZkEtfOaNJN9PHJw1OPGUcfzJL9ztcv0pSBtIGU8X7iENfKitjDOd8l8/bVj
etf7kLT0MXLx4Xau7sxnyO1dxbNCXOSryOIV/m2HDDSGiRxeJwa+srYt/aIFSnAC
gifinyicm4IialSN1bLDsuxWb0KFwEi3lWvnrfoFHUk0UW6HaFCtvOYx17Axrazm
7nwJN4sgHt9dUB6+kxjQ5ZS+EkF2q9fhC3V+lV4PWvd27yG7pQy/yWryOpZLmnYQ
pWxM1znktfrUcn69tC4Z3PxktRJOVPAfKTZ0jGMQ6XNpy1mwaYrR5vCP0nGpMRHK
9F9Be7O6Duq8g+McPO2D64HOSxjK8hswhx7ia8OxPLK6JemYh1SWHOKsLOeoV6Vj
Bpu3JkTLqqHpPr7+V+f0yWD3Yt+JxRIZS7dpN4XMxkGBBCchN1AJcBu8MX+XzGD5
zYMYYZgF4l4hk/LwKeFmkDDLhEG1ltrpnFHvrRQk0DWuiDAGRbteGAMSWzYoBwA2
+mQ/LB0PaXORJFhZkr0FrQxLVjrzgn+zXDNjP57QOL18E96ptFaEOS9lUSfoAnG3
V9/K0HbBaE43yRNkNDFxrbJ/j/bQ0bqvlObxYkXGVRrthyGHyk48LWehrzkemj3e
cFF0UvaBDPAy3GsTFEzSUL1opCcNfk3q25r9FP3U0OMWWPVZVmOzGAz9/Rpl9qzo
WQPHoCvsFg80cDMpNNUtBJ0UTV3/gv9yRkNqVPPOO3sTaVULGaMI7bTXImSLMY69
v43/PZjSpPi0RjPqfwPqqboonfXyhclK3ws+3yxGhPiU/xDlo3iX5LgZosmiifZ4
`pragma protect end_protected
