// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:09 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BjIn5RAf+ibdsIvHchvgqyMQNLWvKTTMogfmhzrtTd/VlZCbphfX4vqyOQe9JSiK
ACKUF7MzJlXExyL875lvq3BOWcTEjjQitdZ54oA0Lss9+h1GE3P62vzRXTZBPvC0
t34GCQhtol9xyrxE94BHMhFwE28S+0dkuRVYF49m9Xo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4848)
c7RilAQmj2JFccq+DfG6R38gksdVrlrOH1GRw8aRhSeNgjOTKEI3PP3VChtLnS/T
f9ptvo9SCOwVeLlJYxGnVAQZ+bN/U7LQ/hx59fxCaESIAeSijUsNc+tEvCjlidvq
PK6zpQ2GNkAT2xwO3UmSSWbWpiXyyuQtoWTz/hq3k9j+aClXR0fDRSYPPwDK4jI3
yJl8GgZCqwtnDtq5bPSjzS4Fyh4pprEgk1tf3khxrMb3JgGuQr5g5qayt3c3xSO4
vCYXda3Z3Sx7o12LliqSZYJXInQqVG2HQXcFERrhBfEtXTBwu1C+Qkifnr8ooQ4R
lK49vLMSfIaXx3P6p6K54uGPDoSiuOx/FKlb0ZiLFpJyX+R0DPokHywTaY8KuiV4
sVe3XHInk+YFP8wZw39AOt7lAHDKMu9dJ+glQZe5Rq8zzsnYTrSgrV0WGbzNx1JX
mld4+TQi9kPKdU8CJm3X7rNYwmIMtbiKso7f+NN1YvbNbm0KVstF1p4bL/YcblqV
CbmNFh9yR4nSjfwBFoHu9oTMpHDUcjsFRv41CwiG+VhmlSvHC7QZ06AxiBn9h35A
ool2ZWDtBg/RY7Hpg0mhjeFWAX/yLys6b1F6FNs2bKYGO6xYKQKN2JlutT3L4TM0
GWjDSpVeWGp5X5a4hQf3dgzQGNbT9Hc7mynb8v6zPSYiICuFuKq3HHCczNEp/Rdl
A2atyF14x07S75WctAC6E079wrtEF/4VgNo6pcrnTE7iE0uN4Mz5vZCBmjcXwYmP
FNIpqB5XMr14SRQJ6hF/NvS47FBDLPaBovw3m9Mdhc03QJQbV/CzUrfqmAETYNT3
xQs+wYVmffiT6HYK1quymJgVoDdSRlHKG891raPxlq/lghMdINpqyKRDv7Fz1RDa
ena/zzU8b1Rj4LGaz1QjP30VBffJB55PWstfVSQ7iUG/yyV04QHI5RMYhBDl5VDr
QeNAXp1h6t2UuiHDarRn3Z/2cpzgB8bOKyk8eoHGgJ1W+lGHkXxJ0fULntWVMLf3
2s/YIU5+oP6O5UHgpiwB9oHyKz1DecZeQrLnXtHUzd/jLUHSPJB0cVfyThQ47tSi
Q2sNKdDGg1EpzwvNOLJO7RJ6AUO4iHLHfG85gQfDzF159twesWfcBGVuFnDYHn/6
obOXrBcfVAtsNTf2wf05CRwVNPS4oySPQhU9kWV395DiUpgOfRFzRG/O6dP266cv
z3gdcX1N54cO+iS6cVkGDIF21CdyNJ1KpNG4CRNIugo0qUuzsj+NcwUpXZmAc7YQ
TZIc1RKkOfMf19dODJvzqbLdm5/nm5IBdclE6IUO3CYyPIk6bVtig8FBn7dws93Y
IhgZTyAjXptGD52TxgjKZXZ19I6DOVlQL4gj42jnlXS4elhY9p56omTnLfcDqLf+
YjG2zy5qwRFpwe8CUVNqRgst2BgDgYaZ6fnqZ4JyqI5eBDySNLK7x/hLG3fe0MkL
iUH9y9qMOj3EX85pSWH22KSXOebK+3nd9pqQJv57jdR4HK1gtus9VjuVwGITVu8H
qnQ+t53SPqdloD9qjRoNcb9w/xTO2J45jTD9XEbrmFykQwCJpMgCcyVF4fveMRdn
OHdQTs2pyRKTa/71AHy5pPLXNhBV1LfbFYmxLlQpy8xpL5y7r+henJ0qpY8/l8kC
TS0iANG7iXj4mLdvjrR3Xcw2A072OIrmJGU6OZwwdJIrdnHFR3erxK9Il0bagHwM
/aK1DxXhgeF3Pxg0Z6lMeyEDR0s23ghB3Lg6RTT5VwPP/0Kx+DG+VZs9BL2I9Gwu
eFoKJSMHoj+HltKGuiSPsWmjD0cWzEJ0ytxTRJ46C74oTgRjGInFlkzZdrJAaYco
ZUg4ojE9EHoMw9TTdly5Fnc15bzMeEcK2o0J7JCKtis7ZPYCDJ+vG6CU07EErmGh
ULdkvp0znsoGNGosIyXmq7QQ9h/2hUj61PiCyp7HlM4ZSTzdyLD+eTC7H1U1USI/
BmJn4KHzVOUAuIDKEZLGZ2iCCXVZSQvV1eWk3jSPATPFDh4pF4ymuW+EetxJXIZN
aRURPDCmcPYvM6ykikBtkynGtIKGHucB6lITFeqXUXnelg9YS/mB2j0OEa8TST47
1zUA2hCKQE+bxS15Fp5P2t5MG+Ab0tTB+0v1Q8DGpsx9K8xTVdy80Q34edyigOCl
IeBOEa24KAwNbD5bs8jQnnFJh0opN1330iehH65yxzv6MuqILv6SViw1C97LlsQ8
HbZl4iL+jQHLDKEfvsAu9V4X0zZXh6l+xz5A5DGsdtpwCDLEdlTn2ktE7vg0NHRR
l4TLjjgtcsU9cA/mnA+Rw9AG2CRmIa2xP3cCkTqfNWsUDRgrsu5n8KCN+9tdVCLM
swDnkMOAK4BMigBHR4Gdsskx8LhOhtIqRiqFqtXrehtQXvgZwwsIMzkst+M9zUeK
JzM0iz3b0yQwJD2xm2AWDk2rtcXCxvajR95pNa4H5PrVL1vursQVX6PPZ7Ljda6f
RHi4Dqel7F4VWRtsO0Ia7mMZDIsrJb3gadbohdRpIyfrYRlsR6LovTiYycNM4jGU
fqirs8khdX8qTSGYQN3uuSLu+AzPkceVcOx0rwe1Z6DlgeIJL9e6lgOaR/ww+JRF
UtoqX3D0Y1DZ/IdBYjtWKDUt3otHUUmFfYBmvs7vCSxQR/X9v99O7BMmy1EIXSZF
g8jJMmIknvZlbSsGt9GzsF6Y54LDNKC9eBlIfwk4zfYZ9bbabAiGQiEIoeSz4jgW
5ZkTx/AT7rTkVt7MCqhFdIrDjLE2mxTRBYNiRJcuhHjrx4L0yB1lZMlr9iBlkM40
zRG12MoaQRt7M+Lr98uXIs1P82VpfaTjdgy18ZK+lQhS/Xaa1TNuUnzQC/EagvsY
8YcAVMpeRY/5c0RVS2FptvObMFT38HXlpKtDPz2TUUMsb6qTakx7kDgnFaPvgrf1
ZYpo1ti1mYwKWxnVJyQ+ciN8zaGniv6uMZSjYrCVISmVB1OQPVLNiV344yZDizms
Gd/MhEzb5z4cYvgmoGiS9a0yayls6jFABRi+YzxrRS1eLzV6ddgnrv09+Ra/rUY1
hFk4xc9W9XdDMEb+TQhvGggV27W8BHDh3L9gGILF9C27ncoBZDZctuCmx303h6Xn
o4+PpK8nFrXAhFWjItsdi8wvuMWiULfthpzbb6x6oUdM89E+W05BIsbYtfYWD74i
NYQFhiqaLp8GwXLPliXk0KLd/BM+5DZCSyHQkNymVmQeMBQRYYIqHP7S/Msu4J0V
tQ69UjPIBDavWklBqK0pJQ0RuEg3QRTwKBrko/U5B6/0hxru6QWW/TcKlZFBge25
QL+S6ie9VTo/bW4NstuK1H+XzIOV7aZPNRWhvCPbxPuS8oTCimYsFnBVwkfXrRoZ
t2/BeCQJAC7ikQk8SbGmqAELNgZU2AQzYrc4HSWjF+BJ+Bam3sj3CweTecZ6a+nY
G8R3VCkMS8Fp4fIuoAJPPJaOGQjACkD9BLRgbwwm2qQ6al1Ya8eu9mmjzBmpkHMl
rJKl+qcqKbEQw5I4SNm2vsTpfBBbquUr8DSAwkGJS9oIBcS+YVvbC1RFi0EYt+pl
WMbkxdCmxFh0bjXRjsp4eJrCrtcsmfzkpGXIFr4aubzVaLrgRvxIJS3DM9iBul3L
8WRDHS+yjjd60xjreqULmC2azxHGWsHnvoJ48OCgtNT81dadi1BHb9CcPR9vUQw2
+MY/b2AaI+etQvHmwcL3/BIZnWITZAn9PWjIgUdriEvwkuxhmWHOfz50ZdKZQ1sI
epZhePYgSs4/ZFL2MPlBkEYramBn7yqHgjURrL7C07lUFU/1UYHxI/n1hw+0sC3v
rWvUuRSetK/rOlIyhfGwqCnlNcvLFpT+5zGpGNi3eFTlFtYxcJcNxxGXzXtAOKUO
rkUyeLDjzwt2wQTSarw6YuISFCE36v8kOCrybZnP0zlLsn4sPgXrRDRe7k7WEbe9
o7xGJJznXBgk9YoHr/ZKtiHv9fcMGd6l1Wh9Ncwn2gdLOrret5WwxDxiEwEdZjoU
Pc2X8t9iht6kdGRme3ZJHGe4zPRL46fbrypcblccZBLeSVCQ5THT/b9bEKdxmSu4
JbUgC5y7vVJrDCYqP+VUkCIpCLwQXgxFK7nR7UPB5ZPJ2rmNo46HjoahBZvhUoaO
DqYkmU5AIbPC7bGUrW46NzLI0zItV+jKVZ70za+5vfZZ2cFU+oUcPO6fvbr+5e8f
+/5riaU2HWSkW5R7d25Oq7k2vTfaLzpn+vn455RHDATfk3Faaw7lSQPBmdWozKsB
M7DICn1+o3OeFk8HwYgCjrfNwmMygs8kauyhX608PtB4Rn6WpKsHYrOhMq8ONI1C
JySQKvbTM64oftcbJFM5Y7Ie13gs2sYOqNbBhZANoyBH8GO1sE+WADURx8jWU1/U
thuITShnqmZCQ/TJqWwS04KNaHTQbeYq0HrsBsHPGhaLsWFJstKbK10/JKqmHSEJ
Q8h9yGjckHR6shV4dNcfniSrFC9HEziNcs5FSlBUhjjkxhMesknvgZJNC+Ff3G3s
WJcAiURjxsmK2BZIHZOOCVdTlYUBi+lPOgsx5RgsomgzIOVH3RY2AEXujRMvuWCq
/BvzLcbzE61Qth8dPXZ8OZCF7DR2x5KiUi6bLB6twCMYOSGtwlWgbv/5JcNRX7g0
HowB/rW9jPD7nABWHYpD6TUER4i7muPPQ/teTHGBY+7WvNfxQ/hwyCJ2a4fne5iE
j1DqoHqSF5zaLZOFKXlnqCJLsmJl4x6egSZ867wvqIDEzWrDFbx/rCDzmtMlE5o8
ntpgIBk0Q1e9gmq4jdMlPDf7qaRRqnOPWbsNX+BjtE7W4us+CauEEzTSTTIAmpNx
1J++N8u8JUiCwUxK7jj6i3S66G3LGpxUfeP2Oz1AAPXTn0vdgupoWI6hltmb0/I4
9NhwXPZOOiS1kYkhrqsuFJz3kNj6U9B60+WR313iovh+xNSqAhWkIq5kuY+QjSyH
kEleSOKhTEmaLZen34yeu3dFfhvjrBdHCakhPNrNAOPEmCH3Xnq1xXvBJkK8hVqc
f1eSz1I7SxM36bYTzkTo3uL3fe9BnzyzUhm3snIve8dxmy5ELfGI+TGmdv/hEfDp
WMmooBj8I3UsSm2ui/9mVabV3I7Y0sSc9Dpb0S51XQlC5wTR73asDIxajQt4xeMl
tA+i7SupmziOFw5HK7KGjTfQ6vTFHYk+mgGVkIIDY/mVmdXX6HbKvJymWVvIHwRt
/FXshqRhrkPRGgYUwXuVGvX1ksZpscxT1TPAKgUR4ka4SQwlRXfFVZGv2kjeigCC
SyROIvHNhHCS8yl6R6uvp31D8EG5FfyH+zd+GrPuEfd225k6jjnk87Nw1TEC3yxi
iejWX0JqJibyUjLKWamda4CjFTA0X3LGf5uaytaX9uS/jFssBafUwh6nLxnUTTnh
tSGQ/QTxABKSBh1lvdItgKGv6aFXPWllPTgcb9mja7RyJNaqeui8stlPxFdjhc+z
bdPZ4ytGWqkKAvNO2DGB48JT4VMeZgjnUAcO7WPbs7SH9W29PxeTOeqo9qvlbIyl
rhJ/vaYizTIIQZ1roJq4fnDRVhgBOXom5pFvQS8b0RZGTFyD179nPs2R7fBMPE15
3IGi3YTQWR6GCBqOL70s3IhuTAS3JXiRlVNiO44Z3z6lvG6O1UVcpee+5NpUZDCt
5A8PF7HqVkOD09C19L7Eoox3jGtelXZLf2H0YfhYMKR1VoMR4DiSPmP1pcDoAuZ/
VLHrMS38AIOLKHyXOe7lqYNePb5BUlzJJ/nkqBs+Rh/x3ym7JpLhUmUs+RlFreRA
RkcDCBQN/zVgf+yUuBfZW6A8btgupLxhKCQ0NErKegrBUzgF5RxVKj4RFRCNjyvu
uRET2OFssLk9YErbSmEZlDhZt8rt5r8Zx450wDpW/0kqJ4kiATXgEt711e7stOjU
k8A0pIWxcCMz9Vd7xfs4Dvzm7xWfowXgvJU4x/h3Numpq4fzqi2z3nsu7y35JY7C
zP9nIhjNCe0WQd2TQVec5N+2WcJsuLJTrIgjDOvCfh0VpEDPo+3bRNrP9HpEMhNg
Nn5gqWlmiJY2RNqAgGa7h/YGGQJiNCzssQFMlg9Lh9kpV9BpgSqmL2zMBs20+V3x
vHsOvKcunhR2tMQcpl9z2EcfdoMgjcNOdUZqbg/B8YafXEVlozAkid0lvAzoApev
8diFInN8EX5nc0+HZMaz5XZcwqnFlOSQnPnehDDkJQzVrZkoJ3BlOu+Jnc6G7Lg2
GNmLC/RQ/kwg5r+CZ3F4105xCVIMKUk0bJK5liTEzsI23gjU/I7/PGtPNZDm04bC
0n7JMVEgl8egYqVQid39PZo/2owau4PJyMxv1wHYfzw48wyVYZlW3a8ESPXmBmqJ
V1DrZgWQJHAL4OzwxP2PmaRuk5/QSRZCUOq6LK5sWLzYM2x/na7ymT8/8JXMH53q
`pragma protect end_protected
