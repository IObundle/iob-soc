../../../../iob_regfileif_swreg.vh