//data and address widths
`define UART0_RDATA_W 32
`define UART0_WDATA_W 16
`define UART0_ADDR_W 3
