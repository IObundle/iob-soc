//data and address widths
`define UART1_RDATA_W 32
`define UART1_WDATA_W 16
`define UART1_ADDR_W 3
