// megafunction wizard: %QDR II and QDR II+ SRAM Controller with UniPHY v16.1%
// GENERATION: XML
// QDRII_SLAVE.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module QDRII_SLAVE (
		input  wire        global_reset_n,             //    global_reset.reset_n
		input  wire        soft_reset_n,               //      soft_reset.reset_n
		input  wire        afi_clk,                    //      afi_clk_in.clk
		input  wire        afi_half_clk,               // afi_half_clk_in.clk
		input  wire        afi_reset_n,                //    afi_reset_in.reset_n
		output wire [17:0] mem_d,                      //          memory.mem_d
		output wire [0:0]  mem_wps_n,                  //                .mem_wps_n
		output wire [1:0]  mem_bws_n,                  //                .mem_bws_n
		output wire [19:0] mem_a,                      //                .mem_a
		input  wire [17:0] mem_q,                      //                .mem_q
		output wire [0:0]  mem_rps_n,                  //                .mem_rps_n
		output wire [0:0]  mem_k,                      //                .mem_k
		output wire [0:0]  mem_k_n,                    //                .mem_k_n
		input  wire [0:0]  mem_cq,                     //                .mem_cq
		input  wire [0:0]  mem_cq_n,                   //                .mem_cq_n
		output wire [0:0]  mem_doff_n,                 //                .mem_doff_n
		input  wire        avl_w_write_req,            //           avl_w.write
		output wire        avl_w_ready,                //                .waitrequest_n
		input  wire [19:0] avl_w_addr,                 //                .address
		input  wire        avl_w_size,                 //                .burstcount
		input  wire [71:0] avl_w_wdata,                //                .writedata
		input  wire        avl_r_read_req,             //           avl_r.read
		output wire        avl_r_ready,                //                .waitrequest_n
		input  wire [19:0] avl_r_addr,                 //                .address
		input  wire        avl_r_size,                 //                .burstcount
		output wire        avl_r_rdata_valid,          //                .readdatavalid
		output wire [71:0] avl_r_rdata,                //                .readdata
		output wire        local_init_done,            //          status.local_init_done
		output wire        local_cal_success,          //                .local_cal_success
		output wire        local_cal_fail,             //                .local_cal_fail
		input  wire [15:0] seriesterminationcontrol,   //     oct_sharing.seriesterminationcontrol
		input  wire [15:0] parallelterminationcontrol, //                .parallelterminationcontrol
		input  wire        pll_mem_clk,                //     pll_sharing.pll_mem_clk
		input  wire        pll_write_clk,              //                .pll_write_clk
		input  wire        pll_locked,                 //                .pll_locked
		input  wire        pll_write_clk_pre_phy_clk,  //                .pll_write_clk_pre_phy_clk
		input  wire        pll_addr_cmd_clk,           //                .pll_addr_cmd_clk
		input  wire        pll_avl_clk,                //                .pll_avl_clk
		input  wire        pll_config_clk,             //                .pll_config_clk
		input  wire        pll_p2c_read_clk,           //                .pll_p2c_read_clk
		input  wire        pll_c2p_write_clk,          //                .pll_c2p_write_clk
		output wire        dll_pll_locked,             //     dll_sharing.dll_pll_locked
		input  wire [6:0]  dll_delayctrl               //                .dll_delayctrl
	);

	QDRII_SLAVE_0002 qdrii_slave_inst (
		.global_reset_n             (global_reset_n),             //    global_reset.reset_n
		.soft_reset_n               (soft_reset_n),               //      soft_reset.reset_n
		.afi_clk                    (afi_clk),                    //      afi_clk_in.clk
		.afi_half_clk               (afi_half_clk),               // afi_half_clk_in.clk
		.afi_reset_n                (afi_reset_n),                //    afi_reset_in.reset_n
		.mem_d                      (mem_d),                      //          memory.mem_d
		.mem_wps_n                  (mem_wps_n),                  //                .mem_wps_n
		.mem_bws_n                  (mem_bws_n),                  //                .mem_bws_n
		.mem_a                      (mem_a),                      //                .mem_a
		.mem_q                      (mem_q),                      //                .mem_q
		.mem_rps_n                  (mem_rps_n),                  //                .mem_rps_n
		.mem_k                      (mem_k),                      //                .mem_k
		.mem_k_n                    (mem_k_n),                    //                .mem_k_n
		.mem_cq                     (mem_cq),                     //                .mem_cq
		.mem_cq_n                   (mem_cq_n),                   //                .mem_cq_n
		.mem_doff_n                 (mem_doff_n),                 //                .mem_doff_n
		.avl_w_write_req            (avl_w_write_req),            //           avl_w.write
		.avl_w_ready                (avl_w_ready),                //                .waitrequest_n
		.avl_w_addr                 (avl_w_addr),                 //                .address
		.avl_w_size                 (avl_w_size),                 //                .burstcount
		.avl_w_wdata                (avl_w_wdata),                //                .writedata
		.avl_r_read_req             (avl_r_read_req),             //           avl_r.read
		.avl_r_ready                (avl_r_ready),                //                .waitrequest_n
		.avl_r_addr                 (avl_r_addr),                 //                .address
		.avl_r_size                 (avl_r_size),                 //                .burstcount
		.avl_r_rdata_valid          (avl_r_rdata_valid),          //                .readdatavalid
		.avl_r_rdata                (avl_r_rdata),                //                .readdata
		.local_init_done            (local_init_done),            //          status.local_init_done
		.local_cal_success          (local_cal_success),          //                .local_cal_success
		.local_cal_fail             (local_cal_fail),             //                .local_cal_fail
		.seriesterminationcontrol   (seriesterminationcontrol),   //     oct_sharing.seriesterminationcontrol
		.parallelterminationcontrol (parallelterminationcontrol), //                .parallelterminationcontrol
		.pll_mem_clk                (pll_mem_clk),                //     pll_sharing.pll_mem_clk
		.pll_write_clk              (pll_write_clk),              //                .pll_write_clk
		.pll_locked                 (pll_locked),                 //                .pll_locked
		.pll_write_clk_pre_phy_clk  (pll_write_clk_pre_phy_clk),  //                .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (pll_addr_cmd_clk),           //                .pll_addr_cmd_clk
		.pll_avl_clk                (pll_avl_clk),                //                .pll_avl_clk
		.pll_config_clk             (pll_config_clk),             //                .pll_config_clk
		.pll_p2c_read_clk           (pll_p2c_read_clk),           //                .pll_p2c_read_clk
		.pll_c2p_write_clk          (pll_c2p_write_clk),          //                .pll_c2p_write_clk
		.dll_pll_locked             (dll_pll_locked),             //     dll_sharing.dll_pll_locked
		.dll_delayctrl              (dll_delayctrl)               //                .dll_delayctrl
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2017 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_mem_if_qdrii_emif" version="16.1" >
// Retrieval info: 	<generic name="MEM_ADDR_WIDTH" value="20" />
// Retrieval info: 	<generic name="MEM_DQ_WIDTH" value="18" />
// Retrieval info: 	<generic name="MEM_CS_WIDTH" value="1" />
// Retrieval info: 	<generic name="MEM_DM_WIDTH" value="2" />
// Retrieval info: 	<generic name="MEM_CONTROL_WIDTH" value="1" />
// Retrieval info: 	<generic name="MEM_READ_DQS_WIDTH" value="1" />
// Retrieval info: 	<generic name="MEM_WRITE_DQS_WIDTH" value="1" />
// Retrieval info: 	<generic name="MEM_BURST_LENGTH" value="4" />
// Retrieval info: 	<generic name="EMULATED_MODE" value="false" />
// Retrieval info: 	<generic name="EMULATED_WRITE_GROUPS" value="2" />
// Retrieval info: 	<generic name="DEVICE_WIDTH" value="1" />
// Retrieval info: 	<generic name="DEVICE_DEPTH" value="1" />
// Retrieval info: 	<generic name="MEM_USE_DENALI_MODEL" value="false" />
// Retrieval info: 	<generic name="QDRII_PLUS_MODE" value="false" />
// Retrieval info: 	<generic name="MEM_DENALI_SOMA_FILE" value="qdrii.soma" />
// Retrieval info: 	<generic name="MEM_IF_BOARD_BASE_DELAY" value="10" />
// Retrieval info: 	<generic name="MEM_SUPPRESS_CMD_TIMING_ERROR" value="0" />
// Retrieval info: 	<generic name="MEM_VERBOSE" value="true" />
// Retrieval info: 	<generic name="PINGPONGPHY_EN" value="false" />
// Retrieval info: 	<generic name="DUPLICATE_AC" value="false" />
// Retrieval info: 	<generic name="MEM_T_WL" value="1" />
// Retrieval info: 	<generic name="MEM_T_RL" value="2.5" />
// Retrieval info: 	<generic name="TIMING_TKH" value="400" />
// Retrieval info: 	<generic name="TIMING_TSA" value="230" />
// Retrieval info: 	<generic name="TIMING_THA" value="230" />
// Retrieval info: 	<generic name="TIMING_TSD" value="180" />
// Retrieval info: 	<generic name="TIMING_THD" value="180" />
// Retrieval info: 	<generic name="TIMING_TCQD" value="150" />
// Retrieval info: 	<generic name="TIMING_TCQDOH" value="-150" />
// Retrieval info: 	<generic name="TIMING_QDR_INTERNAL_JITTER" value="250" />
// Retrieval info: 	<generic name="TIMING_TCQHCQnH" value="655" />
// Retrieval info: 	<generic name="TIMING_TKHKnH" value="770" />
// Retrieval info: 	<generic name="SYS_INFO_DEVICE_FAMILY" value="Stratix V" />
// Retrieval info: 	<generic name="PARSE_FRIENDLY_DEVICE_FAMILY_PARAM_VALID" value="false" />
// Retrieval info: 	<generic name="PARSE_FRIENDLY_DEVICE_FAMILY_PARAM" value="" />
// Retrieval info: 	<generic name="DEVICE_FAMILY_PARAM" value="" />
// Retrieval info: 	<generic name="SPEED_GRADE" value="2" />
// Retrieval info: 	<generic name="IS_ES_DEVICE" value="false" />
// Retrieval info: 	<generic name="DISABLE_CHILD_MESSAGING" value="false" />
// Retrieval info: 	<generic name="HARD_EMIF" value="false" />
// Retrieval info: 	<generic name="HHP_HPS" value="false" />
// Retrieval info: 	<generic name="HHP_HPS_VERIFICATION" value="false" />
// Retrieval info: 	<generic name="HHP_HPS_SIMULATION" value="false" />
// Retrieval info: 	<generic name="HPS_PROTOCOL" value="DEFAULT" />
// Retrieval info: 	<generic name="CUT_NEW_FAMILY_TIMING" value="true" />
// Retrieval info: 	<generic name="POWER_OF_TWO_BUS" value="false" />
// Retrieval info: 	<generic name="SOPC_COMPAT_RESET" value="false" />
// Retrieval info: 	<generic name="AVL_MAX_SIZE" value="1" />
// Retrieval info: 	<generic name="BYTE_ENABLE" value="false" />
// Retrieval info: 	<generic name="CTL_LATENCY" value="1" />
// Retrieval info: 	<generic name="ENABLE_CTRL_AVALON_INTERFACE" value="true" />
// Retrieval info: 	<generic name="ENABLE_EMIT_BFM_MASTER" value="false" />
// Retrieval info: 	<generic name="FORCE_SEQUENCER_TCL_DEBUG_MODE" value="false" />
// Retrieval info: 	<generic name="ENABLE_SEQUENCER_MARGINING_ON_BY_DEFAULT" value="false" />
// Retrieval info: 	<generic name="REF_CLK_FREQ" value="50.0" />
// Retrieval info: 	<generic name="REF_CLK_FREQ_PARAM_VALID" value="false" />
// Retrieval info: 	<generic name="REF_CLK_FREQ_MIN_PARAM" value="0.0" />
// Retrieval info: 	<generic name="REF_CLK_FREQ_MAX_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_DR_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_DR_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_DR_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_DR_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_DR_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_DR_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_MEM_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_MEM_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_MEM_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_MEM_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_MEM_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_MEM_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_AFI_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_AFI_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_AFI_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_WRITE_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_WRITE_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_WRITE_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_WRITE_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_WRITE_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_WRITE_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_ADDR_CMD_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_ADDR_CMD_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_ADDR_CMD_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_ADDR_CMD_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_ADDR_CMD_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_ADDR_CMD_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_HALF_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_AFI_HALF_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_AFI_HALF_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_HALF_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_AFI_HALF_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_HALF_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_NIOS_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_NIOS_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_NIOS_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_NIOS_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_NIOS_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_NIOS_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_CONFIG_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_CONFIG_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_CONFIG_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_CONFIG_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_CONFIG_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_CONFIG_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_P2C_READ_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_P2C_READ_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_P2C_READ_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_P2C_READ_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_P2C_READ_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_P2C_READ_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_C2P_WRITE_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_C2P_WRITE_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_C2P_WRITE_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_C2P_WRITE_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_C2P_WRITE_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_C2P_WRITE_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_HR_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_HR_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_HR_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_HR_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_HR_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_HR_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_PHY_CLK_FREQ_PARAM" value="0.0" />
// Retrieval info: 	<generic name="PLL_AFI_PHY_CLK_FREQ_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_AFI_PHY_CLK_PHASE_PS_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_PHY_CLK_PHASE_PS_SIM_STR_PARAM" value="" />
// Retrieval info: 	<generic name="PLL_AFI_PHY_CLK_MULT_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_AFI_PHY_CLK_DIV_PARAM" value="0" />
// Retrieval info: 	<generic name="PLL_CLK_PARAM_VALID" value="false" />
// Retrieval info: 	<generic name="ENABLE_EXTRA_REPORTING" value="false" />
// Retrieval info: 	<generic name="NUM_EXTRA_REPORT_PATH" value="10" />
// Retrieval info: 	<generic name="ENABLE_ISS_PROBES" value="false" />
// Retrieval info: 	<generic name="CALIB_REG_WIDTH" value="8" />
// Retrieval info: 	<generic name="USE_SEQUENCER_BFM" value="false" />
// Retrieval info: 	<generic name="PLL_SHARING_MODE" value="Slave" />
// Retrieval info: 	<generic name="NUM_PLL_SHARING_INTERFACES" value="1" />
// Retrieval info: 	<generic name="EXPORT_AFI_HALF_CLK" value="false" />
// Retrieval info: 	<generic name="ABSTRACT_REAL_COMPARE_TEST" value="false" />
// Retrieval info: 	<generic name="INCLUDE_BOARD_DELAY_MODEL" value="false" />
// Retrieval info: 	<generic name="INCLUDE_MULTIRANK_BOARD_DELAY_MODEL" value="false" />
// Retrieval info: 	<generic name="USE_FAKE_PHY" value="false" />
// Retrieval info: 	<generic name="FORCE_MAX_LATENCY_COUNT_WIDTH" value="0" />
// Retrieval info: 	<generic name="ENABLE_NON_DESTRUCTIVE_CALIB" value="false" />
// Retrieval info: 	<generic name="FIX_READ_LATENCY" value="8" />
// Retrieval info: 	<generic name="ENABLE_DELAY_CHAIN_WRITE" value="false" />
// Retrieval info: 	<generic name="TRACKING_ERROR_TEST" value="false" />
// Retrieval info: 	<generic name="TRACKING_WATCH_TEST" value="false" />
// Retrieval info: 	<generic name="MARGIN_VARIATION_TEST" value="false" />
// Retrieval info: 	<generic name="AC_ROM_USER_ADD_0" value="0_0000_0000_0000" />
// Retrieval info: 	<generic name="AC_ROM_USER_ADD_1" value="0_0000_0000_1000" />
// Retrieval info: 	<generic name="TREFI" value="35100" />
// Retrieval info: 	<generic name="REFRESH_INTERVAL" value="15000" />
// Retrieval info: 	<generic name="ENABLE_NON_DES_CAL_TEST" value="false" />
// Retrieval info: 	<generic name="TRFC" value="350" />
// Retrieval info: 	<generic name="ENABLE_NON_DES_CAL" value="false" />
// Retrieval info: 	<generic name="EXTRA_SETTINGS" value="" />
// Retrieval info: 	<generic name="MEM_DEVICE" value="MISSING_MODEL" />
// Retrieval info: 	<generic name="FORCE_SYNTHESIS_LANGUAGE" value="" />
// Retrieval info: 	<generic name="AFI_DEBUG_INFO_WIDTH" value="32" />
// Retrieval info: 	<generic name="ADVERTIZE_SEQUENCER_SW_BUILD_FILES" value="false" />
// Retrieval info: 	<generic name="PHY_ONLY" value="false" />
// Retrieval info: 	<generic name="COMMAND_PHASE" value="0" />
// Retrieval info: 	<generic name="MEM_CK_PHASE" value="0.0" />
// Retrieval info: 	<generic name="P2C_READ_CLOCK_ADD_PHASE" value="0.0" />
// Retrieval info: 	<generic name="C2P_WRITE_CLOCK_ADD_PHASE" value="0.0" />
// Retrieval info: 	<generic name="ACV_PHY_CLK_ADD_FR_PHASE" value="0.0" />
// Retrieval info: 	<generic name="IO_STANDARD" value="1.8-V HSTL" />
// Retrieval info: 	<generic name="HCX_COMPAT_MODE" value="false" />
// Retrieval info: 	<generic name="PLL_LOCATION" value="Top_Bottom" />
// Retrieval info: 	<generic name="SEQUENCER_TYPE" value="NIOS" />
// Retrieval info: 	<generic name="SKIP_MEM_INIT" value="true" />
// Retrieval info: 	<generic name="CALIBRATION_MODE" value="Full" />
// Retrieval info: 	<generic name="MEM_IF_DM_PINS_EN" value="true" />
// Retrieval info: 	<generic name="MEM_IF_DQSN_EN" value="true" />
// Retrieval info: 	<generic name="MEM_LEVELING" value="false" />
// Retrieval info: 	<generic name="READ_DQ_DQS_CLOCK_SOURCE" value="DQS_BUS" />
// Retrieval info: 	<generic name="DQ_INPUT_REG_USE_CLKN" value="true" />
// Retrieval info: 	<generic name="DQS_DQSN_MODE" value="COMPLEMENTARY" />
// Retrieval info: 	<generic name="READ_FIFO_SIZE" value="8" />
// Retrieval info: 	<generic name="NIOS_ROM_DATA_WIDTH" value="32" />
// Retrieval info: 	<generic name="PHY_CSR_ENABLED" value="false" />
// Retrieval info: 	<generic name="MAX10_RTL_SEQ" value="false" />
// Retrieval info: 	<generic name="TIMING_BOARD_AC_EYE_REDUCTION_SU" value="0" />
// Retrieval info: 	<generic name="TIMING_BOARD_AC_EYE_REDUCTION_H" value="0" />
// Retrieval info: 	<generic name="TIMING_BOARD_DQ_EYE_REDUCTION" value="0" />
// Retrieval info: 	<generic name="TIMING_BOARD_DELTA_DQS_ARRIVAL_TIME" value="0" />
// Retrieval info: 	<generic name="TIMING_BOARD_READ_DQ_EYE_REDUCTION" value="0.0" />
// Retrieval info: 	<generic name="TIMING_BOARD_DELTA_READ_DQS_ARRIVAL_TIME" value="0.0" />
// Retrieval info: 	<generic name="PACKAGE_DESKEW" value="true" />
// Retrieval info: 	<generic name="AC_PACKAGE_DESKEW" value="true" />
// Retrieval info: 	<generic name="TIMING_BOARD_SKEW_BETWEEN_DIMMS" value="0" />
// Retrieval info: 	<generic name="TIMING_BOARD_SKEW_WITHIN_K" value="23" />
// Retrieval info: 	<generic name="TIMING_BOARD_SKEW_WITHIN_CQ" value="20" />
// Retrieval info: 	<generic name="TIMING_BOARD_SKEW_BETWEEN_DQS" value="20" />
// Retrieval info: 	<generic name="TIMING_ADDR_CTRL_SKEW" value="36" />
// Retrieval info: 	<generic name="TIMING_BOARD_AC_TO_CK_SKEW" value="8" />
// Retrieval info: 	<generic name="TIMING_BOARD_DATA_TO_K_SKEW" value="10" />
// Retrieval info: 	<generic name="TIMING_BOARD_DATA_TO_CQ_SKEW" value="8" />
// Retrieval info: 	<generic name="TIMING_BOARD_SKEW" value="20" />
// Retrieval info: 	<generic name="USER_DEBUG_LEVEL" value="0" />
// Retrieval info: 	<generic name="RATE" value="Half" />
// Retrieval info: 	<generic name="MEM_CLK_FREQ" value="550.0" />
// Retrieval info: 	<generic name="USE_MEM_CLK_FREQ" value="false" />
// Retrieval info: 	<generic name="FORCE_DQS_TRACKING" value="AUTO" />
// Retrieval info: 	<generic name="FORCE_SHADOW_REGS" value="AUTO" />
// Retrieval info: 	<generic name="MRS_MIRROR_PING_PONG_ATSO" value="false" />
// Retrieval info: 	<generic name="DLL_SHARING_MODE" value="Slave" />
// Retrieval info: 	<generic name="NUM_DLL_SHARING_INTERFACES" value="1" />
// Retrieval info: 	<generic name="OCT_SHARING_MODE" value="Slave" />
// Retrieval info: 	<generic name="NUM_OCT_SHARING_INTERFACES" value="1" />
// Retrieval info: 	<generic name="ENABLE_EXPORT_SEQ_DEBUG_BRIDGE" value="false" />
// Retrieval info: 	<generic name="CORE_DEBUG_CONNECTION" value="EXPORT" />
// Retrieval info: 	<generic name="ADD_EXTERNAL_SEQ_DEBUG_NIOS" value="false" />
// Retrieval info: 	<generic name="ED_EXPORT_SEQ_DEBUG" value="false" />
// Retrieval info: 	<generic name="ADD_EFFICIENCY_MONITOR" value="false" />
// Retrieval info: 	<generic name="AUTO_DEVICE" value="5SEE9F45C2" />
// Retrieval info: 	<generic name="AUTO_DEVICE_SPEEDGRADE" value="2_H2" />
// Retrieval info: </instance>
// IPFS_FILES : NONE
