// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:15 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GC2QfIkCUTaIH4z7gnFnTZ/Swo0sgpHl+5QUo4ani2CQVyajJZvc1+kY0KuHcewW
0myInHl4AtDU7vTBFkFbWiBKMvCX9lfCRq7GY+K59XzQKWenlUWF5wHNkgeX6KtF
HAIWDYmWM5VLSZ151o5WxG0NLzwaV+RlH5nUpjVIZSo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12352)
aDcEc5UocFrgIGlosV3WcN5Z21wNnTGyWBV0mZBDnOx+gFupCZxrlhqwPjf10vOC
oZkcdEhXrgCoEyi40IJK+sMHC6rKAAtMtLoq1G0p3PHrYe91LIpjzFIhU/8eI5bE
l2zf6ecipurAqgkXH2dLNd/DC2+AaEMAmUAdj/s7t4G0NIzFvrjEQSfUYwSmftjv
8AwZrTs0BzPFfu7ohwVyYG3Cf6EAlGm6tA4pxpOjcRAskRjidaDgh0SzbAlWjqeG
C4ndmJk4cMnGptdj9/ad2DobTz8XBdoF5fzIq6KwRsgIYZV3dj7n1XNq802ZB2bR
G68To79MBEvFUEBbHpjZYGmBTZ3Q4bK6CKEB+lDLlV/DlsQ4F3ulkB/4Q/irpRw1
+VU7DMP9WyjadzcpYABux5mTLz9IUG+ineMU/c/aHbnExJ3ukf4sKeSNDb/wpH4s
nIc0PWSMoQOueHJet+fungbjk3sWGLSAZz6gjAaKYlKveoNKdGJ9pGVmKe3Fd6ME
HpYbJfYwZ70vJ3h1nKResr8bewn+WRsgBaTf+fOZuwwXqoTk3BubVG/DBYioeUGE
JgmnFN+MWfgVVy0Gu7bPRLM9wPlfilGgLCKAZC09cxPK5vzSLfou0W+5Ma4pacpA
trmZzitesPv168Go5NGjTw1N0wy4uWMiyHK2CnqJdaNTyv0GbNRt0dhD8EVUlcEV
Yl2rG1zI5xSP9ZZgue8e1PulLF9zreuue06a1sBEZC3OSN1yrGvUyxtsnqEhGjEE
2uOlq7HMj5aeCofJJn8bixhWmVBBefQPILP7RAffUwjwkTwWqjYfxTD14ZiGw3rR
5Wf2zZHhuvAzDUzHMJAXWNFA3EJxqln+P0mmwpEs9RCOJtLg+1m0NIQ0tAmGjzyW
CqzN0y8uEWOrr09KFWuKA6ZtZ7XR15onovmXKAYT9TkJ0usbLOHN99SVatboJYpw
CLVnYDOHV0aPdWw3atA+fSrGO48r397NJ6ehPjCuff2o6Pnhnv0SKVuKblhOZjVM
FHf+Sul6jLYUaPS0AiGD6J/+7OLzIa+TVuuBCgIa/OjxhyQNMraNbrbNiF7zTjVb
PG77ec3GQkvEoW7AV7XvPIj589gmJe4KfJ1txVQPZiR65B6QNkucR/NXWD6YE7kV
9qacPbobZDKQevqqkKdkCSJxwBsQNMqalB2BHPSI8gAMcV6T9DKX4k2A1K1MbGkk
cvD6W45YnHCBK5WkIPuyYLk1iakYHpo9BYGDsyeerjKwKyM8NYEkZxaP+nb6do1P
S1k2VeRNy6Z/eoLOxTNS79lgQA4G2+LoMVxgeTILVU/xfpXX4/hqv7wvmlkWgugU
fIQD/8xROjs2XBH51BN9tOgIh3vcTCaksyXJZ5puHSy6TDutN4/Hts8OIaGKfktF
h5fuY56qMp6rwfgCIKbdphvJzfoqumNM7JoL5LKAXl/NWwSSyHpSmb1bE7Jt5FQv
QbX2Cjz669Avbiw1axd4nFyq+W7PynssJ6OR6uHDGym9glQQGpDisL179QoBP/eN
vtloIUdqXJUivp5iAeTb9CAw6rMrlmetJEqPW3nsnbtJC7+mXJZfZicGe53vDQHA
CS3nsYlIQ/PleDZiaH9r1n82IdBd7wx1SEHg9dAfQ3JexW7+UtGeoVGOdtHEIRuW
q05wAXvkXkdsQljJRNbp+rNrnuAFNRTcjw6onsgW4liT1UrxStibBZDSADdkfF7V
6SrfGkCVbObYnKFxooQzCqpelawWNTPzB1/w2zv+oy3bt905ijOSys5qmhKPegmF
vB/tqAouTF53DByQZP/JHNQtFMym0cupWJoCvSCfysHgvriyBLMligmNngHcYHr5
wwlBNCwIple3J2XIydESoxg4h1x+0ckviOC1sHPUtJ4xh49IyrKG7Ixvk0peDSlp
rUuVB//XG8oLxx8KIpmfDjPQBHz0eVswUl0dAmB+uW5aL7eJ4UqLUZAugAh2abkJ
fCo8ow6Kg+gbVXuoKRW00zotIglhM0moG34PaQpbxJnx27kUwle9PopE3ygh48P5
DYorAoHqwDFo9OCiJG3vj/+JXqLlJ8/EjS2RzR5VCjpCwLG5ZOVjvmebuBh2OVnv
pQHnjcCpJ8fTQ7DinhMf8VAWPv9UBEK24wrtizfE/KZIRQw+ryDMJr7zFlxr6xkP
u0kIG/56vmF/jXzpXKd5Dx1WPvIsa+2qUwfjqi2lTS2dC5nLUjWcDpIuWLWuYI92
LsikPrz/wZleiF4fKMBsu3co/wsv/w3bqqS3qwZSKDCm5WdLlopWTKpFV3bAih+e
VvORCprOGaZSgg2z/7cSIeI1RRV4nc5cDJjOcc8Wx9BEDy9FILrx+TlkofVJYB0f
rLEqhW73OvpbJV7KW+DyO88h9Xe+omkdvbIymOU4GzVZfjjztZwxf4ZPn3Bx0MYm
uzLtTkf/KhtrCbwbxXs4igk2/6GODUwHr99xpLnRE/RpwEM6btsMe/N7p81Qm0TC
GACDqJ8pNp2zzhCI7BvnHznSgJVjn1WnG7WzRyDmx3LdH4bukRPAvILHvANyjoXh
IPKonzHDRj0wdlHX70m9WL+upVegT0Lhob9YTQI77wEwjKemYStMbpcQk4UFJnrS
fm7Q5nId6HtcoIOrlbW5LyKPUZOvz4+LxUsrPG5qknET9bsddIloj58oLak6sju6
ccw/Bx6KLoyjl1eer7ke1+iPY7OKq/HW7/GOZoW0s2eTo1eIAUoXW7gjqx2QdPiW
HZ9CkHyZBFfq0TTJWk9OK+/gIH6+C+PCVwlLsiMnm4iNEQL+6OHnok+ItjvU0+Mv
Cxxm9oVMCsx3bughSEDly8JX+GOcsrvY2Av+nQpWtNUHKU9IfDDkE2kFm97umvo8
1tQlthylEUggIPUrkajH+4V/mvjVeBMs7WRi4ekLvYr6Jn9G3M8atQ55GRSVtKMX
VfPSA0q5MWYVzDYlGiiGC+BmznZ203cQ0Q7KxjGVRxsFJ+dzjmVwBgz6Y02Bw/Ym
S2wys0eIA57HbuRN3WfOD6Saw9u9VnJ2339mFpJAFEwryGq+42afCpKDyiW7H9t3
5Ts6RbllexArIAo/zJpRgwRZZwj2Ciry3Hsv+Da54i6JJ+LTMvWIzCynYBUr/PHS
elZIoQoAm7QUDvJVw9pbAAyFEK10Q2/3UuvM/5ivpMEwrBty9TykMcwigDyxRuLy
IlGQXEOFGqkMO2n4OVWUfLiBHa4dgAbN+y2myP1eC0RjIjj6DEn1vlnuAO0adGec
LXV+kLjNlZ8+V/iDYgWN1GmdE5flIz37IzahA9u4pb6zuWFd3B6Us/pKhezKge8u
Om04j+zszUFrRWlQMpsk358mlGnLTToICSOzRzRq2QoIlxB3cOg2xfimQR+kEQV4
BLcTxkgqcMqvFmfC4cVzQ61dxlx92pwsHSUk80/ZxGgNJaq3BUVARgpSnPpheOz4
UJqFar6HKolhAzsuDHlZhBcIDqEHP+eJiXRzemjRv6QlrnIbs2eYNpfxnkeMVOSM
YjSojUQSdNil1Eyt2NLgo6/84AVzWoT7tatoPd9mr8NE1n9okIp00HIOywluezd1
eI9HkggtMTVE81bZ0OhC0tHWS9i4NNPIKOhC6aFAhZutovhxPO3/LIeAm9B6Ve6H
rAg1rD0cGWgz7vsl9t/3b1PeOrH1xw5pa7NR64aeCgoG3OijI9+Imt9wWCXxlwCH
Xn/1rikXwGluWaTGntwqkMqASlaJpNrZSX7q69dsjCYl4DFaE6hnBRhi2GiSvOTM
W2h3WRH2o4S8EHziex7OGu9Lqzbc6PD9foTeoy5ZW7fvojHezPiaNhLpZRL+EgD9
t35nbwkvwKKpIeXkOlrfbyE2abV0/LjJcrFp6sfLsOFBDyWU0SHF36UeGJbx1Eyp
Fa0m9Ol7prQdtj0CwRKMvIesp6gqMqLp/KlJOy1rVtEdQy2eTZYwYY5tzilUCZuX
lnABGx1J0NwmStw+qxdlPYYwCnmhX2JEXrbwzaR94hBR5IxG7J/JEyAR6c2W7sJW
w8pEWJfcKZIO1rv3rz3GZNb99uQ2KiIVv0xDm5eNj70h7rrFwjKSqhmwSxS+JuXy
hWsudRG+7o3HQmp+EGXm+cPov4RrBiZ6nSSGQtS3bf3S5i6DuiHwnu2+MOxHfmGJ
kRWBOTqVFTjRnp1rsnWVcvOl9loJhI2iw9w+l5MvsEvgBoFgyUbLXjyOsGQDq7Yz
auvrq3yXsiGk2YiaJejtOWrap4QUjhaYY42N2f3E3ltYxYtQ0u9WfXBfirYJOCN2
0SJA5kkIoQw6GYVfj3fZgGFWzTTXklxtvAY4Dd0/EP0X++3Jdj14QsOj0L0zXPQV
T58DGKIFytQ1B9KQpD9fwubRNaVQFiCxEHNOMhqUiGRhfrEsyfl2q4sI3hzOE9x3
gbfrlGf/VTaRZOGmWHQY3umMGn8KjR+Ym9wBj630eWZ747jb/AyJ5pMiwxm/GPKG
muv1NAz4neaskR+tHBqFc4Mckt2qn2L7H9kWmBgOc3QLgpILQVKDSmU2SReaXYKA
HvBdH65q4I7vS8sFTJPi9tsCjLC0hscNpea75DZ4+tpuopfbi4c/69Bs35P6pD94
3eD8cuDG4/DLh3pSC7O8Pezni0nrsYuNX9MmfG+NoK6eiXXOfTnWBMnHNm/JB84R
esKI/gH/0o+25fdMlo1OR+bI71sBOJAPyUC4YEeR6ZaWtjOPwHOO3vRD/E3qoj7V
T1VHfhWaA6lk0mg5RkgvM1XuDXcTwcrXxBezh0LCGNP8OA634C2lXC19NXsSH6p8
P4jfU0nyHwPNBh5DO2GYM5GbYstMz8KXvTzdGSe4mNuov254tevhNWxmy57mWFmW
WlB7vkLrz3nV1rUX5fl5z95ZLivgNtEexesqjeFBLohKbwMsnsitRjeqm9fZGiQI
M5DA1Kayn0gAV5qpNR0LIVgkjUvsbQHrQKz04XS4IS+cb5yx9Mzo8lW1gz9zfGvT
tIEXmvvwa60OM/rRGrScB/6VpPlrulg8otvg77UHqpKC4cUVvxmgd+LjPyr29Fgg
JjVePGQZ3YxZG1OrzS0GtE1ZgYUcFxcwouPCw3YGVcVW0adPgPxL+VPkWaZHfLoZ
36Wmdr4rL9X5k84t0IMX2jdFl5/ZJYVSEMknZ49QsB8/uVQTkZkgA5D6z9Asb9x6
+gGcVsoQ4mx//Oo8GsmIJfAmL8pUMH30C3tH1Xf/8kQzlrw1JH+AGVswaVDW2Iju
2emQJA35YpkW19H0WpyzAL5zgAr2jsmhoF5p1Gs4hCTyN+OXjH7Rm0w7Tyovccjm
iVutr3UpdXfHpR85WjeXRRgKxup18tMy4A8kydrwrnnxBYrIJVKrxCbf2WiLfeKn
SSX3a1DI1XDGKFInnELZhYWZq3vuxH+VMjWTGCKA/BYbpxiuX5ksbozN0YbHew4D
gRVl66tpvC7nh1eJ5S/+dHseTFviCndDivDFxvZ4rQJQoTy1V+nw9IkkJSjm9cS2
JCMvQM441EpIUwC00TxIDCfUuMn+W5bq3r5ysTgK6rMy3myaD8mjKrMzEK5JXQIW
tdM+JiwUmn4wCNyu88EmKd7i6K8s3Foaskvj98uUTqJ0SEM1rVBXN/L5IfQXnV0a
7FcbFJT9k7AfVd5ywezk6dU7R24fLLsjQ9DDXzXLSRgncWPcRl1mfShlYd1waoJv
CUe0+7C0B2lPBtA2aeKv5xVdH5nhyJv/iY81GfH8aJxg7G3NO+Uyy4XCTiuQTqKB
AEs2/OolyEZhOfO2GGSq334iGIVbj6DRiHY//WAIx7z8iF+pQocbG8HKG8jzmtW7
xXH8arp+eX+92aKojF6sRtkE/72QhH4LCp8wmniRDPSSeMA5Jv+B0FAtfCOdC7FC
mfp+xVjxCZQ2YtbdLN8DZHF20DpRjF1Zn3QRjJc4+TlGpANBSZNhThqvX7ED8Tj7
6GEWwSpVpUMIMfHLuFUSgi5OK7vxM9t+L/BEm2LQtoHBW5hUDW4iBl7UbGfYhRwZ
98temurcAL/CwBg7j1AJCP/j2WdqtCqL+vm3K118LvGzzngImIjDiiyWd/GlOhim
SciW/11z57QYq5YqEZ2K0wfD8ADiv0N+Hv69OsDxnEZXqkm907XR70FNL51CRyds
81XBwwV+HE8sTIp4to1Sx42ktN2YhrwjnJry8VCoJXM64SIk+BrHwkxVLOhDct0B
J+flwm0EaCdYej5uXrSa6+1fTf5F6N81Q/IkIFWqohMp4BkhptIJb1V5sMYFfPT9
o6yyWhISi4VlkobtyD5uL1F0qiOzTvnbjQsUdCWY7H3+tm3inpmoYz7I/8xE2uCt
NsGcprbE2NgQDjbT9mPBnTiQwZHDK8NM2aApIB1WoNSPQJLLzii1kDMHvRfQupKM
kYlOUrNSGpGCoAzMQb9HyEwxuN/KPEXoKHaGJ1KmZnrwwQ6J3NXB6e/cXpQQONFe
Hz+pqTfMHaFDb/skIWqpzI8Pks+tSMaIL73ILmyCQ9veQ20oIUePMH3sTgxNN2qE
4REEx+B593cTnqbWBwZQgoyGN2uKJaVB0OVpSaOxawXr4VJgw8rH5z6Ch5Lmhe3G
Vx7lMS7xpUABebpI6iDzo4fZqvWO7Prsenit/iBx8xpWawrhNIHMW5FjcDJRhzls
J7VfIpzLI98bJ88t6wR03gWuk8WbKeF42ZQaCKOcBX+hcojgsi55q2wftu70J4Wo
1eWv2d+EdbqCJ2bfZZcRW74LFsq1T6Yh3rL61vAqsNmaETXuRB13NVOnkgOPTe/S
W4yO086uY5DnHYwKmtsgLVdawZC6KAmfIrnPdsS50Zxa73U2gujQcnBlGl43fZj9
SbHPBulAiw0TxqOQwVndJKO91GcrrkPkMbq/UE0T6e8jpOA5Bqjp2iIe2b4C2X8t
lZYcYX36DTh5xLoVrPqyXqRvxZNz4DL3yjAuxJop+N7SA/i1W+9NZKq9COqUSJK0
GQ/fj97z7DivbSML+OzjK29kFR24eA/emAy+hLmIVXgT3BBcH5znb1HmSkgJQPBw
aTDU+9W0SwMv7kxHQW79/qK+St0+SlRyUivhK6XWwsBM8PtTEPoMGM5WSLil8JXn
bxFC3L3+PLwQLF9cl2WSF0apmF4xIjENGQA589ILo3Wq9S6Nc65fFbr5sY0/ipIb
/by+jW4XVL9a7HtTcpbbifyp63tBadP/S7hRgM+Ofhh9WZFcytjBabFPLEWvPqSX
AC9fGvrK65IGy1qkZw72FbgHetxEoyfaCvepERB/v6t2GOKcmtLuTbaTqjGb56+X
vWHMXqNki07yffsDu+r99Uq+TUyQCyzA0i59EIG+8MYAJKb3wZ1TvBy8cWPG66Rs
0DcXa7GkcVSIEltFvOFb818j0oz1hz9o+PVCaRGLNz68vxa+W4wpBBysBQ686CaQ
uEmCfNWhv5/vT9Y7yc2P0lZuY55A6sVAlM6u4aVr/Wkj1+6qfUcFK40Vga92a3bx
+Y3IRWKNAhd4wmT0CAd/dtyhkZd21t1xbqtqKDea8Liq0Y8y31xJSEFbpudH1c2H
OqIG4BDbaUzHDEVsB6ckmsSCP3IpWwtk17lMlqfqpEs+vH0GywT8SEoGhADhCJ4o
vi16+GzFVNfdEyIlCA8XWjpNlWexhQpgO68SkSU839Zca550SFcB71+6iaOxYNj7
eyHonYTZ6W99omm99otmnKIadNhZiuK7PZeBwCKjGJSQ65kRq3iyS8kC7D3vmso3
VVCorG7C7p43VvXn2Px5VsdoBHwHN91cx57Yr6mzDlIAfkw1AWYXbeJce4lCcE2i
UzTtsge8mzgnQbMkLYQDYIh9VujlSO50o2T1W3F/P3awnZgD9lt/mhrKxJ6Afl4/
5jpwYS4lZSjZcucH2MYsrMb2nw0c83y5H6BLW/BbwIBV0XkrvvuT8VmvqjldLLB/
l4zPkracDyhTQBS1DIM21r/pprxO1D5UsS1jUgYxDfmKHxLonVhDj1plyJLhZBbd
MhNUjnBFDFn7DOPh00Uy5IMdDtvid4qe86Yy3Ums0Om39a8Ye2JdqusrcO9Yo4dE
zDbXB+dMUVGwXFue1cYbpIj/TYHuWOuQOKQVE42Qxdl0RUHdFr2aOUNQeZWtP4zF
8yjydvTtWOIjWNwijxUhyNumB24ICHVHiZJpqZ1bZyIqDwyCUX5r2IcR6FV7yC9/
qMRHUh8iEDsTRwxEbu2nRFldP4/7K0KudoUQidvC+5kvS+7qT2oedH5lqYDPLYCA
7Fg/P7O8Y3B4+sSG2prq/+4G301YhrlgWA1NBkikrue90HdHwDaXrcpCRjGVFAmC
+JPC8eu/m+78KhCqgKZ21iSVqYMhwRMPKgxr3BjtLUAxxzXDP/pG99h6asgoGxVM
cX1P/Mn0jkQRKBOfoxsVzGJi2z5YY2jyCBoof8LHFRpwqbk9inEKRmqZ7g+IiEia
Cl7hINxgOk1fha7btDWJ4ovb4i6DmgBcpRInNwXZACRcH0AsPJJWHf/P1CLCyBOI
r7JkOW64pW7aig64rjALsTeWbjDQBBdd8KTceEEcmrzZa9fizi459tN9hmum5rts
HTMRIuCfRCyTJdoV7Gqql4NnamNBVdfJV9n3bGOZUZ5jAK0mP3c2sFjLyl+Nvph+
n8S3QDBiV+NcNIiZtkgEL+oSwywiFFjjvH/L8qkvMyaD9YhtJrByeWzLUpEZXxni
GRmAZd8iaGTd6QBiYqFbbnWQMIAeDWTgzUELt7h+NCyRoI0qNTnNoKmD+3Kwe3fo
ZyDmGrFnHhvR0mpyzDSRF1er5eqm+PKQNggbrrGNl19xj4UrfYdRtySZZ02HlYnl
5+5IGqKY84zMOKnKZzdL+I1ImLCtjTD/zCCGHp6XtvMWn+01oLpzP18Vu/Q/bo3n
i0X4lfOpy78PhtIVztVgYFOYSe9WFR+GSkTnyZO7phgOJAC2bItBlpMTwTasbRwX
2aKy2Q+tVvzprO7xm6KwzePnAxjJaPzKo2GHdBXdTRKjpe/BAllOZKIXYYfXFMcU
Rz4+zKMtQ2tfyLz7O2bvxqInKII8gP6FHcbWkKaIZuRO8O6xBjB85BX1H44kBQXQ
izss167MJh58T7WXULm2S0jLidx45b4E+gpFBwKFnYtV4xR/H+gQmtQOBgiVMXDi
urwZeb1mXV5pcCfW9EkNkEgLCPIwM9CtQr0H/rQaTfP6gkzFg6HiFxk0WJrpdvp4
Z3VDK9gEB//QFxNoiqbmG54HbLHywTNHb2bCwHaBKKupROkCBNt5CUpBY2jUQ5bU
a7RZU5APyM/L8rACaJYlvmElqlN2Az/5AxqYDu8GAOuFaKcpwChnyZ43cxV+pzez
rFPYDa8hs5UOScJvewp+oex5pcfeRnhGAxr+ey2k+fr5lt8VwX8a2QR/q/TYahBa
ip7PG+jheicQQzvYU0z22BAfuNYUXnSvxDqGwAaJoBbgoRsNcetG5UdCH7aYaZhe
gZ5PF3z3txGN9p639pANVD2QB07IWD89FhuMXpVtjAcWfFW9L/qYFK7M0F+CYdBg
uU/uAKJ7M9bjSyF3XLQLQQGjSmRiacHdwONhN7K57KJmOcHvPkD/SEOSRQERrYGb
hroXoWd2GbjcoXb67kG0ZydlCC/PT0qrswS76i5NrWFmVaVtjRpfHr+5ZUFSopuw
jStCwp3YnnltT36RRmkIP7g/kcLyDvtTd699L8v+AoUVwbO2sOMeEUeudh+w/bgV
nk9atZC+tU9rg6vmbWGW2/bFkjitM5nPKkvsTzpZ/ChFCFEcsvVtVrZhck04lgUV
KKg93LdBdKnCJ7x3JQH11r+wSFXhPkLewlRgN745PucU4jXP5jS1JTjroh3FCzob
42FSCO4aAP2hU1bFoKXiXuwc+CfsMAEfoSf6ectWBNE248+IN7Kjx6wp0YK1FHiG
RlspEHaHSGsd2RBT3dZ4hfgVxjTMv8WBOGyCqqC7dx/nm7Jns5XncAjfJHIbzHSd
S50r5CEXDOSJqjkmdtrahA1TfexVDGPOXQ4Zm5zmLbmtz8L0CX1sZtfzGC7owwZg
R1mS/WxuOn4kbb5dCVbNd7aiXd4Mfo13vAF3jO9x/uZwpX59KdQ0quh5Ps2GRR2B
q3JuZM71VEffySD87cpjqhoKaVDIBlaQbgTk5F9Rukw6g0IYNXB8qY7gYAkoWFM2
y6ttm1NijJJ8v0RY7MTfCsfWq+oFPQqek8jKI4enUcnCj+g85AIzgn3Prh064FNq
fOqDuaipCjziMO5RHyLoQq6perDE8NJwhmGTx2i9q/zEjqCPdewMTK+yEQY/UlCP
BprrgqUArRsFWXBGs9mc6GDqY9HP0YquGhvShxV7DHFhZK5HXKtqb+JWwoyT1BHe
FZcT1o+sfhod+LYW+VkPB/v+E+Q0na2HYPsZQGvyABHtzNscbgnwED0yxHbuCp99
XPW9D4HA1MxYU/K4cMxGoqBFTLH2F1gq6HOf7sxfCTE7ArJe7dG8pfBwyE0hXyk+
XINjWG4Pw4rZKkZinr/lhqrc4w0H/8ig6Y3u/CDPkNGE7PoquXKhar3gif2nyp28
Fp3g1fKULPIAIP+LyLFZNKZGTJecTxY7f/WyL/Jw36IWhdmkqaY8RZ1sXnspjg5H
uy8JY0cbF/1c63PJfBpQQ3D2NmYtYGVLOyf2FNYYgJQ1+SdQgwlUz2gaaOuD6k7h
aQf7RUAFYLjIxlsEMuZTiUOV1g06BA7aPaBGBZKvhWnPTirxQ2fVCCyXYlOXqBcd
aYmWOzyY0aUhd+onP+8Q+dTO7nayN6qBag87KPmyCKExYiDUMlF+lBZW4iHy2EyD
Ha8Y+F9+qKyKhH8elwRZN5MdBqlL6+aKwIQPGdv1IFtbwGlmnIKdbuT/RZ28OKgP
N4OWvmeqyhWTEdNKSa/zfMbT3F+TNIsRsx/ovBN5PDgZZfmqGWYLPrWEpsiP3rLs
U38rNb4H+uUz7RELN4dSOyz/5MJq76l92hPxm9Gynt70YG52QN6KAEQZAt8TyvSr
ctTk72pX8SVl8QVFC9zGciZd//ADtGrsH1KoMAp+d07wJXsLt6nf4L63uUDO12rD
eD8ZIK2ccPW6Ld8UoKYKozoF+azl4bql5zigooe+ZLLjDNaC7Gts8aG71n4SLQ0h
VKigwxc2mxNPp4Z4dAFTb+HtmItYI23q7m2HfPnHkb6g3VvNvlMBwn8RUuzvIiyC
AaMZtw73fmdj53ntQpr7OhAwYRwHadcl5UwOoatb2xZe0RAKc1BJCR7hj3iSpf41
wCimQ5eOckhQYPpxmtzdhM86cHlYtf4CCHkMgFRrbEpTd7OXXA3CIQTNcHy9GiZ9
oYCN2w9LlI5BxUgSetKLDbZJblqTcPnDSiq5YtwnbmR6CuuaYrCkKYvWPC5dvngT
c6GBENpMiDY/2SqDsjzSEBcz/Pe6GsCRyUi80MYszE2l/emvb8/KOeIA3/iXvq9y
3mV6bdohNbvNMIyv+8ql2cwgP1R6g5m3BIyDW7TO5BryQlhdpiIicor/tmb6RgmH
h9ZvI85DjskEY9sn4iWAXZBDxVEgE1y4jB4zxmSgIs0t6qxpAuOWP29T1cmISpeP
Y4vyMLC9cSteLFgSeRlB2jrcw81jwHeQaIJqTTJ79SqZuM3SZ4YzdngqKN0P+/G0
d25XOQpsS2G4FRXlfe+YTJSTmFUHDeVMLuNy6fTSuMbFro6Sqiky0vy7WHTfHfE3
UDtrzoO26DVmhqhPnSwyZ0l52gV65mNNCdjjV8bPKK6xKBfUKULLXtgld2DDF+gE
K3sc6OsCSW5JT0c/8GncuSdka20ROVW2AlDz8VDsPkdy2rIvlZdCRYYUvzgUS2bl
ide5By3dn2IBawXc3AOSbmbpUJeu0M+4pNS9IFd+/rrthSQA/l8brTK48WXmhJmD
E1cmddPHC4KMUsbYjkj4ycyMG4Am60R0ypl+FShmMJMdOWRGpIGPKLEYrg+Kg7MS
RT138d4DkKjSG72XUhUu7+kChH14xM1FS0mr4OBN9lZaoXWGtF4UHpPBw24I3fzi
5D0tVrDap4nBB+FOsZqYGmiup7Qu3JnVJWhEyGHRSRnYGD3Pq5HpoAC+HUVQuaGw
5UwjCZ+Px6iGQ2ncGzHJ/GA1Zc1Eb76mAC+y0PM733wyjtH3PFdmSZ4xGjqiwDkF
KNwbJLVZHuiECsGAfHOxOAFVofP8NNYdDOt4ynFEjyY1hJOHMSyljcbpTEIsdpnY
FpZeAahcjpkNOLXLiO3eTXk9UGnW0/oP0iQFK1x5SzWvzPToGyqGnoTr7zj3pdKp
FZVd2yfSqWh+QP542W80g47+hiRkw6x8NPmaEdWkiALWMKTTjxiEETLVVPIONe5h
IYJzJIjkM+2twFeBDglSerZIEqwjyB9rXagmTXJJhXyatZyPNU/ZhPTGnn8EYw99
YPklxlmhn8u7l50BdLdFHBhtQ7JUg8B6JH8PcTC/YO4U3LGEQvdrSP3EzNxoFBa0
BascTG009PAZHjNdlpDS3Cavn0d0Uk3DXQqhUVRd4Im93dQDpzBnWDizIhV0oZk+
BhSUedSwmcAC0ANsfFITqKx/LOyIzx11thU3C/fe267Aq2XQWR8+doYfwkl6oitH
vM2rb/MRKFv/8TMDj6ot0We648imAgbVqZoGjwGeig6AmcRxZ4113et7RiG8Yuus
W3xazV5VXWyFBDILPDtzDpNNUb/gZNQftz3QPL60hgF8/kiWVrz22uZlcVvg1O0T
rnkwYl399PZVx55W5bS0DsgOpVCooXE8nIvq6243+7tRQM7ppGbqIEZ0YFA1mFXr
07TtlTiqRDfxJdeIOa0HLQgvUihLgoGXBpaUvteYCoO9hdU8meVSDyZUf0LFo+My
huJPwPKnC94o1Yhz2SDxB0S2FLwVj2hMPMTFJPVMZlcMWmcTXCWzLNiwLZgSS2jl
Jt940UdiBru+ZY6ILe4nd+ogNifcP1U1DxtFsRTHpZbYNMwcv0KOE+KFdsyKJWFz
lWKw9OY5maWUXgXcGUpa1QawGxcu6U3y1oKPYeQY3twBYdtzWrmGeqX7rbiDvexq
AP+7Mu9u3Bi7W82tDBGu2jCkqm/1D9miXP3uaEPpPSZwdhC/aaEZblvs2qoklF/V
MZlsxqpgu1Bm0uzgWvZXh1e2x5c8xlKkGoNtWpAGwSZ+eyQYGjuec5HwXeC7JFTq
unMBvTRMl+BsvryRfu2Bx460nhd5/NRhRqH2jBgWMXp0RdET6POQ4fpeqX7tF3KA
tbemWEtPoyrkGP58Plu5rq1ka/x4nSrmGRumwgFMNb6KW1fGdnqYIyx61ssNjGEt
TlzLySiiZqKDCmqIuto2xZjPz3NYXaL3SN4ORdtiBlH0LfPrlSsY9C0pbKm1jYud
FS1zYki3YlMbNPEa8hBgn0EpQOxpyt3wQGEHNGEzV0oMNiV8uEBp1E0W9Ytxok5X
2REhKLTlqnvyFDacMdiNvYGSJrkpaN6MC4BI6ZTNa0V8SXXHY+yIK2YbV6sKWjCl
kWDtCnXRGjJ3s79OnSrVAeSVps9O0LZ4PC30kaNTmHQs3TJvPujI990KNV+lAmXN
kkzMUn0bb9dP2nGfTkZJpy410oitCZAL/xGf8f42QErRHuEdS0VMQVSOdluzPQiG
tDiFCSltthj+oFIl3eWxJjw67pLWJuhprBbw+cLkLUa2DmEKKUAeQQ04Op3iVs+g
AecO9ANLGdodESjXIRtq/7WOvz9s6HMT7HxDwbjTYdBYGZILawBM7IUfma/3nUED
YuZt6eoZqxY7YrWZRka2F3D61jlotbN6HAJhjOEbhPkoe1PNV1vBnubFaVCgIW1V
X7XWUJXQkeCYGTc8NZYL2T3MfAFYFVQ+JO3Q0W7mYX/16WeXMWtp7mg61Ml/eMMI
XvCzd9yIXV3pz+DQug7n1tqTy2yOrKfACwc9ShOoXX0hK/iw2k+7M15jZ/Ldzuep
5WgyZug607TPvBS/CJhBM3VRAQoABdDm7st8AL2feTGC01MjNIrs14SNpw4fHht5
d/mZUo3szVhvBEnix/9lvhYLW+FmTrgZXVoe8wGu0atGYH/VgD8p+kg/qK1Q9wQz
rjl05EGMwPK4wTTqJ4JRuig31Laz/dwVz0sv6Hjx9ArREwXy2DMtjZU33WVVLV0A
pmqKrEpouIu2k0n8ng+UuD3pk1++Dh5ACwesc65Xqhsp6PXbaBheGSoMe0b1dctH
f4Lvu4CtipqprNVgvMExR3ukT73SYnJBPylnuC32g65XhX/uUGzvVk3gDQwNP0Y1
QjUWB+aWhV0TTBpS58P+cz4SDkXHjWyiBnVl+Tdi2Bzf5Rkuz6tfqV6GtByFMsqu
oHMF2zYRxU2p1pjyFHRRYtSZcRDuS66iHdmN/Sxx6wyuHroBCcLEaa3gj9If45uW
0Xrgb4A+AtyrIEajsHP4WBKvHAiaEf8DXpO0Af08+NzBMNx62YPhUXVzpGTQHZbi
ieOeYVcq2x+mZc+raSanjnldaBORbNP35iX6f40gWizq/j5i4aO/X0tr1CwdJB6o
Z9qfLrvUk6EH0DgwUXNWnmv0RcEqSUiuXZgDEYH171467NsDj/9UPNV5gjhCUK3N
lTa/qKlkkBrgoBF3Dn3SdjqQ7f+JQSyGcLIBM1h3lphj19yvTIi7RDOhtBc48YeF
DQp7kjk129Z8PkYZMF8pkEaFoEtgqT1ijwAjr/WGK5cqrm7ODns+IN+6KbYZae0Q
eCOsojrEHZN7xioNU/Nxvd3aNkqCisBfg0lpd+BD1eK6HFvPrzq8okVPu0y13w5q
pXEk1lgP6KtsNZMwFjR7XTHYeovJ8xGaiQJuSNKtEjvvg2a5iMazETcbJ/f3hT+t
iRel3mYwHr4uEkYCELmdRqz7nf1RCrMHGsYj1a7pLap4KWHpOVysawUspT/JPrvc
lg9FpergPxVt1AKhLXXe9TJBl3LB26nHVYSwUOz9xPxbEmInZsY1g2In5KHJRhSe
LRmvptWEwqgcNUFsfGWgfcvHcPQUhebkSyxv7sUmWluyCNQCrtwbtazPTFDup7HR
IVEfu0EhaNqJrydyOUbhJsQZhD1s3+XN+aRMAjW6h65ohJgz+8sKLLnAjZm/60Lr
U2qRNq77rp9UI8skH5maZlZ/TiOdRoeavWzqGxX9tRRXYxk+oilaNRgdynCOaX1C
qCQ1a+QBjU8/nx7UmX1GdE0RcNx9T2DH8AjWo6QFTp3B7fPZTnwWv1WbRS251Dx+
Aa5d9YGVxVyQVWtKLjGQdnv7GirQ4nIVjeUXU0GKK6ly2XOTwVAQekVGT6Pns/1z
++pa37Gc/0ttvGJIJwtoWB3wcR3LDP67dOR/a+l4we3Mnp2kt+akzxBxCNJuSWIQ
tMsBTDUwDD382SEmj275Ja+npnFMfVuenkgkWiLsxIv+Kw27ncmh73xt/Zbg4XSj
H+k1XRd2kPyArZpA3J+jGVKE3a/NV2xmtERECWGsA+HLiWqpckdd2FOASw1jJT1J
X9L/I9a7ucY8MyG8I0xrBggXrM90KHJ8jPeaCf2Io7aUUkmwWSmifzumSSX3sOgF
U71HI0+eaGyTuxif4fCdqCuXZhwNKutk3o7fRKvNsvxZhCmX6c81D9f9FGkkwb4R
xL3yJqhfeEJL6v2MCdyXQEJF9GBgjsiZZdD1lhjwWnqOaRY1vHHW6w+7WZSPTDr9
urxlwrNm1A6gQAZfoU2fhjymMrPA+xgfz/8REmMFtMhsfZRwA/1VNH52P9uSlvMX
TNi6PMMLTrq9nN6rDrLeDntanKX01131nwil1fPI9j90cVCQtWBaTx6BZscPBJYM
3Sb2SkXbJEXWJDQQWN08ZKb8af7pEdKCv6QuUWCjrHCfVlUBNVG3vUnGcPDEHqSP
V7gQI/VqZg6MX4eUeoWtyTCpe7S9rE1y1jzLYsbr+lt9ISqFEDvMe+5/2Tg2pJod
Qx/mFqVIqK3t5ERtugYLjMxF5jWpIIbEzkCQFK+qRfQGDatvil0I6CsZy5uxPMut
6KwSuG1LzW5U/vqolgoa3PlMz/Fuh/3D2ECMGXivhvDMEkKs2f5ZI6OHUUyLFJS/
brgs4YmpnhqRbIVUjFinB3miAgrNvdJyLKfhFd7/D1qZpeCbqLODVSQ7ezS+VodA
yHgHZnCfXYX51M1RctKNqRRKebNqS9oBfgEfPhqqF2uwDANZy5zpwsVoQoDfmHce
/0grb2QRdXAFDLX7E9zm/61sYWt2Fvgd5gUc0CQYbTqziUCkfTwIoA+j0g16RHZs
ERaSCTkJ11LAu2nuqbDMjQbW/ihaElQpKUll7pvZO/qY+vsm22yStlKB+F7KNhT9
7sjkiYftn/P8flma+NBBGgG5zrJgHDMusJ+LjQIg69zBOGVbbo1cF13fKxta0Okg
VYbB+zTmLVXuglNtpLysFa0TSYMsV1e1AwMYUQ90k3LRynY3ro6VG0Q/QTx/gwtE
tkl+F2cyRWsnaoTiFGGoxw==
`pragma protect end_protected
