//
// CPU TASKS TO CONTROL THE TESTBENCH UART
//
//this is a temporary solution

`include "iob_soc_conf.vh"
`include "iob_uart_swreg_def.vh"

//file seek macros
`define SEEK_SET 0
`define SEEK_CUR 1
`define SEEK_END 2

// 1-cycle write
task cpu_uartwrite;
   input [3:0]  cpu_address;
   input [31:0] cpu_data;
   input [5:0] nbits;
   reg [4:0] wstrb_int;
   static byte nbytes;
   begin
      nbytes = (nbits-1)/8;
      #1 uart_addr = cpu_address[3:2]; // use 32 bit address
      uart_avalid = 1;
      case (nbytes)
          0: wstrb_int = 4'b0001;
          1: wstrb_int = 4'b0011;
          default: wstrb_int = 4'b1111;
      endcase
      uart_wstrb = wstrb_int << (cpu_address[1:0]);
      uart_wdata = cpu_data << (cpu_address[1:0]*8);
      @ (posedge clk) #1 uart_wstrb = 0;
      uart_avalid = 0;
   end
endtask //cpu_uartwrite

// 2-cycle read
task cpu_uartread;
   input [3:0]   cpu_address;
   output [31:0] read_reg;
   begin
      #1 uart_addr = cpu_address[2]; // use 32 bit address
      uart_avalid = 1;
      @ (posedge clk) #1 
      read_reg = uart_rdata >> (cpu_address[1:0]*8);
      uart_avalid = 0;
   end
endtask

task cpu_inituart;
   begin
      //pulse reset uart
      cpu_uartwrite(`IOB_UART_SOFTRESET_ADDR, 1, `IOB_UART_SOFTRESET_W);
      cpu_uartwrite(`IOB_UART_SOFTRESET_ADDR, 0, `IOB_UART_SOFTRESET_W);
      //config uart div factor
      cpu_uartwrite(`IOB_UART_DIV_ADDR, `IOB_SOC_FREQ/`IOB_SOC_BAUD, `IOB_UART_DIV_W);
      //enable uart for receiving
      cpu_uartwrite(`IOB_UART_RXEN_ADDR, 1, `IOB_UART_RXEN_W);
      cpu_uartwrite(`IOB_UART_TXEN_ADDR, 1, `IOB_UART_TXEN_W);
   end
endtask
