// Data and address widths
`define NATIVEBRIDGEIF_DATA_W 32
`define NATIVEBRIDGEIF_ADDR_W 2
