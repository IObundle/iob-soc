// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:08 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W9lRhNGstiMAWtPmpOAwJhPXFf92uJtJgLYXtjvUo9XHhoGB2uhxPeLcB/p21xxM
8y/PL0g8YpcPOrY7u832pCv3TPd2OEdSlM/+5VhRj5sXLZ1AUsPET2UP7dmmKxGa
BMdf6T58SjyHH51aJWYBbd9/frEteE+k7hln6ryVnlM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3296)
2KPzLuDndVBRaoppTc5xbkSiIOzHlFxMtCMIMNOI5ie8mB7YJRdExuXgUsPR9Xcg
ypLPOEE1O5HgDCNMYYUrtiSJRyKM05UWePFGgIBktg80k8QREpdg/cNFH6VZGw1N
leMgI1dNg5iuvXEqIBTqwQaH7+B24cfNoR3tRR6lXhx1pBizFYSi+oMRUP/sHI1x
uYCPVoMyyNBMNXDC+RUPy757UCgyqgbL4iKensRDC0tsKsXKQBc8vbz+9YlQCTqt
81YPw8hIp4VK573gBQPhpfmBy7N19h2nBdREaY3R4TyTEbc7BQe9qhGRQIBOtkwr
07wbV4Ev7sakVYhIa6Rd04KtJIz1B4QY5iJbFaDb7+MyKyoNB6DMVdWexb0MZOjj
KI2Nu1RKFpfoYBKbMQZcq7VT2Hr5B/1tjhcTFoQAAN7ER92tf1mve+x0lQ+8gM1I
gehgkYgjNUXfJ7xMKx/MKC+LyPzsLMy5ER1ozXtZNTYI54BbBoMbDp2Xy7lAcQhP
2UXXD+M0gL9Tqkk9a3Lq+L4O+RVbPFeqvf5TQT1yVFTGzSK+5POJVmm4sqBiBljb
T0Z+Hnmx7nIrH1znZiOUElEPVj2YIBpK7yI4v4jp5ttnjOOswMVWAY/nlO3qQZIq
CEehsrXDYDkyzff555bZxSpw/cNViXUMlj7ttFSG7ApPPY6AOTNE/fUwhP8ti+Rr
ZsYoXnmLq8ZH6HHejLEFj9CXv2juULEpZ+RmBzaKBLTJTUrigJuFSaSfUFP0oY4U
q7FzvAk7w3Gz9ILZ+fEU2dmOp7VZqIjrrv3N0AkRWljBlqKDJPjc+D6QYBWNckx8
Wl9+0q7aT8CRqN4m+Y9kzS60TAImWdgO+noV5ptCinM73sd4ov8Yw9ZSZJnOfKbx
fu/ElBttRJ/adR6T0GygJyNb3XsTSbxG1OlxeZ04vVfPIlHbXHPmiZbWT4/p5cLn
Gt0a9csAtlE+672h+JlbDYMWnQflcOGCp0RBoc34n1L9cwjXoTkaRmgtlRQIoOe5
zrIQy1S28Tnc8bM1JQe+Sa2g5gkeGfK8QchAQswLQqajgKz8gtjGH2G7TS7q8cHg
Ovlb51rnQgU3xSyRZpYCnmC0Hao4UUFsSaDf2n16XUW9QY/mGGBb247MlC6DvcGk
MjgAe/D8h37zLDq4htmXrPWRBJcv3TgQvkkjwqUSZ/eRhQ++D9kMj7rVNLauCZMM
Lamy18K5lvdSWPSUAKEYA+Qe2/cn0Tv2bso0aO+pyJRDFjtt5atwe+mP1k0D+Nxr
t9AQHav+qRvsowX1/5XAtTw9JmYUH/c5viTzTNafoySSx7QyHqDw/HQ76CbsDDW2
hPJ+JF3oNuIqjFwmvZ+RO5xDcw8jb5tIRisYDd6Nb7/+evSn4L3IZ5emgV7rkvZW
b/hwmZe4QFW8ZRlufEnrT6TelP2VsAxzcSAzmKT3rLVkSkRABK+yhRhfk0aUyO1F
XcAraQz53lKUefFbZSW7a46mHLEXdZS+X5O/ZmaX7oQRog1RBLusxaTbnn4dbhcr
28iFThVOAhJNnkWkYqhoMFcZiFQYl+LvJtwZ5CClez4VoUFH4Ngu/1j8hoWPG0S8
Q71l4mnLzV/nnWftWqK0PapyWv86M7PSxtBhDVpEdwyJVd2PS8o8kpyMFHN5vZ+R
5aDGrhMH4RJfIBjUZQYLoaqQltbjktifhEDEYY4TLeXtlSKyfFI7IMK3gKNEppTL
W0+N/LYaRRRbXl04qb9doB3JNqdrfdsCrXGkXfzdoFgrdpNNsLlVC7cUbcL2eJAy
1T0MYYMR/e+5AnKFopwwlZ5pqUtBl2SuLbzJwXkS3aMpgh9z1V85534WTgDoJr+L
dHX06q43SxNQvIP4S48V+A+Kgg7MJp9K7bs2YdQv5MZuMyABKCweGvhjpvqdp+Xr
sxfoBBnA10VPcjZmDsz6eMX14i0buJ44Fpz02+Vi23iGe1SKt4w0Di0fMhx2FwrY
YhNQu4GzqcHE+cwwdLUXUYCKZmhKY7t+TKyBTgeXpvdu9C9PFg7LYiQ8rKz7lXka
lbvR4KGowW3hBbylJ0Yn04Xwk9JN/80sg5eMrUD7WCZ3GtuXD8ODAg+n4gulbLVO
1MO/9Z2V4008Vchwz7aEZuzgI7WiN7C5t0pczxzXZa27yItp/7pDNRKBTwWw3Gd9
SIjlBLJmX3UXg4TtVtfNWhFxwBErkfVTq7KEvXJ9FHaztj2XoCklm193R0BPYhPY
kBHDtqrVfJ3dRDoaSqglqUGXRco0MDOUfRX/COSrxlMmnk3hhf2Aanx6zHL0ZfbB
aTY5/LrgMkbUVltV0QC8mVGD03zotqGRM0N2yisKfMc0QZZNeMVoWRdJVpJ3OuW+
SSojDeY7Mv52jzMuGQTUkkneCPiwVZ0PnaNnzfMjAs66p7I0NVWMchCmFUWk8qqX
qczYG8xk1hU0an5KbD9Z7c7jixLo0+f1GoGm7roCvVI0A57Dj3TA1SfL+L1c4iwP
ISByPoiUgRmu7tC37r09TLH/L0tOQels7f8JF6pE2IKNt0Gb8Yx7HzS1TeSWVje9
rwLiwpwTERMtA6b6Bppxwew9KaY5WJ9vzDq2JybA9q42LJ7eJ8umrADtaEeaT8cQ
ctz35pUsAP/iyspT+aCuC9CTnRLL66jbUGhBIcmtPGqr8wyw2szr2LWK/gnMfKBf
N3BgXLVf1QZrEbjeo2cL9uplNgPfrUV7A8MtkFQdU2KvXx706nGUdQwUokzpiXzc
Ycwjgom45X1L/OccErXrHkfqaAn5+WwxwRKALsyLevBJPTDAwyG6b5uEYlNZabkF
KHzW806RnRE6bLCCsTqXKt5C7M3RXGEe0Kh9gGZ8jDWCn57GPFuUNzg/BdREW0gc
yxTFoSnDpOd1WBxpxqyCyByL4ul4UvF9Sz/2mcHy3gve3GHOFhAv6pJ6Fd4KruAc
4JyLj1ZUAjWsuwF9cnp0NZAsuYVpI7xMhAEhWAkim83fqps9SNPvpW5QkRBAuNSZ
3wLmNiHdF29h93O7iWEkZ030IVpm+xCxPln88Esrz3/4I1Mex7wv0jKCqpBtlbTD
0w+BUfm4scJcHnTP8/idGwevQU5FU1QN9Suvfz/CD5wxwQf8bIUXs4YCwJCraYAS
qsAnQVgBFrahLbvmMACEmDxbhKUbzuUhUzH3pP4V+wf+Pj3tvPnQpRHz3THEoUCx
nAvinPkP3ywinrB2fzikAw9b2UC6qusr/5EMo9Zy0oDDBKuYclv+tZhm8flCLLgt
/ZSkvw6hLT9nfozPv1jY5Pek7IOvlI2FPTIokOZchflexG1/gpMKyyObd7w9ZbWl
nWCnSWxlkaY6ViHAGPNNKdgE3NkdoNkJk+qH6gWveXj/LDCiuixAc+omgppCzwKE
/wTyMvB0gHPtTlnc8XYCqpd7pnxi4zllHwqj9qQ2iiy5LoMQHVcAMi3bMvWzNRyj
0gzifICUuhDMIsmVKV31Up3KMQS7xOETaZyN3lGhTXFvM8XhjWl1BUczLHLgBkj7
xuROQyX1kvyatLUnWAzwGpooV5bh9xzlndgl/NnHHQhfrnlz1kst98osomNbWZGq
Bcve8lt+M6IEvI2btijCSrb+Jw22FTSM/IflwJ4eN7B1Hdug0ydDQ7KdOClz3tWc
xplMzNCGytG3YoarAm4GN6iqFDvEIUv+X1fqGEGA7jZg7sSPmBkSrco6TU3oS4Ku
n8mr73+FzgQ020nYBPheHB9FgGKNOYNhRE0TFMB/DznCYGeQR/EC/+bGZ9WqDGsm
RmCGJU3u0CV2jaYIRPOKZfqmxSYTZOUJwq9wh3wa85ROfHxMpH7arSMPKBKqMkQT
/1tzOdoesJIyqh+ghsks5YYqW93I6KAP2P2lQyOQNv69NKq3wcQnol794QRx8gjM
sX1zwrqzVZ8wCYoPkbfif1MGwkdZJ0u/LtCIsr88stZYl46Rj8+w0PPC5CVcXMSl
tvezBbB5JhPmxWLZtkkaMCZ+SZFSY9RRhc9cLXxxm+hZWddO/3gHxdmSsJbARli5
SqNyioNpb71ZK9gHAbV1lIPRBPOYHDfFZDejr3lkJT0BoRT771hKFFMWduHXnLkx
SXoxRUvKRYr1LnVgjXxPODSIJK6muEH24pxdCAYtBhOxcGkYe7HEqbWd77LJ+6dX
HgcT0sSOspvkAQoDctE5JZ2j07j0LFEhGFjmtHXplBhWQIZKYVmirokhLfl84xzk
x0tVO8uvznzIZBfIYPCmG8RmN5taYtncfI4Me0E9eeXTE91R7T41KSLlw45ocR4o
QLtg74MicXtFngx4jnTCKcgNKy+zWcQI1DDDnyPQixX443+SldLA9PJovOoI5Y7D
/qVnL6BFp7V/GVKyB2VR9vbU0HFExMfDni1D1AdZbMA=
`pragma protect end_protected
