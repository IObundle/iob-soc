// Data and address widths
`define GPIO_DATA_W 32
`define GPIO_ADDR_W 2
