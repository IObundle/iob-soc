../../../../sut_swreg.vh