//data width
`define DATA_W 32
//address width
`define ADDR_W 32
// number of slaves 
`define N_SLAVES_W $clog2(`N_SLAVES)
