// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jeL2ac2p0rtOEjBCKJ6A+hWj785YCsR0yNErFqTPX3jFb0H40HvCQ0z/j3GJHuIW
aFUb5GmmNSuYhGgzLF7aF8TDaRpmx7tQMLjS8ejF8KX6HcxwJh1XyoBBuAaCdA9d
nxjuD78QX1+ahAfNdl1otrbxbePJFgD2GeLRRDuAhYA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 176752)
dDKW1jp8amNEYRWlkjo9k85jL1hnATI2RFWP9yCnelq8YgQPMVMEJZQMGbVIt/9T
60SAeltZg9d8FAE7hC5KxhhT0u3LCJ3zFpz5IFPK501YKvVUNABYmP77hAGyZh28
UrmU4zwNUFg7VEOq/CH9jmu1Dm2syj3/9h5TIPkz6rx1MbDUEtTcZZ+8XJb56d3a
7wRC46C+qHBQ9zymEFQYgi4/rGV0sYfJp0Ez4NfflUDUjFfP+1AViQzAhf6rpmh4
bF35nfFBBndOeN/r/ja7ijSIO8fDc9xe9OeuleT0BQupME9wDuSkdbUGnpW70eDe
VK9wkVrdBU8TGptgyDP8sv2gOUvdQoumZ21xatfdPCOyN22AXU+72BRWjwRyOMkt
5uuLDBu5XJJUjpOqVLhAY6kMS5K0BoJYXL5jY3IM6F7jTvr86CcjJ2ejU8W97I3H
CQvSg5jN3cT/uWFQnDvAV8CIqpyHBSIl7bVAsPOTxh6rGBXjC6eMbyM16LijGKrU
FusYW/F9zJCRwjShNCg3fI9Dh37XM4HuIMFpVIZ5p9JDQd4G8vQdrAMI7IjaQDhV
3PHruwXNjo9hK29q0FntzAVsLDggqLpdw9PZm1qqDgJHm8ZkbCsaHdUeoLkghmlK
X4xmOVRoi50tmMHdA2hOiwP07H05RaLtaoYRsWGShmU1v36+IPUW2s591S03Al55
YEvJtzUmZPKh00bMx3VcFDgfTN9It0Qkdzxafksz+2+bMKwYsrPYENeGilqR76ht
RVd1Qfh2NuNf859G+GwHrdkRfgXWuaJL0sjGay6sXWvIBLy8tdpXv2CVOzFNKx7s
VUsgUDYWWjRx/XEhwy3M7LtYMWspZTNBg+TMtBUWDHgBAi4V2Oa/kp4HWD1+h1VX
KTHDpU00ehkUY3b457SYVTFknWIkykot8TOGcPV2yi8WUiB95Y8EOGUgxrc0rS/H
9TGVaOXryyyOd3/RGlMoe9UjxI0LdJUFYeofu/mgsmNYsRl93MplhmUz2ZtdwaGf
5ZQuw2xlpKTMoupVTrBVS1l68+v1n5Z7y3I0njLl/ej/FojTPukAP3p19g9iW7oR
KFJ1g5ONumJH0BA/hdqMWOs6oSOnLWJmhv/rIFBm0YblgLKvpThhngUlpt9PbJHA
RRpsXbEIigOdrroudQgl+vfGaQ2xP47BWmuVBY4UafAXinLuBqRITlB0LPIN7vZ1
x9GCf79d1rJw3FsrprUph5r8YGWKe9d28I22DkB0bU6Xre3/Oa5+SUC4QKaI9Fv8
1n7IX4ROTeOt5s8l9G5VRg7/Buwc40CYpjsYly6prWR8EblxVeg2oVRHVdeiDCiJ
SPlLd1u1AFJnuoCJXKX4Ob9htZKzo8V6UWrlfM39sB0BWQiEIXMZTrDRt9HTCn/g
qd7fJVBegWqTr6+RMX9uQ8e8U8isD5Bp3Q/TeOODM5DUC43zjk6LLnYXgKfiREWM
k2Z0XEdJeiAwqjqU3gEZoSG7QggxpVBb7CnWRXxDTj9rLraihSU5Z//+wlaD7SZR
b9QdsJgEI4HmvF/7SlMITJdj/yf7tp7HB38AzWV0ugIab3BAgIwoZiwCgKQeCGM0
UJ0yIRSyzXRRScGvqAgNknqYetYmUJNC7v96t3dnpYjOyklXjyubYbT8Ui36z4J7
wSfD2KrTvPSr90/RqSrcprgEANaPKhPXICZfJFLsbc5L5a5htLNgk6TaFDPbI28s
m/LkLJ8CxEpdUUrQs+vrcCTiI05ehJrOLN/Ro2I5H69uIjFspJO/D95d4OYjCrN6
u8ZYuELkkanlV16WIZnYL6kjInLk8D+4xIzp/2TLu6NV16UOuK8Aw/oBMXp/ljhF
SlE7Xyf/QR1clxhS+JIKkktY243RM7UrexhTT6LlyhUnkAg3uDQYGFW/4LgozyW5
UJA8AO28dCxogMiBlwvMnepXBRr7aso7Hl8RTaL94bfvjDJwbY2YiyR9RvwltqrJ
SnUZeP3DIDwmafH9ZwdgCjGudhHi0WtZmn2UyGceUIznr4A4JMdzxIAbwZ9epCge
iFpQB9hHGjB2gD1Finrk1rdSWFYqWTpgOATvEt31ByD6hKVtmJO6O/FmJvUf1KTB
tfPv5n81nzdHyu4fVP7MXwhoyNlbbZNBcedc9n1lHo+8YZInhSLiDRmxDRsRnEvN
lUXhYC7Xs/BiQGf/Rx1hU/7GGLOtEyCVDx5Hh1NTDjOLbZSNwX3Dq/39z4s1hx/a
LDX+HW0qdNJ8sMTMBQFT9TRBJVBXobEh/DajLJPlo80Mysb2g+5BQmp30MbeJUFx
l0KH6HV+mzRQ1Pb30cOkGwD0F7rI3Nq51PXpWy7EQQhfajqRhI98ygThLf69IDVU
fvRVZngRv922EiRrZwiJkipY7hMkTRS/JVQ+OWU9tv8ji/Pq5Ur2VXbTDXWgw3Hy
6YRPWQeyfZUN6ufGQ/4gz51ginHPZqL5Qz7nrrC6BtVm8tlvG6bXK6lyy935R0hx
OrcBCmtjzjwT/BKlJTOAnj0UR5p+In0iYsc5YlfBBEjQPDx5wDU3ri5fKry2hv3u
ADwdfjjBRXb4NVWRRtfmCpXtpX1rlD3D+qDulVp8gknWh0rP/05xF6Mg8IpTXXuf
LoVH43qFYJGNf2AKM9fl74ti521/teaQJShbIqlQQ5l8G9ePTsGsqPbKQngl4Yrw
ys4BhebqRyNqwy+Bd/W6G7SSWAHkt5Ua+OdzjWem5KTAcfj8Ie1bN0bBcIS+L0c0
85YIs27V2xoixBZMhlkoq/ytM2msarrk8+r+Fq7yRkwY0cOhQK4Nr6tiekgqpzue
mm1SrxLgOIT3LCcfb42mFjFgnpsIzWyrW86UYHs3SFqsPsoa7ERrjim3sPWaqhA5
nLV8cnlPFW86Vu+0LdpgtaE6BisntmQtPdyRhk8ZsSB7kJu8Cs1Axdjn0PaatI5Z
RaXJpaWPbXbQYVpvy7hofMgE4/nlpDyAjU2S+7Eg4GnOeMRmcLdqqT5H563JlM8c
cXC3/KOXCHhKD+MceEl/1QMHO88duTNt73Ju82ZnL4I2/ThxxfpOhMfW80djWMxS
QwKjogROq7tOhmFrvojB7s2fmSA/KB6QiBbqglx85n3xVtnyatf/soety9jiqQbv
y+aHuxVDUhjZZMsClyv1ftyA7/EZhYvjggM9JV7qCcXPYTykPRdoLF7I3+XmC7eZ
fs4MZzaNg8dMVCnXV5PeNzelKIbQnMbsn4Pmxg0fqlclRxkAvqWjlS6SWXUB1P3y
th2d1Q0GW69ibMQ+VDB8S+SFTpCCQI+RFTPp8RaSjyNlt72/YPyb1kDwxkRJ512+
9jjJfU9h7YkxSFPhhq57X8IFt3MgsppzOkSZOLSE77pzQMol0WhxxN5fFoqD2y1N
rqLmzyBRSWk0sJmIN+iIsE2y4jcxzGepwr+Qw1WLLh6lENd8en7P+Ir9ao9XbzV9
wkeCM1dM0pG5t5TwdZBnuU5CWn8wkSKMj1G1aOuWyVkyCoqhV/yBSpGsKDUV4Z36
MEaWo6mJQvWMGx73rO0PKFQjTGik/p3xMrFXACia+KWzDYED99YsfUJQ+/I74hdb
VsvG/HhVjN9vKwiAA8GTSlfdRkCfZMBVZBP1/FAay00B7bzMmBwastj7CdIlqkhS
bdGYFZptLhYv/+FgjKJ9JqYRlGgaPNSM/4F0VK/0nnznYXcgllgHqE1PYlGbXigK
dYxHGsYygbYMcTQwvA+GW3wF4dhFAabdeMY666QhWPFax2r7mw2i8aqufIwSiPgg
6NVU+duOsyMNO2lTLiH43np4Szh3ZA4BwxZM2liX6Piv68aJ6Lt3zcKD8TxRYFsh
vSCHiXbLqOSyagsKs0+FkKXhUTWIugQUCuH/pTQvTQxQ39rJOf9hisoqaHhhALfL
EOq0dBBduoajV8JGtwYFIcy7bAtWJ9Jobx2KVrNXvzQ/pOR+tRCaZZv5bCmacY7j
qt/n6bmmM4eVW8eQTZwLqVtjX7suy1ZL+DqSQexPO0guMKet2+MRn6Md3Gu8wu6Y
fXH2bUE3VA4XZKz830OTkxRym9GQCvSfL17NzNuAmgmkNiiSUGwlg5WqB4JYVYa5
fuzHn+ffJIJf3U3CTFhqqYz7FG275kcqgeyKzltwOiX06dGZk6wn3jsqUYYSh9Zh
P7kN0CamGxMrwNHaLJTKV9VIQu8FeVmi3MOaqG7hBfohDTZixqCyR7GrMgUD90SK
Us3w7P+e+zZH4GXywhis5AbZ1CeoKUungDEVTU8d6T6vTd88HssTEx/zik0xxi2y
Kaw0FPEpEh41zTiOFGrm/DEPu3PbKlR8aWcz8kj4FJCGnl4zq8vO5d/kj67hwDQN
LEOsPKCfD06Jb8tbV6b9vA+d8F6zWJVsy1kbFczclGGS6RLXwp/QDdjqja/1oNBs
E8Ley8i0SpqG/kSOL7/HJnXhVEGLaPHIHKUmIAbfw2U6boZaqkxSTUsUHr4LEUR9
RWFb1wi7AsXhYWFnPnLbcFRQX1XnQ+N+wFxSI6vVyaEfCY1LNnFugYnpVmBfhQu8
TD58bMdNbWI/bISIVhfeyj0TfBSZ4wNjpOpAXZrGJVcM7CYuQIoGJ0OjlkJAnfcT
LRmk9rxeSEdTB4psFYh83zdjRYiFzBgn4Eu2AUNRsh88VJ3kRtkGT5aqClTIQICv
byaeBXUAJl+pi5hvzCEsBLfOC0v5s0ntwW4Fyu25mipdUWfIiXVWlTMGm4CYwAyj
lfDfw8sirQqal4rCpzNLC7eejf9Ha0naEx5WBvjo1gaLOmaC5Mh0J5w2zcPiRK30
R1Xqoo+/XMlMXMzkrRVJ4Oy7JktJ8Nv3ms0PDI05pcAMNSa/y5Zp+stcVI53mM1S
1bx/rHyNnLD1qgI+WRMMF/GQBWGGOGSLTrucdKNeQ/iToVlx1ydn2mRCjRG9qAjJ
HnjQmn1n5Hm7vOI20qtu9GYBCsHH6EjkX0gu28u55lRp/OTOVF6zKgcWkJ9yLYcA
9oFGlK1+q8cII8azofBTavFk6yo25MdYLkqCUikjiJEla8HnGJLlfKuFjDcY3Mdo
6GoDO7mjXgJBm35i2KBamrrli+gs7h+mKSiZ1taawMeEPQ2GNHMHQfXYJd5tl9RV
6CGnYeHqLsZu48DlECAsUg100/p2Vw7E38T7uc7yGz897I6lhkz7Adw07k+aegsT
j/zj/ge98Dusc/CnvYYdkKlyGSeTGrApGOJDQtAO1B7ovE+mhKE83ECC6nkXUd/2
HK9oVwkKTI+PS5K/hslnNd9YVqDuQ7FIYlYNHHZ0d+DEycvDrvBF1oaL2w/NISCI
onIuJ2mmt440y7xDVONaTyqRPQop6FaJM/iPpQ/KSUNU9KbkSEu3/CauoLMUYlbg
nCnKxBKzqs2+ityAD8pt3QN5YxE6w2tnfPb+EnoPSbHO3Zh2mrD7ykVa+eyTx4Yg
w2P8VMNd+hfC8sDAB2Vi5P5emc4V6jk64PcFxmc+1jQYeWNrosDnNDGFn9d3tpik
87NjZzN+X6nsPHINFU7TgF5YgAPTlc+4ADugWZobMeRokQUveuMCTa5g8Cwj8gFk
CfGkOfdBQUIDy/Wq9sbwELDoFx43cQ1Tk5uIqIQeUcMCA/SKn/hrcadD6rF9bh6R
LAkzzOSkkVaHmKHJ9Qgzcnh7kPA+/2pplyinkTpx4R4d23ZKr5lc6POwIIBcSViO
rw/0ofJaKUB1FmTXSBcJwLTew6JmyKCW6V46DyL/bDpcI5wA+Bw5aM8OlpCM34hP
DlWYJnc0x/Ww+fQZtl2M2WcYsU/I6nH3d3JDQEO9nmk7EWVWVLmZjjDsijxvGVTd
5xiPpXoR+RHikIsMcWINZTkCRjlsODy1S1S77YSoWDrjeoi0r+cn7VSqwWx+dzYN
VV7VPskO6ZI7LIDCYdBir+eKQ/MGoh6Gji9mVlR5hmfhJxZwoKcKb46JxmKUSdK+
NM6Jsf601Bu14kvYHaZ7ArkGHyI3WAwBTDodJMtISCLdbkPFWql2cM5FYPtCH1DP
dKK708MRqCT1hjudQiDPk4zO1IcT0IlYJF7DU6LIHfhL0msZRDvK4Ocf07pugIRU
J5RIhh3EgdGpOupQ8TdkGT8rnrtMDSjdK25j/EAkfY24Gzp5tQk3lCkh3Din0B3D
miVkeO2miiqeKd+FQ9l7DI6MFTeHp+aBVr5LP5dc+aNbqZjcTzq5AajvpEvql86w
5XYjge+hWwysovJQiE4aalpHFjRel34AXuOml/Wzt3q8MFA7YAHxUP2Rr1bsa1UQ
cG+W1olPeX7SKDxG8qEtRt45UgwYtq5hAavR2AJS5ZUXXpT3r4hpWMikRWT732YC
zxex2NVxXxzvJp5ROBqXFyKx6f7b53v3HkL5dxondt+OXHBsH8kpV3X9uLyg/2rD
aq4uiz9zuuyCfO+vX0g68ufFtr2B4NZf7tU2qtqs+mpDE694wnepNiaNBNfi2FGN
qjomEAJ5q+MzBzFNqGjUuK/kudQi7QDuecgWMJj7SxRjfetgxPlQs9bJ6MZFhiD7
YttFrC63vnJZOnFDOI60rLiSBmnePfNuDYIWEEvbTcBzcVR/auImBtv7nz1eqjJM
UifmxEMUedJEzVwUlgCV1ufQrMz2p1f3V4AahDXU2Jz2KFVs46b39X4HyvyEZe9Y
gC3aPZR+VVw1wYIViC97zESJgMB2I5xIQlwdrBsOIFoz6H6epFfAE/mVudxwDONT
Fe7FOgkBQIaVicry7llQt3t5XghrkOXXMo9di3pqmevdFC3cGba+cdT5BXhofsZi
7kB1jCyaR/SvuRieansW56S+SazmbiavuBXVB2ixe4LVDUvyAMGED3ZPZUcLIceG
qntjcgdFJSyhiZs3ocLfYgp1gsWAI0Topivc4s9492dDs+t+k4csryMR3+J/eSDL
t/OOa86oeWOrCl6QXZoJCEEjewE0obk9seYZk+I8DdXGXeaseWVfq18MqjmjvqmM
QBGW8TH3JLT4Bb0EAR2BHhoCcnJFp0orJJR8tcUKzzlSpOLNvkC2xolbcKzBy2IB
OlCGjR9AtXtgN0ZzTHK/V9DHs/g9eojCa4D83WzHh1uyo8oLZMJWnALsPf0a3tCR
vBHc2KZlz2q0tMQ2bychb8l1xsM+CuVkbR4sTkNRs7u1dmDZaoRKsef8wjUj+pE9
5dxNYJ2LLCNDTngYyoFPpClTujVS4afrSBsMbi4ixXqncEZATGTC+iY1ITsil0Ei
D4Gd4yA+18afL3TLTSnK6tMBzF2hvsmkB6TI/qvSMtz2sOegZILerVAn+CYw5l2m
o3dBbr+HwP+HnO1PaUvB5bLaUI+eB0Ccy1pmwXchtwJkUn+3ZTilH/xN8UhMyG88
R46mbVAtJXqMjFr6yDKN9MzXPhRvEltkDqz+M8OyvKEdYIngjuCgBQZbht/9oWEx
TcFhvnf365BZJIgCJgeCttA3Hcq4mi217M7hPiSIlXYskfIaGOuWX85efHFiNR+m
5ZSAafZh9dy25OV32weQxE7rRJzUvCWGQiELaJAEs727mYVKQr/0v2UV6ZUW+5ZD
mzMsfdrX4nXX61w9qQhgQ4ohWeCpuLXrnZt5BDTq61KlCVSvn3J3xwv82Clsjorv
35du5ssINBf/ajg89euJ1tfJNNHVbwU2vlED+dACo6Di2WxdQfbXIWpecALPlb+z
Eq0bgOEYyCA7srk2+yBj+Bt7GHa0eyoMFaozpqUkTjAlsvDMQHVQ4nvHMBEUBXg/
oZBLQCcWGDlpA6gnC7wtTybBz10cwCF3nGKkc2gIYHqLeN6HBYrE7CFgnK2srBpy
J6ztBSJNABw5kkJ/ouY4I9/VpAxX2OD/u6qeb29D/cxcF2Xz9UAUr+dhw0Nncq2N
k6jRROTUrr1VuSH+hfUDrB4drPKBOWSdKUD3c3UCYIBsFJbnJSh9YhP5kz7KTYDN
rN5sIy0E8I20Mhz3sjW19AerVQG9PyeoJAiBeOylmLREGJO3Yod+nT4uS/da77GG
LXda7RKQD15rgVYUF+ubzRaf5oa0p13y2fshdPeTdk8VU+Ey2bprVoS6vMKt0JNt
l8vME+JOgTURwuD2EfDB1P7WIgNBNxStvnyHdQ6apYhAV/pKOSl4G/8uURHUlX1y
XoRrT0NpJShLof5u0LfEf+RpzsVNMB1EcRf0gRHU3xGvP6kVMFscFJK2SoIunrCw
nr7BmIxA6x3akXxBce1fXp5+iB2MKtJyrg7rPBCM7rbq3jXeUz4CFi2tqxhRBTEG
nm3JxtCS1iQiHmVKh0FebiirpIqeiqua6D5ADqu1toAjJT6Y8aEV/4mA6iFtdvMw
oFtOT7SFeRTPdIYWXkyzt7tfAJ++DOahUpnNLox9gEsHbWj/t50+LGpCuRyt3Wu+
78aSmiT7seQFqKxVSHtYhfZ70G+9nEnzsah5OM9xHiSnITIHEyBvp1VRr8rwE5mY
2L92XJBD1YMeO6xtKhDcI1uv1urnCX16LlRMAiko3WUZvvhPZfWRBu2XbGESFMiH
gwY9jrEYYtaFnrqzobg8eMyHC8MlfiSduNPdTerif3xbA8hVugR743zPD64+fmqw
M0D+fdl+817NMCqvFXmH0fCOh/WFcyMIh7sRk3zenVfdzpYv5L6bRhrLv7Kuk2W0
PezVIZUpbyfdQKFVOTxOqdQAP7DzxtgC4W5aqyki41QnJe8UzJgHyrzqARRaTB9v
67G2JPq28vQ9ZynSyhBJxcUejJfW+DVgcL2eHKZGIte3OZloi+bb29pESwpYl/S+
/hcMGW6Pj6hZ6cJY5eNy7ylX4hOSoyC3qcSlS/633wAAESwsssdkoMMfuqBpci82
+uGZa1/eOWTjPXyYcBi1vmnuUoEWNBmGf55EZG2p0qEeiJN9R9mh/asNDxEqOHGb
LL22BjV0vqkfMyoKKG5QCgGY8riniLJlx5tK4GuKKHAX3qVPbDG6AeZcGJuYHuwI
ZNOwYkhuLFXZ1uP/O4v0xppKw2gvoG3Die9eCHbu1WScE1UF86amYysBW98vvhn6
oms7RNnUmYZkyXjj7XSZq6nthqWR0+4anP36MWxrEddC+fyFwATlWkY60HcNpQQN
CxBaqeqWunOyWOONfZP4aN9EnZ+mE1A1wyWRE0Md0F9wg7JUWPLZTHJ89yg95lY1
ibouyXrKwC4vGke4VYxcV53Ckx4NoV5yoOXjKx5NbCahAH49Bw7wUK+vutli8Uf9
IxSolP4BF9FNT355LRoNuouuZvUfLaG+93hUHQMKX9JPuIkrONYoTth+Z+DkXf3j
9TkZNI3OLqzKUR7OOjIC3vdhM3CZIYLsGqL1VvQkE5uPn3vocpkP6BbhZxyhUSn/
rgkiJ8z8+fQeRdg51tRV2m0FcDLb1GFkjh+Uohsey9AE4rr3pThpDN6ADT+1QVPP
A4IEjmoJ9ZLvBl2BWelzCvUxYCHiNLEq41dDWeWI1kE9ePtsXO8W++RrNTrFT4gD
TJj1H/34MYd78iVXB9LFK93hCtToE21uIXtUiKrQ7vACE4KWCM4ZUjEnCmsNk+d/
2klW+8hSl2FFG3nC9p4WuVfrJAgQbcTKuEPJ4/dKRN7XFHWKMlONyA4A8P+yrZp2
DS6wAiZW+lQC90gd4Lv5qXCjgsyeZFFK3E/r1ypDqIZO9+LRoF7Y/3hW5c9OaI+t
VFlx7+/9nz8qto+WvmQieO6eoHNEVkPZSm/DTfdng2bSdcb7Tfinu/aoShIdYHqw
/dzEHEGwXAgnZFF9wil+MixP5K3ZXN0oNOCu/QcEpoXYJqhWcekqzdj2bngeBV44
RPP0Rzs1oSAdO0cEzQoIOEkXSZoD1iNgKaSGcN6kD9lgdi4pZ0HWkDsqIQFB97Se
R4kaPjAU+Zop+Ql0wweHOngh9NXnBxmEwR5JYmrIl5qUhR4Sb5TsD5mJgrYa5y+Y
m3HpZrNtQpcJwctIdZpUoJ+bRueEMH6tWBfl+XjsxPrXrjHUwVcwQZLy35476y3f
ADqlUSdLbnSHERTOHyt7KZirCnNuS15Y0tcvxWHeU1vq7Dv5xSzjRdhCriB1cVtl
/5IceBU50bREGDSLusmLOeLWyuxdkj8VacHP2mkNKi7WmwFHtSI+hbGsyBb8PE15
ikZXZydwMdIJ4y2M9jmaENmS6/h+vnCQN9Sm3whcU0o2TRK5GkE/E325HuLGHgtr
k6SwX2W5ya7+kapmpP4huFC2XasB4IsWhrg3QsVzv7KHJ0+7SlFd4pj2w7ta8Wyy
pVj6QxiKBrG9mgqAL6cndKSCl5IrEeRfo2EMY5JOpQEQXqQWycwU8NeR4Vc6eRHw
20e/9LQUsTdg57TzF0psrdCk8L0S0I4fecdhmKkIeWdcJOIDpK2+C+y3luC4nIAn
mJr42+C73SDDYBiHHQodJGgioErFZfbeMoNGI/HuVC2YPIUQpqGWe5KwnYault1K
P3NuFcqcpW+D1aAipYGHsWODDf+A5D2Nb4FFGULeeeRB6rTm6ulv88tTbvHWt1rj
n3stbbth2yBt9z6Xa6UhPKsfdaHDBBnaS5dxE/CBvvhE5+uKiJlIeNDsCJywTuc/
FXEMsniNva6DZVK+bTZUYbP5Mr2pPQsRRQ4ClXEx7L0ImO5vSrxDd/dxd1xlKBwh
HjgInib/GLnHTWkdHKbPFFJqFXwD78xWzusI77raG+LTt+CnKhXQzkrDPTOh9/XI
+jz2YWmn/kOdQcOur3Eq0zniesBuijqMu0EqBIItv1MUUnMYW6MGKL83vIaPHrOX
HW2FkOppP98wkbfL7+GW6ayPkC5Jx5s/cP3STQV/u1MYINSlJ2rqmrTZtVGBD8t5
lrjgNNWfxa7wPlDKZG95gBNGvi5fetuxL6JlwUMtnbGkHX17zWWmP2Xlb5nL3Mvr
49N3Caj/IQoP3Hh1NG+Ya6nWP0sI8CE9PPAyhkkAnBCf6Da+bPBiz870gDwF5gqG
hrPhgTg/+hZY0D46jf4rngGoAi53gR8ENmO4CCUwp7Bjuzi1rmStEbwNCnNoCm4d
yJBSK4YthtltYWCeUl7mLXaZLwNYSzCWxgLDAAc/VmEfpKMBntE6oj9aY1FKQq41
mIApggipGhUlqCCnTTaHnD6g3n0Dldnl4j/5CqVF4TqjdsYmLFDCjY3YVHE0uZbx
5hWJ4lKqa8UqBiNvgUK7BKTGgvn5dXyNlQZRnYezEgoOUaVgguDxvNKz2t2mYCeP
hNNupcXLr78n7jdQTvzwn7Vj2cFqHqdoslKHM+zNcg1iy54u+HtgiuCcl7UcuOAj
FAhcKvkVMtWup+T4K7epVKBlmZIefbb+p4kVhLn+O97ZS/i4sErNzDBlXxkIFatb
5yxD2seV+308JxtOJq2QRmW1h5cydAXswLJM+/XjOha3olPd0fIctgQ9bdgBFkJV
RRPqaUc7HL8X/PME/HSS2Mjncl5LdUeuHjzPmRMIAdJDfCKNeCwhdBptyPRnHew/
8xZ41LHGMipz+Eiwjay3JrkBxnq4C7MSvhIETCWZ0ryw4+87MDpv81ZlIzhj0OBK
EKohbupEkJTku2izE6slesGTRftV+IAHJpc5k0Qt9wFGiBwSMFfmr94ERDnV8FAj
hvQl7RBdxhek1+TTW9vZNvge3wu8cwTXUAnezklxP2ndH7SNr/lRrU1JATHYDFFs
b5sUMszWf8eXL9inmzGOUtmzNVaH382Ml8FWjtQaCs5CumYVZqsVNWbxAHwrjx4z
MnEQPR7crKjTC6c26Hr/G3+coAd8H3Zwn27vZ31nI5zIREkM3hqnuB57NO60+/U6
+sk7gjjop5qbSMbKyanDEK+f5tRoBwVXTibnuUQd0cgB68WN0dUWIstdWw4gx2QQ
M6hIan9JIcS5jcoSj4kPaUFTpUDyEsoGNNP5t/GmdaAUUYLmIO0hTTlZ31Ib9CbJ
BLR1eDc9UQZibwsEzER3SirHFoKWr6s2TGMe0BWNPXcAE+nPbfINL6zSlMBLrod0
6L6r50hsoL0IIlqxibY5QsSj2VvPYHW5GzLHHZNGTh9fr0eC5L/vMxNn2+xJYeZR
M9jSm1aEmIc7qVOF415cipuNSaYqTD1h00uVa9rq+VpmU5grTmYr2sRNrUAx1dRM
zBaLmtan7BCn/XyDcn4pcmQqP0zZ1UtJN67/2CXkpjEbjSNfmApwdmqeO5sjXW6v
cZsRzkE52M2B2/BFqn25yuYU++81DmKBCpNq3rNfgiQTaCbh0gAjNrcxwKRkBhvX
06+ZOzakHm5NQuSkO2Bnea3fTaFuDYLx9i+H+U11+yPp7kyFvubnGeDTefkdAQ7P
ljybgQnAyAL0sXLRhRaKPR7styNH4zH4INA1wt4uSFLLQOnNQgC8y27FF72lxx6p
x5vMRoSyXyggsFV2qkRMjWsX8ocHqZZ35/8tZksY/fd/KXwMOb+BCwkozrunK3qB
PkOc+qkjEPiAV3xwyzAmf8whQoO2pPnbVyR/HJy6Wm6uZzonIlwjYChZJkYAlvUB
rsBhFNCwcsXk47OXGnfFCFPVgXkbv4icX/hYcjXOTa8OJu4Nl8UmZQWx471QqAjw
jzkxX1tIbq9nkr6ygTbKXU6tU81hvZ8qjrqh1gRP1XMAUNJ2z/ZkqkT3um0BtdMP
8TEErqEcePBGJr2E/DJkvTmGiaxyrqJrVys2syaC3LL9dxrv9iiYMCONBE7AHXV0
lwY6k6RJbYwXyaVkWhyevlOtBNMcsyWskKMaAg+PHuaWis81sKvAWFjc5RKIK+hE
fCR+G/UPodIgS3YsmNQSFwJ9uBpMqf/qRszpOLFofC7Luf/z19sA83hGuLBs8GpD
0PRCTVMGX0heUxhV0E8wbrEFKuWKGM8stLiLgxKeN7hObl9/LN1JEIZ220eu6R89
hXu3Pmfea7gMMnYnxZOLHyg9T3pN+wxozgynULkOwh2yCTLlmmkN18Iu+faRUBTa
vCkUCnb+VRkJm42e2hVM/RlE/nCF8G0zOG7/k9wBpaijclX4Gms7VSjpr7GllADo
njvyUGXdVhVcSyf1OQUxjkIPAVBH/2VacBUHkffZRb/UdXFkTewYiO/4bBKxyD3B
l/GeVW611pyifqXV6rTaueclVc2Jb6lucySZzPIAI5MXzJfsjxY8ittO4mxiQPwa
eYOVQ/0z/3T4FWWCkaEZSTC/2bvRR6upcJHWyY+B1Bx3JpleRSQdbW4XqgbhfZlf
ZjH9MfU9Bp7IDpImcR23Wd3o22DJNM06etRipMpYny4NAWomvt7deKauMTAEIAnM
KLbAk3ahMn5xfGEDwHOCWeXQeH3zckO6kEoVzPSbLqS1NfDbiMA6uEICXXzlv5no
ta4NWAEpGL9Tmq7T9tDWKI+IKsgXwlYKbo/ykJnOpBo4FRunTHE4gCoJARR0Pwut
bjUQOAgY8PctS9XMBEKj4LHNQyby8OWFfJ3dllVgEKNxnz3kSYFj5q2Wnurn6QgG
emlkbFj0IzTXIejOUSUMl/5oesbYefTyed1GYrwdbdVqr6BEEdXVDLaIG/eJSGxJ
i2KvOCbffnwAlxFeSAzuv2uZ3BeK+FOPq2VzzoE+eC2BVUPuh51RLDk9xc8ANMMa
EgrGJjXRsJ7EQrnx0Xa3pVuG0HWwXb04Xcg+RFeezG3QxOnMNImaJOIjXBnOmeWa
NE9MAGWX201m4TESHh9aLYsyN/li0IEnaIZIwW9fa7ca1T4kPEhq0nb6pAvimnc4
Y8sz6joxk9ik7uJq5YqVYaFVWQw/84nxj/vvdJqCpOm1U9KFBc+m30d7lu9T2wFA
Z1TYPWyddnTD2TUA3tmKHB+/6hswerh+Fb1THuikXffpB/a27PRFsQfSxa8Ntt3n
5KGEQvj68tNyca7kJHL2mrmY18Bt5X519B5OvIK4Fi7AuJD1JKyqu/dLgeK1D5z8
qkCl1QupeoUeLU7zqUKVebNKIlzZo0OhVm9mVqFjb76TBREDxr4nQgDZsd1QhYRT
CFOCVr368rnHe4MsvmZIe9MCNUUzv9sgYf4s1LPDyShzrNIG+T7dv6j4mvp4d7ti
Vsek9OoyinNUG+H7uSDAMiLx/DeYQ9PzJCV9I62D1bkwyrYB4WwnJyb4T3FWuOtq
rCcpi9F0mspJq3xxgDjTuvL1V9NNHt5vXvS3IXwiu29rKy5ebOuz1isqpt8ddg6e
vBsUXvxU/cp/vj4Yd4IfwzIMRK3B7s/tZqCG07Dwcdyeu07FjdS2e4WWC8aDLcSV
4pQZicLaXyOgv9f/wdGgYN3Na26O8oV8kjSQMZCyDB1fkD+OuIeBE53nP7uLieRB
63rvdYOpEeYD+0cnA4HJMWCBkMWuZkwBvbjZcBLgqQAqd5nQp8m3EeaR0saYi8Jp
Fa8xq3AYbL4QMFZ34FCtTHUbcF5bZXYWNS4kgilJZXw2FwFvfnGcQZ8dKt0mdpHr
L1eN4ereTLRIUERzafIe303fe2BM6HeFdjaxv5urgxV1jvG11AmpCY5KH2VTRl21
3upqLgZuqNBATBfBYDyZWBuRSxZWdkuXUULOidQXorzOo+0qPuzsbYkVXoPf+HD+
MacF23FJIkRy+o+GCCm3KLFEcY8tdLR9fZwaBOBtLKwXJssE5/dQpHA5x673fjjt
y068eRjFwiufR5biOXW/pAGFZjZ9OchoxTvzuMtemZUbJW7roV8mgv0sL9rWi2jn
OKmPwBTI6+jN3w4gQGgPIX/0g4T59MarbaVFC+/tMwTHA7tMKW4O0ssEV2flKF8N
n6v4CnSuDQz9d5lMx+u1PrRIoNDDmb1XwG61x2B7MUIFvr1VWVzBvCEAykkuzFOv
fDRA0TJ5NiLhbKGgAe3bXr/8vwkXvO0Q+I3gq57y9JlYd1qVed8zTJ4LHYVNytGe
Ji+guoryRdnNXlqgY4foKQCIDHPuliA3EEnCZnkyjkUPdxPe2h148PEhaqDDrWIB
VAxaTPsZi69yzLJbD+RBPPc8eTd5fIQlJn10XJupYQvIHM/SHav8pMPkShV76wmt
VTmz5fAQ4NqC2xY/Mv5qHtImf9ORtULV0USp/mFin53yPJUPsHkv/5Cv+RDSLPtN
G3vvqjs/0rgCDGHMqMwUeyA9YRMQeiKAxXaNvKbF3KuG4m6x/cuTPkaGFWI3QQf0
hhug+NjLvQnszluUAERPw1f93554GAlUSH0/9PQORxHHWqhjVqGQaD79qAkU2atT
rrjlAXMsP+G4AAG37xH2FmDyOQHSGrZ8oHN/gTp1P2fOlrdE2sRbbxlFmz9L87iQ
M4QcGPzvG/QIFURbNJCTednQlfV9XEJlL8zlkGgcxpxY81MZrXWIEGlzzjLuVja6
CKk4nPo/xA+jlhF0+AKQLDQlrl5ALtNZuAZgGHrecf89D3kQ3TsRT6fQyw0WhNuv
ovXsR0kIz5x8FzFCtPxLyo4i9KGcl6Kqaen5Q95AP4CVwCc9ab8YR08jhhLZ/5it
eskPNCkh3r54U7fISgqPQX4glI0eMrQlCVaV7bhGS1USBchhmYRgXYopDUCeB3r4
BV9X/glOIwJQJJGwKz17xiHY0kcDKwwyg9t34jFjfz9P6ftJk2jc3PZKlzN0KJEs
+3j5pR3fd2hKW8py8O65L8CZRYjVy0qifdv7ISIK+3TXpP/Fm+nwfy/O8EV15ZKc
WbnCVDQ54pV1RSX1Y+QGlnRv42TBUgIsCZ3aVqetGsxMg8bPgipc4xU3FUzGY+lG
A+DOW9Lqu3qMkbD2PPiT4oWkJCUkS1o4+gwqPgFX7qgS2vTHRcNUZxlKipB6Wsxx
PuKavTZurToWY+zN9ocGjtBhX2TBzVWQlIimONvPbT5wmntMSP7GTsUzJNNi+eSz
pOq4Vjort+X7ERlu7kf2TjTuS78h1EYPlBimUuvbPcrgnmivXFG+VSL/syNKWuN1
ees/hNfMsPZI9oHOH0g9AObQ1wwYjZCzHU/w8ITcmJ/rLR2nkoykQd9ZDMWtOGYL
xi4F6S+216vNpKtgOKr6YQNOCofLs4wSbdDbcMBOt38urfZCISU4NYu92EgUBzeB
7nAn0UUtgrjluKk3i8iH+L0H1xW9B8ifUZzRwxfkt9txw2hEMm16VB+07xCUsbdb
UCyEKbZZz82lqZPXE6stQgwBKbVRnFFMApkCmJMcGrqLEkvTQtjafwjCPDWUaLeS
vBDd0ouISoh4K9niGd0ImcdZZJJxU5jY1+WGAyyYefCm0QcbMb4G5enX3DuahcwZ
NL39jR+RcZqUvFJffTQLQ9c05aufl4dOZ5nyLTVaCpHudGFzZSgugXPZjpPLSuyU
ZZ833tU9AVS8aC+7Q5U58JSeXu4+pQ+m5VEAcQt5lIFLrcNpyL6yQG5lGotxOBgq
fevE6UHXL5chjMnEJTYiZEaevblQx1whWM6h6JrgGzHXtIDUj0R39iln5Aub/Rie
pUAyLUxbuHymvI63WdqCa1gX+07JLS2pUbMJCA3H29RGvcUXyNruuLMiDzCgEk6N
1vtRVJo2tOMAIS/X/XIBFcgoHMrM9gNqCNkml2ag/ItV/tNo1kH3FWnpBPcVPCJC
FURC0w4DQIE+ODKddntvqpsdauTxoRwOpWSj1+PyaroWSvTVmX81zemOe81xrIPA
TjEIB5ndOYZmJE+AfeuqdnWbSVRu5TpDUXkANi0PYqG5HontETo+CSt4BjAju0MN
/KXqlnbNB4spEtPhlAx++EGdZJ+3ndb0nWhGfMyuzrMfmfefc0OEhlcNHe2kfcLD
117VNiSddF1OYdo0R2TogEt21zoyz/LVP1cQluYkFXNnEDOIf4UvPItVgMVdh3Tj
YO0vXxEVDNeDdji7nz1wQAhRY6GbhjZPC0V48t7aTA3NYCtJlvTXHs1ynecbZrZ1
lnpNWstIV8Vj2/gb/qcdL9aw7BXMmIQiwsEvsoDTPPocZ6xIAstFzD9qqqWW0Kh3
wUlaGT9nh6KM6K57hbDR81Ces1WSBsyP33ELUWwhG9vLdspHWmvMHChN+eXkbsHY
xSYoXSDSW2L6mcXBLjfYqlWphei6E9KdLdzc6KH1ZpTWHAw2fZZIXNwmrdPlJnsw
f+waOHqXvY5pBAlKCeU7NFJgS7Kxf+D9ZtaPAeODMLkKGYr3tm4F7Jkwz7jgqsx6
fqWuvJAnEitNS/4i8IcgLCaJmODM5T7Os9EkHp9SklclEJwEcrrEEYiDmkdIaG0M
+Ci9B/GD1ydEFehrp+dui5dvb3MwbMGW2Z2UqCXXvgUthMDL1Fg25OrPc39+mNEW
67ZEWrAN2Ds9Ogy0oeP8QaO90Q/rOaDXxV6PTR8vm1eFf2y3I7SMC/WM5J3kav1+
Faw4ank8MBDUPVIOnlgXvAx1YUfYQziVN7pcNEbOnrO1WExNSOXrPpxr86wWjAN9
kUvJoFKay7sgp8kD3c38wxJkJ5ELlb4d1mJ+yssI69R7CMoeyomltwsgkJnjm6wN
VtXYB2/9W+zrOaFrXb71k39A0xep0mBoxfuM+CSyLoJQR3ImxKN0NYJz/JaiEh1b
1Fs9G8bh5FPB0VD7lgA+D3P0bqh8m1k83q/2Xw5Ve4B/CL2I6xYa2KiFl8he3SHW
17jjjY6D6WgPHKYyC7jGqVYdTBuxD2HmUxh9IsJDll9HuaAmycrshfMSTmmN1h5g
5t9hFh4jO/CTkjgrmOs9g9p/16aUV2UxCCq8kxxwr4UYW933dZt5XN3F1W63xXrF
dHKKnthkZselBs5Vhym1cH9PQSTPYSGdsdSfb5EkAh1oQGX80LAQh0+QH+EPYcri
6PjvaUYl0JdlgR8fYpzqu+czPcvLcbAE2Cb5tpN6a6iBmfIQoUutBGAmo2tKPbQ4
wAqW0TJ8WwHhl3IFAw0MRFaA1wrsqBdQcH7D5to0oJuJWOUK5RYeyNBBi7/c7WGV
J3z1Q5UKQgjBEVJEj6Gs0lBXIJcI4JqaTtfzJqoqGqKNSvmlCH8EnB8nb22Vej3B
ggnojRowWYk4h8aks3s9eOlCv1nOnI1NDcDrI5eQHRDTpxp68sWWC0lpEYfWGe2O
BTM5Yjk9/ieHNIPYauk7XwNXyHQgR6h+7twJEZwVjHZerkO0elZlUUkh/Pang35y
hCIobwUmeURf0WtqLGnSZqGhBg+uaAxrn3SZLgI74rcgr2+RmOMwRftI5uLWc/k3
zWgIIHEV0KbfYA2mbfbftynkfEclFhAayPwIPyTdomIMoYUeuS5Jrxy7XCypYcWe
EQm+aAOa0LLL6xQ4dReix0SO7jp2b9S3YysPHRvhkTLkMjPDlK7RO+LRaCflkcvC
NixStORxrE7nzfRYPL6dc0cifF2Mv5j3uTdNTUJZ5Z1wd+UEZLV6crgJ4SbXLmHF
UdaX4xSAov+UX4tPGTjXJ54dPjzrjH+tzrNNDoh/Hl7C8zCo/c4vZj0dRZ07pKig
05lGYDqVrHaUQR2U0vw63Dltz0G46RCB4/ll1lrVnQvIMygzRGuyXMKWdJHMlNix
6YfTBxJFYDVUrO9/EaqPoF74592p4umAh1r1Mah9qqCpA01GaWXYUKB8pJNpNM6l
lmgFN/dmzi7rmselS1zJ+Ovrbgai6CFgfbibMrzpwKjHIm3fGVNj6v833S87TaIk
sB+VzPJPGxRbDcFnC0HF9njTT4FLOSvZ/8ExXdsI/hZxLtHmnBq/Z0trja/PQO/J
/gdDlE0YY2cperbShkRLPqlTYvr70ojGwAmqfvu7EW9TqNG2HOmKDwp0vhp2563H
PoRlz6DdGqT4vF3fyu85ZeAyuIJArtskuoLcQ04gkFfHgYZ89b2OpDtFfjU6PMy4
i7dgttWMincfgbQst6Gf9WRYiOwCVHAZ2owbAVpuXd2Ga5PTMnAiLT0Hvji2k3ib
IhPi6fC6uDifTmxofaZa2EqbucFWvvn/QA3U6dQ/9aq7sCSXt54QklnPK7bqJ0wh
gTsB9bSQQNYpxk4aBv/DZzuFlBhPgqHlvEMZ+WGM4/YqN6U+D28wHCbZbjrmaKFq
CoTe2xqezK9HdjBvnQ6MHdomtLFaMQbJRZSwXYCpVG5DOB242Nh83LBxPCT4IxoU
J6o/KbSzTYbvNzeO8p4YKk8ANzM9qzJkvT0ePdxH2wYxwOze7y142ZI/dGs2gTi1
dHwQJsNOQtLIMdsCt/j4GSisZfk6MmrAJdEovGp0iER8k1ziov0Zp12pXJ7q0YSs
cJxqMecT7DIm7oBVM1DMqEYPrbgZokFgVixeuN+uOW9N2UBV8+4dlxZmPcW9Du7c
g5dGg2m+CSfOfx7MhqYyMddd+XyPrc1cDvGp15ErmlNKgHs11LcNtpKARx/5asv1
cXtFxS5kQIxa3syIpy3/0C25xYt5N0WFT2jLHri7OHq77N5RkFcmc/yr2UKdlY6l
pOL2p1BGmxZSEPz6UPl4bHKg9vr1oIqFMxaOCMlP/AuQhrkSCFs/0qqJRjnBu3az
1HtKgFd/Qkms67TZy+ktwZYev1lvcWmMZGel/JhMRBLekP3QO/QI31MKgzZ7FJST
YUlop7DTcW6j7xPqDIoJcvKMT61xujCLJ04KTiDWDF5eUp4JihSqNotSacgsuUqa
xuXGYX+R5bu1Qy5p3TVi0VBqDi4PTMVCThxv6/zCP1Hs+Vowc7IZdSw9AxdO5yF7
NOmLA42dCsiBvpyh1JHgVE+u8fSaQyxZVW25PcJsBnpRU0qbqLMkfWj3Sdm68U+R
qYsh+i0jXeUCgUCE6G+sB0cJfFBY2+F/meVqHZQNmwhazP6yJezSXxIrWrcs+jyS
88UuK68DdXaxO0mU1AbFHHIl/95vbeFyzKFUwIQRQnKeEq3HSo7DZqBew2MI/BZ/
UBFSnMBZthC+LIGWsK3Rtk7sEBeCECAwgXKbf4GsOGoYyWJxF0+bzrqZcNRCGROz
WbehoetvJ0eOgiVFrtQGLtPR3BZcc0x4f9a2iRgGH1k1Mgmn1vQvbs8nK2xHL1Ou
DQpX2WxnJH9H6m8Ts62G3r/q9AcED71V3kLv+eBrY419mFLwHseUpzj/el1fbMx8
3jYuu2JTkhjSTOOkDs1YIdpo8xD8vZ3HTt02emFKW1LZjjMD0lqQ761y+zB9I/9C
5+VZBC5gJw5o6MFEEO4u0HHeuHOPWmYEhjwRUPRCaE/SxIVIonf1GaSVI1y6iJyL
zCBIk2jYV2Ydew5gKFhWMIQ3QYcQoi42SmdYs1zZTa9P1aHzBBsGdKDJqeZU0XXH
tWIAzKtv+1tf1CFifEw5skvsUapqtO+bPznyoxOlwLkyBk8PfByGKoHy75Lhay4D
6ts/JIftmzV5R0OpJNMpuptvE3wX8Dgpe6LNO4Vu+bDGKUBaRxPT+lR0knK3MUi+
UD9pSxN6PjuC9v3wvhKbH9JIN3Mq3jQpXu3codv5hjuIWJpWRLzXeT+TXgGAvc5v
bcqstmWtf/BEeWKyz6osqDMaQz4HhLkPeXlXzEo/s9GQ0ToSQzhcw8zSXoAYIWQv
n14WytJvkOjVRaOla9dr9/lAeqKjV7wtgmjjKcnWmrO7AaK3UFCbbm7FH6yRtoca
6UKyJy81p1zXP0RPik699Z7TjYXX83Tz+UjihmwipHfQt6AMHfOY2DcO+CplDfH4
0HHozQmXgXmDTnSA/qjd1xRb/5sfL/mXKi4Z3YYwjjDKtSL/nBiczCZDoamUIkBE
4IjQkkvUVfQln4GQG6y+77jtMjoftzbA+9RHttxWkU3TnDg2p+W464EmakCEAAvb
B7m/DFw9zDHYi+j4HQVJBwhwMn+GpOne+YJmYBeRiYe83E+/UnlCrSOCpuKRgcLJ
CNdLEpoYrUCaNsV55j5iCGL7DCyNwSTM+OoxOzmrB/qCkolFz392pNiBKjTHbrHe
dfVPdONgOp8XwiLehzDsmHiDzc5aFbxi7odT0HbB/Gs5C3ptnql+Ya1Eh9jSU7n3
1dxhV79zztUCO7yqzcp1i2rzqwr0L0GRKPE35cCvf74qXKUx27BY8LmeSEO8HHAn
FAinOM2bBNKIZI43fGvyPYqHbud2yHIyHUUEOJOujP8EpMVKxS2uT+uYIzvScH7h
hrBS/0k1hYrTGeTV6qKVlOZRKz8Y265w9uMIp7FzIhXxVCMPN1L+Zu3zkETdk9yX
zxKKKUo+fb/4I9auiLS+z6U0okQHnzkVTp27TIh+byb/GF4gxi0rtgGVvpiBNBth
fzmBDFLNeECTGFlHpEDRTM8n5ox8wdbPFr2Fg0v5ENzx9ERiM/GdY/v4Hp3yP4bM
MQobeLdoHnNQD0r/FzFQlDhCXfbSsVZfVmyCaNspyfhSznPuITAjVq6zJVn+PGJl
TQ/E+YNd2RAb/V36migaH81gOtPY/WWFxXHJ8T44m4YInnzc5lv43RVt7TsLoum4
vufwj7YKsjlC+83C+8dyGLaUoS0CpRLC6FkNdGpkC2L3Oq2J7NeTFByavA+riTkS
15fHfuP58PBqpIR8sRsgL437afWIQrVM1b/Ioz54kjqPkBrynHSW9HX6N9VYNzfm
9mzEs9oj5LTi/G2CaztrfdjsPbA+X3SL22U59R9vAC9obHDQgwOA68JlRYvQc9s7
agQt5NPbituEZC7SBlh8j0Ypo061wBa/MX9ZL4N0pYtVe0oLr3rIInC3YzbblWWc
lrcSQd5C9HMUOF9ijntkppHJssL9sKjs34omdspEj3fhJZjBi9nGZirvCtxHMxEP
abGgOKhlZ8qdjbSgdnERsARCWh1r4Pob+ps68sxYG1R6goayP/IjGdByZkvTish9
IqgDDbvC2BFS4JMDdzM1px1VbbstMXFi6eYDLx3Q2jkooPOO4im6w3McjJVrANdW
04ujB3yXdH1uR0mxbfm31Vd9vxSdn2gOtc0rbGcuNr3cI3AGfBSZb02ZdlC0VFT7
IWm6Zd3Owq8CUUVFSKJ/vw/W9XT9kgc5lqr/7vkW4RCKxfdJfOOEnjitUJUvCCj8
QGFlLe+V4z3MXsFTmQOCkAooKSzOwTWa59YzN+/Kgdf/M9crWgXzkdfIUoUqlEPo
bQMllxYza0+7hnFeq6+zN84eQTYCs//Rtgqy4PK+1LQmeMEgAipmbE+tPDcIaqPw
4QMmh8UVQjDYmKq5tzUnFZGNJotYPNnUi+Fs8TWF8DlO9KjBngq8PT3ZfPuz8Y3U
wBPAaXJDjTVAj5q+1icqBIB7OkKxYPpAHHRXq49P3CWSOxkbnxOVP8DPboezrYH+
wO8DTBwZkX4D1Hc0S288M9ltoIXdqXq9RXPcsQNvjvaYqdTiKDmr7i3upuOGwXGW
SWZQ1qffzCjs8oYwTHPSnNjhWbQyU6OOPYePmGolhLi0XvtUkLhLjvEWVW/jHTzZ
AdteR51HCNec9NCzKelbwIZd5p6VTZoQXrLbvKzH1ozr4C+Ger5NmKe7PW3xSL91
O7Ll2sOdQXqSLPu/xjX1f6uBbJQMQxKMHZvhws77h+rncF1PtVuxYfnOdEqd80zw
VIEuLfiXwcGxPjzRQKt9D4YUre3LHXMB6Rwcr4iAlnw8XPXTb4kbXwUAIg90fNTu
wmkdMLEghv+t/15vcSrS1qZHDeqgD1tD+bDUlstXyOgCZDXv0coXJMpPlaoVmwx/
nxQhuBeqDU70ElytB+3HSDGOztPJ7KeJtdijGlEj8s9zLFfENJhmWwn+TdunzWjt
BXMOD/lQcrLBKv/dMQKM3uaziaXlL0rTJzDP1DFi5raNVncTdVXD/bsPBxfkOcpD
GPWnBMe0QNj4CSPRAl2GAbSpVZZAzhJ7cD9ZzSHhIpP2iLAJ61aG0pDq/3l2+sjt
6V4tv7R2YEqJ2fWU/hIgdj/6ERNtiSeZMMW4oNzF82Zh3PNpQ9+31tHpyxB1+Xi1
kFox7CbCTl7JcMvqJKvUkkMgREjFM06sQBzTYZ7zX3YAHG0MHaGdLOgTU8ju6RI8
Zf12aahXMCL0vGxTbnAj6IwFiMjJVjT5j2SyQoSStUt2IjAwdl1jVpCSEFjtudF2
uzGXtBjLGTvPYddo9JmXZDpu0BviNxppeAP7hCcwpn2ilYcoG61LZ5MCPhxqfyxh
dLJe9yQix6NqAlWD02x/gmyYArZADk73kpjBLdHbtkFL5Ga2Aj1/VTnkcvVibLfB
KhfLAhWhMLnVxYoZVwUSxSxiGH0AV8EIUmELVNBzWEPM5qR5XwP2zqvjRMAOjR1i
7ZH+CAirjxxkkvWCNekJNqSn15DbXBtZbZN1FrjbrymsviH7TssogSxM8+fp11R9
Gz1EcRbR/MaiZVeLchO73YpJDur6D598hh/ADbj/MOrRY3KRzi/rruWxG+hdWgn9
i9JybhBW8sLjajm9C1PyvCHk504LT8Lk+orskCkNhdSm2bMd7tZUqw2EIz8m/bSo
jom6RVT5sj5yRA9uJasw1nusdRiHd1An89eP+qNAsHaf4/bywNamwml/bHFYfPEt
YFjTK9TUSlgq/eZyQezhLtMwTt3uCQdL43wYP/qS2/CShsIZn8Ffx4Pp2fTvuOL0
yFDgIHuyUq2DMJzK71Y73XH45/rZ87bPwI+e+zlJEzZLJgED1vJQzqm7VWSsYCEp
dnFRXQPEXIx+UMF2oDjZpLCdqm5s+VEe0Om3bk103i2RNnUxk/vyBr0bX820r8j2
OF4LZWQcDyIpPhgWKquJ4DI+63G8XxLMZyZBXB1c1MjEMnsQ9E8+pvNAeNdZye3f
VCxMdyqTJ7huSAKK6e5BwRlEJCEjDqV5DqtCjNkLl7MaLos07g+SoaGfrV6IkZT6
Wjdr/qLuDo/SehMg9u8V/GPRnxafk0jEsiBTCFbmdGUQJjMOWdGmdUR93qaLuOK+
p00wmDbD9YMJotHnzsFBdsX3jl5MzH8lsZMdZsOFkYeN7aG4V2AyUe5XDnBwbBFw
fZD7HSxMtwb31Lnnd6V27lxHpfiXaDKjCWazOMuFwGMrnEACXkGxU0EFMj+bHag5
/pBMcKKAYugoWyJcjFgbXE+4GBdRE+/VvT05LzNeiRRBheEi1ShBYq985seHDUU+
d3rH7Ir76OoB6/eIi4GzS9Z/KoTFAeqjXnyfHLXCGVGN77PBUL6RH2EOnUWrtKWz
JadKJJtsaZWZpY69P1j8Ss5cU/XgilViI3OR5G/04VyOdgj9eQPm/rOaxu562IqT
eVtPZzr33vRoVuAVqk7Ulyw9w1RndG7YhNC5s8uyNl7xnuV/EBWy9txIEH+ZD55F
tvGMoN5sZBn0xyu55Wkdat0F0wBotrOIySs5bIgggPlkq0TKpXC/mEeQXslEx2iT
9mFb524svyLdwAk7Tr0jnWp/KBVJvJiuod9+GkknvOy66Xkqa+PoyFXz1r2dgChR
FhxlgJXM+PItWGlpj6+16l+D/QpULF0gRI5nM7Y0DHeGmzkBgUbH7jpyD9d5pgsi
X9aWSl4AkrgzryS05jrVIiT9joHl8d6vW7CjeN8KjVkFe14PIYpMY4L+Bl0sB+/O
EB+rGPcsjDp2C/H8AhDKpsNOe/EwyZ1kEFzDOnc9o22tAZvaToIGIWONtAohEya6
EzbdAzjUbcR0PQEWqY0TqUoq47gVSmT/z9oa2mAfNcTBypFXvF5ohJ2KpErH7qM6
3KGiv2z+Nb5ldQkyrFMC6gTwPSlquOhXOh15qSi6gV+uRtSdw0yxvWrvylqXvpKv
bRcAc+KSaSPr4I/XUGg0/0iGZEl8SbJVxOaP/bajOg0fMA55oDw9IFpb3IPVJoT2
gD9b59Ln+0aCMS4UU91l+WHUqDd7Db1u3pNpE6O2cmuqY1inYCWnV7B8P0vgQhfk
CKZHjE6kfr+fgnTPNFfBlBbGzqE1nqpUWsVGqUcFp7mX+HTb6xVCOEtT8TAwyWcd
mmivMOlMaNDzVP2k2KgQe2wjgJ+nh1QmFf2U0GzC9m9sDxk9lHm3XOMhQHkv8qec
zdeK8lr64hK7j15A3FadPJK7JTwdijnkEwpT5Vpb4p3A01csIUz/g45vCxlInkpr
vqJdezlQli1WuoDp+Y/878hYwgYYJfp86a96oWBi/8U0L5csdDkJs2HmHZ3MxkRv
Ws95fPgGaehI76lwrBaUTlXHeG6Jpzra6voryNTkYiJSDUiRjF7B3nL1KSzQpLOm
J5ZZAfaPJunrEdIcRAgXzvRwUGdiib73DYM9r6Rl8a28xcN9idfMCdMOyllOKnam
0ETMR2ENXRJKh1FlDZwMYCVZFMjuKGA1jPNfkfCa+pIc0coNjWJ26pL3kuwJYmzp
4k5ICrZKt6MjdhV3sBJa/c/MrBomNDXX8/A3FhWSvI0Z6SuBVWmgQNZURJy+IycF
T8xxNuz+c3lpv9slPJlRyTtlfAMrijRw1+nxglX+AJMUIS5DzcKIhfNq5bNfgDpX
M9SATKhlhjJiChqcJkLjNQDWmhtWGd6g2qwbfOBoD7kHiIr4vUWShc0jpcd96i6D
QDiNWaGSphroNOuSA0eiqt/S/7+4mv1Xz+LsqvOzsBo08Lu0WbeUEbr/WYbC8zjB
SUXN55vWGPo5ZqZdUIwt9lnxEJ4z3REoHnCl0m33YE5NK+5u3D24Z6jsA+5XUtzV
1CsG1i2HjXVBAdHvKVKu9/FacUhP0WhY0H71zf1A5NquGManz54dvF+Ik5gGY57k
zZOK08uICC/dGqk2vzuGhhFzVrRrKIFwS6j+wE5FnrlS0zffLOFJQL/0PuJWjkJ7
7zraWjZ49AeK2ji+foR2Dawb22+8fViVzNUltrI5WDntAg94iqtryWrTGJPxUaR6
juHFH/c1LLCsNPwSkSv7gT2R9j6BnInVsq9ecyK52y5gpUmtYzFMI8Tu96RJoaCF
QxqZZHhB94Q048s5sPAgkpd8/TYMufruXOIdCHPcpUSN3Ce7dT2z8AsgqcITr6ba
0dAl6D79Y3OD1Ck9AbsTKdt2Z6/Q1kwR3Efk+dT53EcTC9ElBQcosm+nl+Y4Ogr9
BM/zK63Xr1rnyZMSJvnmXCSVoJWWsgJ6SO1YBq437ugjfezMca0sdRyTqgILttcZ
WwC90akiSkPUaJuf3aqBxSDzsclUnl3S7BBAk3oGL0WTs2JVhd+I9wQImpKi4fON
L+y0ZRuWCSbgfHyvqw8VHbY89eHhWUR6xf7W/SFX+h/Oe1bHDHImCxl3JR06M5Md
2U+lVU+ssGwnI4Z8N3LI28wJmwwXPtoAn4KgkN902eI7pWwrml/Ou+ZjeWkwDYTl
HPCsVF0hgiAlfqIJ2J9rXwRnqV162Kep3NVTsg7iDu/CMKCaIDLtK/MK2EdG/Xem
9PQzYixlVqZySQ6Euc1XI8jYxDNQpNXsFBtHL9CZk+mR5dqDBWWBesynckEHa4/p
SallnKU7+9aG1IaPJum/AC8eIRxLdx3zmjtfKCWA/zWBXkb+UQbfdakoXnfSjfL1
T5O71MZ/LkIVk3iXioZ9nviXZG6XC5hOE15RTN6jBc3UX/QfrmESqChGJatqKugX
nYzeekGVnNPJwlA4HAVbdGaA75r2temsMLk3dLKmoAdPPq7oEeaTp3Wu2RmeD01m
2ScG3BkK5wmrDXxXcINNOAf7LfU2m2LzlrKOkRKCzwjfwhvF3ltm03oBgfHCzgx0
kqBqfnX4XPahErmynQCXgv/1dEq9sCyjK3u4RADEWBlHf3y549G8hHwVowwfIRLg
EbOzbqc+fQRRAhMJmQtaZI74BsZx+cP6t/axV/Occ51j3ADuBkj2A2TaT0SdVNNa
MhjP+Mz5XdZbqtUyQTTuN6uE+XhoYdFuZCIMgAQRpE1e7OW3s4+4Z4PMs3rRpO/r
nYzyOiacdNOZESJBqhQOybiItu0lcrzjJnWysnDi2EniXIGQHHi4HfJARegNjihE
N1ut/s2hERHH29hA+MstTkIa3YX39CGV34eyGCp3pQPueHeHU8HDzfScYUp0EWYz
Xra+0aK2HAbrRvkYvoR+8Qs1NmN1budhss/8dPdFj9GZ+P1QuK0kziTtgshR++LA
Tk9sMQOJ8vtk+0HJwJpgcFLK3/Bb/vrlV145oBa789xYISCXufdHEh0Npdk5vZLg
XYWoPHFWg3gvwSODdxrb8UCehobmxrEgsAEx0/yRilP1j1hWglWX0NXKZh3OOHlX
Gtd+Kf9fedh8T0AS3OCm6kkNyx1XXD+FqWSFiMznir/+dqWfYg/LxWPq8aE1Y6In
slEtDHIRgRhOu+XHtP9o5T0CnriEHhqTQZPk3HnWucM59UnnwGN4G+wP/7fD54R+
9xd9tMa1baraiJxMnr2UMrw4C5pG/AkA8TIae/rovghB6vcSziS8W2KpbJfdTIdg
t9aB/yyXQ3H1+s4nfcP9AHHxCtM9RVE7HBb7F7LIZMOOnBGcvfONkv8g8sIpY/tU
jxytozPY1m4XPmGcLD2Szblh1dUz2FeLtBMzbkYn8JIXyd+h4aVazMhy0qOZU7bq
uRO1ta51Jn57IbbfZzXCNqI7zhWB3OATv43/JSqQ7tkrmdcgUFAgPatZ5vdKvQSy
ByoQj2jCcxxCzUpqK0TV4QJj3fW2RfuJ17Nz4ZjjyRktSU1aBJA6d04ZqkvhWPp3
OGA/KsoXzyz6AJXSKQdzL606nF/Jc8hQq2j7CDz+p7HS7q5Aja+SAmZ7MNj4/4oJ
+rlvkvNssYszFH73rOr/hOx1u2Q8tok+PcbKCj5j4ugqLLVHSnOlDYpMYggy9d0f
EMp1pH7qMHD5ouOJfYtFjxjCSiEgaJFRJ5ShXsEOtOwj69pjSCTqSiUT0lHvPYpH
CVXjciMapxxIB2Ld76VOP0TZOh0fYL6bDgXXiiP/V5caLuZMYlQ9aYTgeUwIKQco
eAlT54Jxj+Yeg2tcRTHSTDW8sG6uyyz5WsCG/P7qbJRM+nwaYgid10v1mbvXH7+p
tqzH7iKST1iGG3UsDNuC+iDNyHIHEptDDFTc2PJZhBVah4Q3iuPbGbZ7DMWnU6IZ
9Dj30286DMoc0d6afW1X8Hzluf1ZmOUbubklTTWaMo1YfjJb+Xm4WoSAIUK6QzPE
sc3+GD/LMH2i71aoywXeC4gz17sDMPMeXcVqTe+hKHNoXP2HjkQLCOh9FijPZqJt
8uuar68Tjvun9Tu8o/XCRo0y0iiRVXyiZhWV2PSB7ckttXuAZ5Lhjjq/dTSB/+nX
syf3oScVAfxMX5KQDIsK6hK0LY7laZSdbozQyzAwoIpODyQVQK5jga79aNXI5AJy
qVeVMZ/sdz55wuLkCSDKwlZngINFrz9PTewnligM4ADWhZ5nR4vifJRIuohRR1aM
/xlKufdkKK4Co1YlUlq5Jj5/kKsnOZhyYd3gi9A8hCEG5WPjuZq9d3Zfu9UqbqO0
j5PIOIw7q5TE6mRQCnh5CtItlpWXafwQYSChqeoif6HKc/FYduxZ7sioCOGH2ydo
A0D5HZLCj0aABHcUs3PnbrXt0Ufy8iO0VKxIdiMpUHQK+E0PGiYNM/doCtC5W+jP
OvYp4I9oSgyjPrwsLzZEzI6z5qjUsreyKAgwds0uZD4jNQUMHI00xJ2OEgiaIrUy
XqFjMUQjfnggKSxmd0LtWvpGIJDV8rw0TOaZrrCrjuxu71t3qyWXRp/qulGXzTuE
tDwokkcpaa7/rpOALUt/VjIK0RDcx/lGd2X9WKpPPPlBdDSresyZvq5zXpD7RmEf
ljGgJFgKaHw3TdQygx3cNmbWakxrAh+2We5lluFcbybi1aVr/0Xe3cyFZp8blDeD
DJwIoYCWUM9VeQq8Ab74DFw6X8Ijv4FSd4m4XnL+i7Id82uQKn2Q8Szl8pvNpN+e
DPMbx6p3G2kDFYXx79NPvyje3Oz1FaPumRBr/3HgVwwxp8/fGZS99inXuWk6wCz+
2hVJFavwsvhvfYkH5IWklaLNxCzthqL+6AOeKGhUZaTJ4NlzC0Xvogmj0fK812Ny
Gnc8qQymMTK7JCBR+qzRJemUerZLUUpFPVmIdYwDAukaLsBUIvg291fDufhYn+7o
ILq2rILv+8PtMVtxsNMLs8K0GzBKVHwGEYIfwnUSxR4Nq0h8+S/NXc8Is2fy0tBu
HHR8uznbshf8WDMGleY6fXfPtGYvXM/yzN5Fm8q2pE/L2MPbARZ3ryDvcOAuhpZU
IM5iH5TCcsQakEUkWvMzz+MEej5qg5QpzEsRpoKWHwLZpFJauk/vn0nTwJdAv0Ip
U8SftnqSKmCHTptMOWDRriZTXQvA9smT9phpsLnJKH+UV/PEUBWc17AmmNu+LOuo
5Gh50P6hoqNAfIkwchTQcFNyOAl8HcNGwNFUWm+j0/VNDs4BA/THR9qg/eRmY2B5
5I/8UnThmpEFwLZoNtG3r2T+tPYmVIxWc6Q9L8h9w596LSkITqsM5EXG/f2Do9s5
umc13r7NAc62/Bl2SCCBMmSiff8AtPTOR+6GKWOFzruPmFtHL4LmfHBpoz273mL9
VFeMUHLe1cGqR80eNnf2oNy0pIbgO6te7Mt5DqEhS/jBpH9K5mN8o3Q4eWZl9H9Q
BO82StWdgPs5MraEb4p2hwaCCkGrTq9I+r1qHk9o+A6YDkDQuFhTMZWIJtZxABj1
wtZ0UmUyn4rhke4N055rzVwS5KWm76wgs3+HBQLAcxjNrfYPePGU6UHFZEE9zsl9
bRmLHtT6O79gxsFH99lcmczW1xf7Zi0DxD8PVHhaxML1ShQMpVSq08VOMu32EEh4
hoQnBxyC8ArpgbOW+fKvWOghi6GPQ4CMUTPikrxJy2KXklLJGZ6B83dqGnlsJM/a
cfpkbAo+sh76M7Nnhc6OIDg2xr9QisFfO2h8p/BLUekSNC/iiraaEVvGNqrbFyDr
FRjY0uC8gh4SFjbloI+xRKoQenrbLZszBwvLUf4AP7CdIu6U44wMafA+UjbbvyyE
4h0iEsyF/q/ovUdGtKlajhbc9johyOEFR74Nai0kCpmWWjcXWVOg3nhfAnwlV289
sAa9Ll2H8J5W/4syyFnHutJ50xINnGZ+2r23QX6moOTexlF/hmvlZxb3+WiUQp/K
9mMDMCz6efKVQHVM57Tzav2lQhSO1hdwvjZchTK4GJluN6Y7Er/Ps8KPaipggJl/
1uDPDjL77eN5DdWg6W/wSOUvyW6G8+rZdCoUgaDuq+Or3Lj9ykBp8oDvNovSg5PM
4RE6HsDevaQ7WMetzYSln/+UJAcnqKQPa5cvVx9ZtD9Wjj+Yl6jNC1S9R9wejDTU
TruCSEaY9RimbvSpkXSyHHw0aCEPX7c2onDQnZxivTxSWg5VSatVgwijafhCGQSh
QmwTbJe7Bq3d8JVeMHuuG+q2e8nY0Ae6KH7DMsC6WqkuYF1k/pdx4jhqXuqh9RwC
9nebbVQsjOmPoFvNF8EX0d6bjCO8ZpvOEN2w6/IE91VBHwGnF/JspNh1UHsiuNVZ
smT4SowoVtZ29B62zByKxvYl/epAvvhdhrCgk/L1viKNDsKgr8B7O9TcenlKlR4+
Z89TGolu6AO2am282/c516iEwK3Ki7voF+3ANopWNvK/yU+KiRtZnyfdSti1WatD
RHqTnIM57R/GhVC0KcoiC92lwOQIDXL+7FJX6mKWmFwRQ3rFrnSTENDfOSepD69A
IAb20U9vIFImGZaRJWJSltYW55hrZAPXZeP6KXFWUWQcF6gShkpwGE5O3aOx2eUC
NjstoBTPC6XUG+53/lfL1735VZpUzDaxi2mnuHYVxSsWb792i40fQeJNQdlBJDSS
ye2I9m6A6V2iWbsBrCZjjRYhO/UUpGgbE1JZ4xlrJdoEZQhXeL7dtTbMBPvs10Rr
mASvXx+xS77lFbvipNmOZ7D+cwOgmpKSsGGs30Ta0u1bMOJ+oPqIHjg4a1s3dJY3
FNxqHnfIntFUeIQltQoW7BK4JiKJH6xhsk7Iq6v0rDqfhHeMD9OppF4jUkz7a5in
0gFRq6Y2o3guEs27ycLYeddX5XEFJrau/IlIlDaclC4pgluHeK4HrUvViUcSb88y
bQXeSnbWT37Vmeg0ZO2bx32xOXcV6l0Y89aISwZY+y8bPAiaKEa9ix+VLBVFpWQU
i0ylYyuFdDm5QQ1TV2XdVOA3YiTAD3d4g1jbqq1UgXmcwwysSPEQDernmvHP83Qm
Qn/mJkv/Rr0PNnzjPTvDv6T5K08EHLKiNSC1OFLGbznffDe3eb8KrA/nfDcB5Hij
evGa/4Tr4uQ9REpjgQZDbw7gcKq8tTBkt57xI0Gk4WBjyl8viGGXGxOAkdMNqD4b
5a4lVslFm11PTUfKXBpb+AMhz1+UnDFw1C1pki4eXzVSKRASw/YlVTHKmFOrfI9o
QlPNZDghCtMZSNeTCJ5AgCZ1jJUwFw5E4IUx0OuqdMf7M3VludjGot2wVEx7QUpJ
1Xb8pJ/uTH5C3GdnZ63IV9nUdToQ5wkGkKHxWap9r9erHsTY7aGbkCPoavXQHyM3
J20LQGeilDYCvtHRKIOtV/M1rCyTQHeAlThOGdpnL1S/Nq3fdP2olthb36EaGgOy
110iOUY54dGlO724IWSp//J9WaCoeDG8MzX+aiYbJdM8kdc8Plx08V3+2by34hIU
+903F0FHkwr0oD8oilv5eH/kd96z1icxXge5GVAK7mcqA4R3nptyzwkKw4zWCXjO
d24nls1DuHiAhmUcZI3EMEujAK1qoAy1DwLAimMnR/NI6wsg59gQK6yzJVSa/yFq
329xFjQ9r01IcAUUlCDjFgkseQWuPlqoVRK4eYnOzQvCGO91bd02LS+RFh5WWV0l
COx2XEzHVBCIX84ds1K2XILVYwiPccDfcxCQWjFraOK5q2Jj8Ledpi68ypbQJa11
Qk97SCgegZsZHI/oXROqVgSBbQ0n7KDvm1P9M+e6W/3r5oM7GGCdGK8UZjyAqVYC
3qJLF67sAclxlx6WGR7/6pOh2p4YvROopvd3SjjMC/xQjo+R13NK7+j9W8xor53E
aYfWJLrTP+27jknAAq6JqRViBDmpnbRmPsaTR14LnYmExsxvOX+4U3O3gSlf5bGN
2wMX6hULYVt3viq/iHiGvvqGlehiy3gfU0EIbk+VA72OrxlQmh+2K8yBEk2iY49I
i1k1TDFS06ttDp+quJbRK+GV+Fa5tpOgFM4o5APSaY/7xt13IO+K3ODN8Wf7m4Zk
pHvxENnNTQj/xBlEeG1tWHvQp1X7xc4yH/SA3fylOZ9JyBcbYA9CcO/u47WlMwRG
T4oObmat5IteFZkygofJDyoWUV8w3ML21h4vLua+/4X5HV7K7tkPDBEpHSxz30jR
yx146WiK0HLUtXl9anxAKJvq3qbOkH3GFj4hDJmL0q0xlK6JuQ/eHbcmvOtbfNtl
xsIioka3Al+vLJCHGSEGR4HxABeIO06fMPq/jTO0KybnU8iStu+itNzvhTF6vU69
wRfi56f5mS66zcIXC7J2Vs4bF+Wi4jRNWCGlVUlDUryaJkn/p+YYknk1HFNuq2zw
XgNOEN6OFzHkcbVYSi0s4AaFtux8RlTE9iCbjgbOIZqg48fO18PlSwQAuUhqMVjY
ZGMq/FPUpiTnHHcTR7iTd2mbEnGrSAxtRlyjZYy8SrYSQ7wD1TIMv7M/ZjJfDGPU
88e6GGhM2taDxJ1sd1glJtOhbEXeYnbCCRB2DNk+GBIW3lsuH5FNmLaafcvuRcle
UMViZMy4KF2cuh7CcdXuBOBf1rO9GMGXbK9acsuUeNwCzUllBJ3Sr5N2swYlZJ49
VkHBH8j3zaZmg8t5CKMlXTCgJnPXfKs2tLxZ3i2dIwZHV4ATPRqVy1jrY05ip+zV
kpM7sVUxlaziAVlF3f2o9fQnf5Xj8vbROjrckH9zzKGXx6RgtorkLKBuM7J43P7z
nzJm7VDt8PiGUv2uXFSmXvpJNzcr5miTCPXwW0wqy63J8RDWOcQExgYalk2NWpD7
eo/mCRBhIniieWm5XycE/b6jDWkawOXW1lqWO1KKjDHzBAI+XMotGxs4Gup63sHg
CSdpL9eoFRBZv+0mqqZQ+cixouNOAMH3TrFXQ0gOUimE2XbmnYJOEgyHzq1QTrC2
+0u/sWOCzYcPrQrJU3bGpetaFcZEoo+ebj1ouWCxSch2T3ryBO9yvRCRTcb7K/mT
MuKBW2xcO1Ek6y041cIqiXJtAoOsuefO6DuGDAdZJbG6ALteafonmZdGlYwv8azt
4fnzpcJFGR+5c4VNyOptVlQcfREK0VWXTNXr27uH2yw8AynkYlK7ELg+gEDMkWer
U0ndPTn8YqNABS0/82iK4RmW/qA9YLyRO9kUG5aJMBZpB5KqhfCNOZ+2cKQCu5vk
fn3FSmQYeoIvnJLckIYTqIAd17ultWHwQ0o4npJxvuPK+hnJbs6kT2d7y5JOfgWq
PE1TEMtJjGIRMaV4iJAhMUdhfzO+HAwlpx1bPO1hoIKNnJZBQym6Agpkec4pKJCx
5cmvT0mk2JPw/ekI5qinp1xfQhnU1RZWrzEEzbR8gRQFRXOKENqZQQ0Zp7e2UX6V
jAnqyNJcc1+d4nwbLA4jbPztRk/uiuSbhrjDHFYPz77IltqaI6vlM68X9LmHD+1r
rtzrbELnyctFE5j886Kd7twQ2gwWz0NpHAuAALobBy5gy10ImshxmkZ5iYyfVfQy
t8pRpLPd9S2JdUY8WFNX66mFQ+FiRHs1r/fCMjA5gt61j5IvzYgdO/N9F3NgAn/A
yyYfBM/VAgyJpnx+Xm9Euq4+gLcjIOfFyqHGiPSaiH1iq8xtwLj1/Yr6puqa0+6s
NcrU2OmhuWrVZj+lnleNGmJAEXi8pjtl6da3jP6A8ryTQ0W0MzlaBPPk3NxfOReq
eFazdWSpd4oOt87U6JvKPFrIfV8veG3y0fHy+M1pKFDNCHEO3QIWw+zZypHsqhN5
Lkp20W79EY5TT41KqaZ4HX1GTdRCOB9GJBnhE4BSD8MY5doLnysxV2mIz+7pPvH7
7LruXNq67x53GP0fdWmGLuxhycDyBMMvzSVOD2Ef8Fj1KLGnCvZs5KSuQEfPUym6
Tbaeo52VHYevSiGZIqbK/JZ2P5YE+WcHGGwgbZTjgtmo3bdNyNwRfpa2Et5rZafP
deFOuePkcYHOI0ZK0lSp91fHKK8/4OXRcgAkQROSqX7x9A5EnGgvY/2kr1w5fjbv
KFW5LjR+TA6GY8P/i/5N7oehVsC3h5ZxP1D8b4Xo1U/GDR+5o981fsGYAu6U/mIw
YmKCr/xkVrmwixzNGYWqZjkwMLyoB2RH53WhGP9r3Dbjwepv8uwQ0dOrpx0F0oKk
/w6Gn7hyFTJDsA2pMfL46T0eNvmFxlSqMTlx0nY71kXM9Bb3nru+j1lbbbJILkRs
Q76PkcxQrYCeUbvmHSvI0u+zYz8g4ryV+6RPj5RR6aUxUwRTwkPDdEnnsLc7e6ht
UD0oA+TNp2TBDGgYNditBQlaoFjI1qlTCArgmeSYPC20uqpcBzci71Bbc6ZtKbQL
AOcvTsNd+XpS5c5gfIAup1l5fk9xvZ/0ColdeJaMDCob563WtgoCQAp0opUPpTeC
rncdetOpHrdfb1ffTBuzIxd/D/OQUxWkUAPuJyExgLge5K8JnfcjoYFVRrxsATJ+
e7mviA+07teL3HBFA4fM/cF5ykO1DTmz3fbsJezwW59i8JMBUveKUjZPGBPQbzRC
05YbI5poeYOez3VhWS3yl5ZJ5PN6x7UNeoF8FSP6YSStyVG4aFgarl0iyI+q/F2s
kzorXyCcHAhnjtVGE6ofOpTkOnDA0/dQuLWyBSaHNbRlVUUyzKHnbWHj4H2L+K+/
0enG4J2xRT/CnlAKWt0MDsdnyKiTiSNZ02RpzfaERVUoWqnsqqCL/VPnV7aZ0nTn
HaZGO9XPFgo6I+m99MicMUSiIhUwNeN7Un69GYqnGIc2PHHEaQmY9IOV3zKKyWiC
dxMiw9TNBw84im7/QuNMFzMELVZWak9EAhOuqQLDxGeeuUxvaONviN8KA8S+N/Zc
30wZW0YON/URev4+yZGbqotXvl6h4cLo6XKkFim4WyXqj40j3CeTc2n+wPe5Hr+T
Hacxs1DnirmmvpFsJb0wpdAtD8yI4erfctLYkEE8tBJ4Qk3CAaFNqxkPmucgjI9D
NUHwwNBIO6HRwK/Bru1I1qP7vh+JOsdK4+pFPg3ZTfd+881OL1OBsJCcjZCasPuh
oMEWwkcnicGYnflSb9CRq1UsRhhde3wP3WQYZFphUQrHVtOh5Cnp0bsCVwPDd9BA
d1WY6R/d855Cue2u9X4nZxL26DXDrOppyq5EhYu5bmn7m06muG7CZ3O9kHLErbsd
JK1r6i1/OTgxrxY515gAHdEMEoKlo0cFMTwgfBAx5VrVe+y5v2M3ULSzkrB5L8ef
JnJgJsBFNJUztPz8yuMmCMDua4MglPN8i4OTYTCLccOMlu13I6muieRb4JGreW8g
OlC8NdLTsR1IU2qfIfUFu2my9tbuTSRaGHuYdOipRFzZ6BLhIQ6o5wSF0aNM6Jod
NZcAyZbQp2en49H6xZf9sIK+DqnWE6Qbk9tXD2JK6Tm0Ut90g+qUdZVzIfTNW2sU
mFpKLj1RGsv3SWkwxLqPmShFpAO2BA/pv1BbYKktTfW5QsUGJP5yVLrmr2nvC+YC
V6Dn4hh5Y1V7NDva55BwRJUeMIFDY9+P3Rfne32fM069R45gEUxXB/NUqhsYNQgf
OlqlRqEczMv3HM82hMnhQkmY+kjm0nHgvdaICvDti9m7yEYr0sIDsuLN31iO9Hkb
BpRFezoXBnBwzz4oV6F8r3WkJ/Q1bshTzxnXgg3pk7/46PmPkBjE+fIlAqlDPIp7
tev6VfMuu0YqhVaXCVJ2FAp42zIooK6A35XZaPXoqLcj5yIzLSLY286Img/TtQT2
flaOziJ9f8wSrNrzxOetI0Vkgc6MFg79NwAycLIWQAFeCbUdwXQMH0SH4pJJDDH7
eDW+Ma/UMWJrCCWC9f8x1ue4t3QSX4LcQg9YnFmJxxSEeqIZSHNLg5S4M3NvNF/g
fxhJIOVVcXX8WVpEh1IuSlvDMgJy5SMoB3Se+F/QCzlX1H6yV7GZXFLCICjnneE4
pAsEQpG5sJ/kcj3Au1sMRiBt3ASI++hVoAs2rgUgJCA/JHuwBPt6JvFUBG++Jlgi
7EE9hnmxQYR6NDZc8k7gcAePZpqSM2toKGOa2Y7UZuyANVUsqRR5t+JtXIITRrBT
26qozb8U0scONUTf2hhVWQ8lhhNpoFt6E2MSU9LJ2pfYdUm+hIYy9bIdauWo92Dw
5/CxjeVAM9AcRiqFiFV+TJBmyENRfIxzqnvaLxZW4tcPUNcwBIArJqSInY7zSBxY
G04DwECR7p4uBRy1uWhV5PAk5A8zQGIbkuuHxQEnXY1dRbEvOPVu5NXoq2EtGObL
12QYVXnlCeK41pNTumelUIQIOy1wuQKHzbPeQb/iEc5hyIo5a+R0MnYetFKWUC11
1MiO+uk5ywgDPjTHo+uMnPpMEbYXYOzBaNgyI0LJg9hgI9QBq0s88X1Xme6YFCkB
ioA83IJ9jtURMF7AdAyd2laILzh80O/DIQqb64Qa6/HSEzSol5Zl33KjOneEDSwd
bwRNHbuVQXLVjUsjpg+t7GkB81jLgm6MDeBZfaepCDUxhgUYlrDtAvsu1sdnjOmH
VoFVClH936JQS2SAkZKSH3nK0MWZFeoT6FHkpJqxbmnYSHwbpk0QsTlRxL2pDV35
IKzGjx0Nw6lplyguLRLzIlcKJnpuof8143mhkxPSOWWg/wZ5g4zpxD4RzJE8GhFf
o2iP9BjIKAH7eemdvh5Tv4T3KM8nahCnNuDhQ8FyhPduaECxUCPgE0gy+SSwb4wM
rYy1HaD3NGwQrSdkSxcovdQasw0QVM5sCVdkdz8irJLTcau/ijM5PwztRSuZHXvn
KXFvBjICFdSbUGdwFpDIGSd035/id8eqq7WlrsSMT311aiyfY2mAEtMxOs2LXRgL
qP1QoUJWDnT54jbAVrcH++7abnoAPQw/+SVY7od7lADdrYrVkhsI07OIQ46dlNhS
olqxNGB/HWWzgyHFOM+Fv2d8vckJE9cK1mtPeVN+M7h1c82gIXFpuK9/DXmw+Wuo
ue64Eet6EAWP2zpPfNgjnzvmISN2B2gJFrnuPqUOUTAOFZnlOqlahgnr2p2dB02b
+lC1R0t8812Oy3cN3T/OjYnaniUV6Q4jn4d3uEjhwU9lzAZzaK97K+shr0Vk4K03
U+5BjqjXZN2jYoRW7fc1VKRKsZSVbAQbAASK/cRPbynKddFfLtWSg9mSLk7osKcL
7t9VL72FTX6Pgm68mSdR7rv8Vqr52jmpvWMBW/rPwzFob0E8wFsJawUdlIaqFwuH
SB+gDDZ2wJ7yL3k7Tlzt9jJCeb3xpodW0ZoYPtpv7JNqiKquTHPNiUASQOPA29aP
C+KnRGR8+2R1rciga01/FdYfjUk8B7+fOHWbhSD9QXgTXT2EDyhQE86uUyZ2OxCn
9bkLcXhGAMAmXTnoeQ5GXTUkOqpKQYG9fv9ks0XaLAlLORs82/XpHO5cFCsl2zMd
h0xibdfKutLHDIEHOe9poEvI6BhfTG6b+5DUaDp8a7f9+exGOxDKqFNbJMHBfujW
MSnjGBWg4xjUc3XWWXFa9vb3KHw3n2AAc7OSx1NAho9dV9YipESTDx54+rZWsHAZ
3hiyEQKa4MSP76RUFsgoJOnqI8dy4o9vk14wcpmKQw9CPCF+dD9ZEmkAnk0ISN3u
CGdk6hV1sMSN6OpgFj4Ie7/qJ+DNwyCV7F0+JAFMjDJJj9pg0otF1yBgQY0qY9A/
3gG7irESMslfHkeec81Y8WAw33mhHcxxq8LKPbiHGkJhE+k1A8zCpTHsBq1fj8cL
T+7ZevfKkQ3GD/wWibDcjS0O5yVRynJVcix9f6icjXZcH3eoaxoHd9X83yq6a4Br
/mkEffhAUpmFjO+KCtWQb3SsSlEI9j7PchdoySLFjRWynKmTsIgQQzLRLdOnEwKb
hxuc/RKKm0be1zd59UVtfPA/cWHlu/IdKrRTsNtEcokcxtNhObw8zcTTSmzCAir4
Ku/n0nYLEIFWyCV4cLIOOAACkIC0hpkCDlJg2IX1DQZdSNucMHf03VE5C88ciem9
37HbDcrIpFsHgx640a4NGF2uJeJj/6bRmM9R/D1jTZcdSTMwC5MBZfj9Gm/6Dd6J
XdsdVAdXHZQeLH80psem66nRt42DHF3HKMRUpcZaKdZzybCqsOeQiq+oQX6KbOFu
wnzfUu/8JCA2hK+jC1koG1GFoPTlAdgpuMvww6a80p+t/oucB/Ymhq05h4W9TgCL
dnB4NB7CQ1SY0wkVtQgDcqUfZWZKb9H/SgY+LJohYMz50EJnAIeLAhM/YY/+Dp4E
WAuQiNbkOWYBs5qvpVNedKYDrosA2k+uttHskKswzUh/aTen8ADbxd8PLo1MS+Dk
NSBv7N5t97oUdupWvD3DOfRV/mIpsQ04WQrgNCD45y8eLMZ/JOSMWFE6MlxvyUtg
oD1/7cUwKOIwCvYdiTBAg81v+zpyoUb7nbl8GSsPhOpABX6J91P0t3xwwrVYYEuo
mHPxNaaFmqZwQzWD/2q8I5qlZW64N6dm9m0mCL4q+v84dmL2lRRAqt7ZGhHMNXn4
TFcSTLf8fqLVTicl6YcffItmoKS2kWnjeeUMRou+Dtaol+gvxNmXxvZwxPUN7Amx
6y7GkLwJOsljBHxPafk/ggmMuWxlEi6qzyHgsK1SDA0Y4KVtERI1Nb48yCUQySa/
visuZkFe5FyEaf9Ec1sjhylbL+t+Qo7mMyjAdUr/0d0TwfpNBWbGqhvrDi9Z1Rta
+ZETd7bHn5Wyz1Izs8HB4OHuO1+tuH/k0VSjWFBxFQ1HJbqtCqZkfpdp7OqCbK0j
+BD/JrpPUyndPck4s/zWLSVn0jvtCEYzaWh/L0rFg+vjfatuM95oVMJHVoO5g9Nh
fg24Ehe5Et53by2ZdIFihvlTPdxpMC25TeUFcAw9URkhgm06SEWzqhfLDu3I3W5I
RaYZehJTP93woC3djpXSBqKWmWTcGg2GawItg7B02bbbaD6P/xz5LRq8fIk8uiGM
xCA7i+7LH09p5VXY32f7nXn1yVV0jUwe0hGBsadhTdA8B9O7x2HYmv6qIbmhuny2
dpM7qhjiaKvC8dn8sAch7aG7HWDR4uKmqzCRXpjvibimeChF0B2YkHuS5NjQnVXP
LmvUkgpK3HD6EpydlMemFuFdCwkv1PqGBILZ73GK+4VCa7MspgIn0PLiGACW/S+H
fbqYoMSDqyyyPr9BB/UdR0CLjgCpmJPmPSJxDCYV7KBSY4/Dhcj2bp6HzB/LpCda
LO0FWmNgE7MkjJJ4Q57oJN0rvoXVHVcUXBn8CDQd6vFSVy45LkNHuLXZyhpSRcsb
VXbjSzaO+2P2RuhRfXKTvgQfFd07r3powB7aCUFwc9kIpcbosetDYVsxN5hywAJt
NDFxhIwTwOfv3hpVMsJ2srQBlLhY6AUvtf89PtGv/1LSgOnlcAWlQdrzwrNps//W
0qnGzA6jBQdycpIZ47pcUV0eThi5rZ1zAzK4XEyXGsu7CGj9RQW+s4LB42ypJxMo
STNMIGuw99gRBRicZPscPDjZkav1etHBXsMR9QsFMiUmKEFRZ9Y0K3kKm1KfOBJD
igt0Yt6TwUxzEYzbjNE1rNkXqAYIp8i7RtLegawhL3htiI1CVg7w6oEroJdCNKbC
ymhxwJLVUs5JZ9kaCBiLfdNsi7AylL59elBzQYmtnZnicuUoaO/2y2NsKEbAXZ/u
3ln4S8cqqtcADn4VHZEqtLMYn2i71V04yH7S0rVoY+ky/et9IdNrUOWt+RHrtnm7
qxfC56SLalnMqSAH2LB7K6unaTYXSfr+hkA26wz3TXyPV9EJbh1G84q7OB/31BYR
SSWmkgwBWcVzDZs8kMdROlzgvK+QhVhwoUIjfwSdU1wk4l5JWjQdkfl1OzSPiSJa
9lUf2/ypMEhFlRNxNC5kU+IPQREL4sDGepSLN/7T/2pPWHbkuxsdP4iHL6z75UZV
IiMSu/rv3qewAnH1AwjHNIWnWPYce7LcJrB3fcTTZ0yN4qIki9000E4+mf476H04
jJy7Gr9JYdkY6Zl8pw6i5Gij1zqFhoF8357pRX9oHuPbO/t/iCO8WdjEh2JhNceX
PuwtaRREc7SpdpCuRuIeTy1M/W+LyT2a5UWNiE4WQCiQ4Y5vFz8ZhSzUB5r33XiW
rc+sIOmBMNGrwOQV3OI2OLFnvXL+xLf2iUYStYuhwJ5NMRREA9ZFOE2GqHTNHht5
P6c3FWxEDRz0iea/RO4ox8GiuSaaUdDqj1i14CG2kO5CAPOzrtjRnFHSyCXZI8lo
6g3exDFIm/mvbGcuob6Xv5KU7tzliCRbI2qhg3UhegQtUSgbZhlIpsUS2VQR3tmY
lvieV14Ii7c4PZnNlB/nCKeINW9nJeIMXa8/Nv1lIibbAfZWmQva/ZoXbmE0Rjh3
0jPTbAOVR0l0X/LJu+4vjYJ/hmOBDe9FPvJkmTz4LCFeDdz9amrxavPYb0UO1MBE
cXHWXYl1SZ0eMnv8k5NKva8xhO699Symdx2tgR9wS9/YyDc65Ref5VP+dV8tiRh4
nsEi7t/4JeT7Bv4pXdTkNuycbaI8VVOouwo/bUjTwvxkHmiKCeS6ugLKitozT+xP
UgDFs4zpklw1WSfWnEdZw3Ec8y2hOe0QHuyHZyj4KqjaqlTPgzsetL+aVhsuHhFU
RJeLUh7IKJcuvRB2h3Wc2wQaFc5HUuSdSktxgVnTtG/IO5RnPJFjppQvCAqWoBGw
/yFyzO7d7e9qs+ndFeMoRFigHHlYZjSdN75dYCVrNIwRFxfh00CkiuI4Ug3qjRUm
5uK42hPwX4BNnV/RJJ43zYqcm1XvAJthbbqcgmmAwrBoqE2UXeKRia5+LcO8VF3Y
Kkr2iCV46RqOWKzamtQoql+lpl3qFZkrg32D8ltw4DXfsdzlXUZ5hi4Qd2W3BpSn
uBT4wA3S8i1Twkv8jrdxpIusAv4KKRlNXmTetFbIlJ41M2VYCXECfkWXtVmgmNhI
V39ikIVS+MI/iv14O6hV1RocSZrKThtOVssuMFoov5XNrAlzYPxekWADD2cdGXM0
GQlt4XRGIH0xfsoRRsIWIjVuXSP9emM6k5UDvHSjPW9AbJrodqo0o8rqIvGiQkMa
C94GMhlQdkZnH/Ettvs+eDJb9/FI/RrB6YyclMNriuX7HkumI89tn/96CLbeXpAf
uNzr1c2QTqdmTyiLoiL8ywP7Mr0nqs520XBI+fpnSYYLXEzJAvcAoUcjv1STtsPo
O1cdIhUjeLj03muk24fkyvnR3yTW1U+YsFDgB0frYeaioMoN0A1JmREEpqCndqq0
KJT8ug5mm0yIIUiv83KTuHNzaRkgRwJXIodJSBhoyrHNwp1tdVIu7m0sRrzocQNS
N8dCycoOIpOQxZ9LuV63Y2ofI7G8sMp8XJGCniyyjj3Js8dR4DkE6dMLKKOVqYeL
NxHJFYIEFtWdL2tDAoZmWDUFH725ox7HKczAqd5PvZiEWsTnXJotm8HqJvx+jbVV
vMRPamd1M6k7yv5xTkv2AE8HmL0xqxu5paUgImd1g7AM3IMiYiPVLDI8DQ0uhYK2
v2j1rHyJ0PfmIYsYTPLoVyy0CI09oxrnx/wxLIfMzmYKWKc1CKKh4jo06oVhhA/4
ZGm62jxUtlIgAgImjTwe+lIOXYDJs86SeQWdvsMhnH9BnZ2WwBIw2hC3bT+4FQzZ
1kcl0HdlpbQIYYlM8fINkpKe/0LlneFuGvkMCLk8yA/TIGyvj3W+p8T4cj7eZJ24
Ip2CoK9t45VKZBQp2h4j+FuIaOgfFoL0wg+D4Adr09HCk4mI2FmSAC/4DO/i9MU5
rJ4eBYE6UOoRhvWo0ONkdXRGKHAHZrJ2kxvwR7xZCe9egBflGpA5VKiEHM/RBOAA
7btF0ogvRTNf582PrIKEL0EFw74gP6gtRAnRTbYv8sMSP0VaTRzmcPwxn/xlBxmm
bD3eeR+Cv9RTEOKjiKGJ1OdN3yxP07LmpJF2nULNN0mND4hwHmnYrPS4g93fUR1L
qoHVznCBXRdLnpMFzHUStidPFahhNg+7mL90G/IA71vkO9JSBvwXbW3HKTsN2ZbI
sB78/YIqOAyuln6swN7vvy0P5AXp67S+uZhtpRe2Ry+n4cwZR0mwCNlgObJuk8oV
/Ykv+rvUcZIXX0O4xBDruL7GSNrdHy74RLIEGCHXjeYig31OdbbnDxuQsvyXavRh
5ND+2APNp6LrzuscaXZIOYpKIv3UtVuHQ4RsirQit/aUJug2/g/UXtwdiygj7/p/
9hfH5IfsBvfx/IFtY/+YGumsvi0pSjG4w/APCYjLb+rdXKKTLTqRouFWwAwYvsxw
QY2yx3OD6mRIbRewABDvxSABflq9b6/vvk3bAHz0nAAddc9T0sPiLa7z3uo7nx2K
diCP52n6kT01hOmCMNjyFCjxaAn+0Ot2tg+6/7pPQViXe1g3ba3mXDFF19ZQSnnc
asvQPookQk3YWbbUQFrHk8v8lYOlnizfDx8IdVS05sUEoANHQza46TP+yRRuHQoG
O4h8iuh/QXkTrIEj4fk8VEOn+ckNvmMhplNnDp0TZtPfyqxDVenHO2O8b5qH+BAp
7Mbmz1Ln0jFjMwiUY6XyogyPIE7aULvSJheSsS51kw8XJVQaODn4CY4ECCXp9HhZ
z3qcoLf6JR+IwTCuXIhgXTsxD94P6t1VlX2YxBFB6IUZS1tDAN3fBoaAOUh6P6AU
PQdq4jKa0cl7qpCpmEhalz23f/d6GCYFeWrR33YZcbK3cWoS9ZV3vhMoxvt0dzfZ
KrFzNeUOS98plGuSfhOn6i+SrRbXhJFESce5ODOcntiZYmk1ojWF3Q4UzBLGT2qp
2iueZHxcM7/wWzHArQOjIIsvqPmYrlMjg6Dvm7iDMXBf0k8rR6YRHTtVCOor8DKk
luMPaMxF/1H7LIfT+9aE3UYpHDq22m9mvPJmqurk5HdbUASKmvfZCSYUXV39OC2v
53/sUUD22/u0MLr42Od2GFH/7mMPYZ8lwR7AxrwZkj1EjSkgymABeTY15WegDisz
MF0SqCp0M4QahN6Dzqs90gQIVXWRv6osGF/DOGluP4QuSRU0D3/5izjN9otfBVdJ
lMROMbpDLWzEBKJfhIREn+a/f2vlAkYxwClHTiIeGDsNSP0VDK+1OUjr1d5ISCxe
KpKZ4c/FaE0N+1Y5168i2QOYtfxw1FORYbn32b7zZGwSNUE/GRH1KIJmjBZ54nkK
Q5N7prAlry4nuShZbO1P9qZIn2en9YHuDT8tBttKZG/6065ojax98YJ+SzE5p2Ci
Otx3nVljbgCjU2OWlPnsXEZR8aSxQuLtQ9Tc2FczU9IWBZb8P8JtLkMMypbBz0hg
z1y/9yGQDQT7zikcSEnKb93rHUrz3EGSlc9veks5zL81tJwrb2pSHdBkFpK1udkI
63Ko1gMkMm0TKOhPlamLuMlq8tMUjHyUmBK4p4wYNXUxNJ8CpP3cdX3WiNSzI10+
zQqdN9apMVkPlJNA2VNIm6eAHXzLNi8A7SbwxQpmPZe8hcKrnBK/nPltcEoRso78
YthCRjZLjlH3VwUmu0uAil/Ti2AEcvwaJF3lGu4n0na2ISKk8fnP6N61KFG6raSc
158lQboyGqEFHbF2cnTHyR+xO+uOMcZpeCZBzmsJHETdk8SP15acIjx2Ohj6r48/
RvASyqG/IWVzkusZ4piM0HNCThImS0ughwPoihkxv4e99/1f7QjBG1vvnU3I5RYo
ueIsnbIa2J1Tjfp89CreHleyAVFifRlud1kSaMYgeQGsG52cRxc1pDy98bdP/hLL
hJlXnQ55nSwOyiMR1j7Sc4PgzR6On7ZGbAzVbHWs6Nh2O711h7KsBM4+TVyMBTso
HrMhQsGYmCt75iRgLbEnOy9Yx31wNDnzzndcwc15cC6iaHUnl89/Nu47uIGqJT1y
bXSi9EOPkXgrampzB2TC3Ia7zHPKVheuu1CCO6LEjJkFI8+72RoOduJ8Q0PSahGM
liOEZE9jfiGFCnJiKdiO0Ikq8E3oQXQ/ffa7S32mdrc6NkkhQI5yE0ygyRyAM7fr
6/IifbUQ0OgpX5CPpfb5cJqQHohuxWsSuoQBkIWdXqsRMc4Rj4GpSl39U+ucpr81
66Bt6zPk6HJK3Nlu1Ezyjq8fxFZBj1p69G3TVMwtfJyZA8VWbSvP/3dwjCJXdFU9
e4i8SYA8T8rBziOh/8KG7OV8+JqBMHznMSJPuhCFIaNYegRWRFZ4GNCk3NoJwAEy
DJXberCc1ji+IXYi8GdHHiRZJgF6akn6hzpHJB21RuWPPU/bFHjZZxvHIovTNPn2
uqE62s8T12LzRLF0IL9swyXeFlh03HW6c04B62iHcUl5SO0MhIJaOgkux31kwzNm
6psaG8OASeZdu194T4BSfJAPcidyxCcjUEc+JPAh9dSoSPXAhMNsSRLLp6svC3ev
ozwmLdppxV74wyUFPOx9Wdd0x1mioZYj5FKAo1Jwfx0ioOtQtnkrIw14QtaUv37q
WDzuecOqqGlCCDMQBF89ZEoxzK1JPinQ92DHcAR/klZIqOD5Yyd/m1T0VGwYB4p0
EQWfml8fHUc7qsoaFG4iiU3uozzsXXWdlENEBgljEX7bZJclPWOGrqfACaeg0jay
1CfzrUJr8eRToTZSSr3z4DLJ0umKc04e41L9dfBg8sjcaIwZguRIkHhZA55iAPG5
GrOMVa5xOzLa18PgbnQYvlU1yk1S3ecpRa3e30+9OoSvN3PoxADDpfvk+DOqV/gF
wtUTp3wC24Jz1VbYZ+SrWXGbhKxrqdXfK/jkDlhgoUJKqwtKyi3szZollwzgR7bp
3xf6IyJh8NJ0dghI4Cs7Kw8KcLVNuTCM4AxHNWNrvGh/kGBV5dvO4i6ZxNyXSf0u
Gxa7JMFR/uKAq2zWif8AsNRd9TidEzzBZjBOBTBJ/+7MrA9PA1tVpx7TwKQURWXY
kRajCh88856sVm8LA6MZECc3gGGjXUx/tURy8KY2R7B00KM80LqL/xMYcU0YITrp
vKm8qRhjNuEymUhIIHMoSxL/fwvdjfygWeO7J3XY28rb8lnz5Y//WXWtnIj4Qr63
0fAxUeigH6vDfT/kvVM/JQD/bdgglrbq8ebux6PDqp1P7JkYF8FeQeoNHGaNys2k
31cUylresZZ12HxrZVMtvs7XHmsKDK1mZAdyduAJLL8sJsZ6w/zpmDOsPvJVqMCq
F88qPway+DCEHPZcxWKuBvR2TdLU+cHLazh55NQsDEHGssM/ALqFujva+KE6QOgN
1Nuk+qj8KzNtQXTszb0oFWG3aDXwqJZIyV45iSGB/TflMa6GqV/H1MvYQjwwyM56
k3rcRMJyQ/jcxk56cipH3hp4AqeP3emeKzRwCGOCKbrQfqdnagi4KLAaVk/xJ72g
HDgp7+J6AO99WaKeJsUiC42CqCoIWs8qIjJoHD17kt0UrnCr08xzxiBh7gcBl7+C
17wdE7DjyccYYjz0B6tcIKk3Dddk/SMfWE5gyh4N2Gt7NfKPE0Qe/GfbGVm57KE7
zfUzDppD/OfGTgGvwT/rncYZsQIUA9iHRPs3tVe2xDIC0CP6lexR+Qb7aZAmaN0i
GCs1Dyw30q1Ym1zhCemJsoFNrnIHy1updHr6LEtGh00YHC/y2gNT+EiZgjhCHqRa
7FAUvhaXMOgFUwvveuFspF4bKVgt+hRvKePUalr1JPFTcEHPuXZKrV2TFXRXSheS
NE52YBA2oB+dUXTGTQAwnoZkwlcawlAeHfIFbPZj/T9Wbl+lUnlRiL8WnnaF/CXB
PQKHZNAPoDjMeOzLvZpjjWSX4vUdK5mt4/R6P+qG39KUH5aXzFSiRKCJL9gA+MfJ
P4Bpq2fbrMTvIeIXUDLp/dC7SsEhbbKhFkRKbeL9jluACJxJ1BQNwj5UH3FcGgem
o92x+6hcE60HZmE9PfSz+ApE7xIdMKLNSmb2jLVG60Lhs7mIBKGg0Urukolzu98q
j+ij4WZVjm0JduCJYkzH5orXnVvW84r458O6qlsJoSL03SvzIi9L1ozVAvlGnyI7
0C27n2uHmtEd+uGfgvQKn2U1BOtWDHnTDCFuiFiA+NiAEJi4PjQJJ1pWoehG1o97
9vKIXONCL2m4MVWr3HOqsw1WYxr0tQD1TkRhzhAisiei6l94XdGsBLZYaC5Hv9p7
dA6zCN2tAICDpDk48BEv4swg8jdECeav/orF/49Egd6qIoy/pxwbrUmvRs81a3GZ
efX/x3qaZwzWiUbbSoJbuGIIHQQ80solqe76LGhhft2plH6QlWXXUCJeKAxG7N34
Lggt2X8lJy/Sh7jXfZN+rBLs+8O1fja/bGADYrFDrmhlFuFtDbbLXyWH8Eg9WSi9
oTM3lqG5ZZrQfUawF+1Q70QsSiruzmFzssxHwzBNqsvXGFtnTN0aQl0rtAWD9Ko+
Bki41v8VwiLQ+GQUhkCRwUDU8OYseR2AjhKdTGdbJharNiPUw33MFgBgEPP8Eclj
YiAiZcXn5NREGv6ws7UBxtNqjBmUryUaWfPe8PUvDM9K1FZF+/yo0K/gCN1ITrmi
UmGRlGiY+37ispAHkJ/4m3K4v7+9+avUUqnzwoXq/M+gQK6ID4iHmuLDnkEeIkjT
3fOcs4PhJVUZbYZtSbPzT2xovaqwX6fIL7dgcNNNoAzWrJbv2xM9Ysttq93LxfCS
0ZbxeaKYNwz7co8J2u12SVTDyQlM7WmEBeiVs1XR13Y2xTiy3VCqwZ/gxEIqaWk6
Xd0V0CESAtf6xfdKBxANCZsbe7EjRbrgjuBB2vHaUtElMnkDwtsR7vzuxnZSR3PZ
s/1PpOpaikcRWTuUIAnFrEjba7jws/Z3TyVGM89jf/1R45M8N09joiXXn4hyi6bu
5US15w3irMmMX4bjBbtq1MbPqhMd4hBQo+btHtRcMRBrJSI3nYSrtzSZHCzmU5he
QeMUHp/iNqCo4Y19BeNkAAbKqB1+RKEsMRiOG0aR01GcZwnlihfPgdI+0NZsuQTZ
jasw1eIMXl9DTwYZWar5WS3fOVS8E+8CmdjdR6LlB0UNzg1bV/05SPlGFA4jWxKC
Lxa5rM8tQPYDy28gWDIIYGp8dMg4aoTHiXqobi1upgWmvza3epN+ZXAe9UMc8Sdg
ICgRbmnBJ1gVYBb/pTeeYLspmopP3uZLlsoLv8gqIbd137qRODSaR7f9ZBLyvSHC
nS/WFzVC6lBjD4SxKRTNRBU1+Yp7GzyyULvey3+FnqEZfnDj/e7ORcZrhJL1/KSN
/kOvjDiVmiGMQ93Qe6A1YXwVdFelD2R3P+2rkN+GOxAUcGbBU8Zb5xAJqrk5yrwh
2LUY+ri2dQ1KiIrsnyRlz4CAL6EQiDzhfgr6FWhiyp5jIzrcDZ2JdRvJuRI1XbEC
oRvrtCnlMLHvQY0j0NPRuVo7//7DvaVtmrborLjk4WwIk8v4MLLD6CORe3tu8CDW
MpfCLE4+yxQIGv1sl+E8aBa0GlZxjJQgNLe3BEkSDovBxvP8L22u2XQLJZxbMqyS
jWBj2kzDKuNoDGzYtoWN0l6XYxY8V4z9ebQgqtqb/Q3nz3pjldLhjgvcgz3tDneQ
TCXS6MlVOGBNlrSiTGw88jcFLvPm5jHi/Odx09C8ChEQWfUfLBq5eFiP2I2lsyhH
3F1GpOFAownn05aVir7hb3ILrQ+8+IxxO9W93M0Z7Rs7bMGaqipzjJRn4ocKW2EB
gXynBPJa94jBWsuIP8vz/4N/ELwD4Ef4681lCdEbmjKAfb6oocu3yQklvyOgwGi3
kJxIvysdJpP6bBiA8xfTI4RF9k7u5vDL+TZCWS6UrMPLnQi40Dj3MUN/GYs3ymcy
8jVlWqTFBipwCbfM1uaBDGIJmrSRXner3D0ZhQqe+mO6CLitF7ytKOdvchruYVAZ
GNBCZDPc1tp1UWfQq0VvKBmrzaUcrtB2xmnbQ2mCqbHlFxhz/FPo7ojaMlxkgAgo
iruE2ulCAPfNSpMLuys/xOOzouXf506/It6bd7NxwC7U/3jvtPT08ZA8fhFWuBV3
MzL632Kcdo/uluNWxivDKR2q4J/xZUYC3YpMAkDmTN1H+zX0W2hHJ069O6sTePDb
Vdxw2WI1mukLk/3SNorMryUWTQC/HjYag/FogXnHtshQm3oX+1KsGQZfhpwM3gIo
P/3GfEYM6sYiNMk5KLGzUQtwQCAbJvLE1CSXe5u6Kf8y9I+Hu0FK6+4rF3BJ5atE
2KR0iQVjEJFS7NkqRoGfJGcrxtpRi0cJnNx29U82QJQi6QG0rlnRiUaxLDEUSlQL
s6npLtbUtbLo1Pk6687sbuKQAzUfnb8pbrx4ssyrhHg22aee/nnr7eloYnUfhwGq
3ksqXo1ddo445OQ7lBHaXnTTy4skLdGZDa7mStrg6ztwzyVC1nHGTgw3133NJq6O
buQnWSh1cuV3VPJCYMunMep9pjWVDjMO4EdGuZ86hEczCCd7V/YO1XsILCRx9VQ8
VSBqaPxEaynap/cpT/n2Jdx5nHq5Fy3KkauJ/cUDqYjN/6bBHeEDIQUrWerulCBm
dHOn3p4qFYG761JvstjRoQah8fsQi1m0eQWA8IPQUmsVZuH2uJ+6AUjpieiWOuCr
pGvRcrhdl3EHpIGEw3cHaaV1BGSErWVKz+kEmkRIKAidME8fyaH5dYbokxjzyW6q
/9q7VXZ2CzXtGOPgxVdeiECBk1Y0atruFburriJZ73dx1jhX8L8po2AB7WAoPpkP
rBvXwwJT/Js4fvj/VHbZ0q6Q5JOlPFSOetupZtv17gAk7JSuYWdHedHnHKan6FPE
TwNU8xLy6ljKYThjsRubJ8w/TZv9I2efBBVJHqEQhr56uM9IGPfKtwXgyOMgPhaF
NiOf0jhe/Wa24fT/264ibNZZQDuJWwFEhj07PK2WkB2f8isO7fVBnY/vshbJfCiH
iihGcsBOosH8Hi5I+O9+mfTXkjS8Eyuz1ARLEp2+DOlQ1X707QM1mnnHM5N2ldfL
diJoA+bcGvTe6zr+k8ITrFNvqZHMrCR5oUpbIrTsa5yww0kJP/O4N8sHl0S6Gj/X
iXBiBirsPzMeQ57BUSodTrxN5WRsikrPPs1kqDCn9DmNOjmbaVZj9GckZWkOi9zE
CbJlsnLxjzpjMREQki9dD4pYIvLRRGLb76QmoQ2XIjIJBqhTwMANjCG8mPmQskMA
aLMi3fVEpBYQ0s9JjAzectuehp9cfDvevCoqjxPPIRqOQpLTWCU2IdxjP5V4AmjV
EFydrti8KZMU/tuJNxU+TTHy4201A24D40iFyjV/7piVFzDWDeMUoLXTnCiQZc/o
Efg/hFXDEElPrzRUJjR0YiDymorDZ5/R0mlm/ZE3P7CJZ01BKigIGdZuKyJY29Cv
dGM1bju9d2xaBnALsZfSio8QFj+30sKHh3tx46xAYSfz/2QL0XY8WvmK/Q3uN9Eg
ofDL0dCfMtjXOmg7cNVGEjzXLFsHiYkjYRTDtR1Z9Ty969EnWudlV4Ysl4n4xGGN
SqHGTKSp4BU1nhHruqEOE3ywvMe3kxWRlcwuzf+6GYnUlPgZjJkSbHf4Xe1PYnWP
k+OPJRmQzUmrmtU21sDErGAGfomr6Yt7VexMEKfgQy2h+4bphSv/Nd99+uhNTNfz
SMj4MimoQTbUa4lUDY/Nk8q0ran+ea426X/3Jj87oRow8z8Gf5DjBjxc5aaqP8Jb
Uxk5TWd0uAicWWYgjrwhr0LuwSXiX0Yowr6bGhscQSrIbl8cVZxYONIvyWHoTfYu
lD1gGz6GK9jTUoo89wZpvkXuoAc8mvfeVfGUHM8WCrZOGFpMOB+OEeLl6IzAX4tm
MepYT0uIeCzoF2HD1Ym7lSpv6w/lCHXYOklB2/0YMlGezDyf9OBBMPDYr27K6sQT
WRIf0i2Ed6c+NPNX0Gq+TalluJZNXLlP5UvzG5Nkx0X54S/Hk2jDSIbqPYQGLAXo
YOh0cBSShSSorpxwUHSOJ1kGDDnt/0JSjuwiwhNw5jA9Hdxu9M8GuPkSvwHDqKhQ
eMhgxo5tTxoMXMainIpU6jCdgTpcYa3QUXitQ9Nuh2p5Rtnnhwbr1Tkwi/1rcR5F
0kmMEem2ZJnoF9KZF0y3aiYpA4Zgl65qF2y//XKqBVfZ9hd6l/dbzN/hosSH2s+9
AW2ngt+hdz9Bu5KR+dRWuyQwlIV7IqegBz8moi1O7G1EVODkF4Zo/I2NK0A7UAtg
KgP9qviOCcVNIgBs0S+C4iKogb45OS3J2rhqw334sAsWAiPsLwyl8Wz0xtErOVcR
W2fnQDrdJdVbNPSZffBdef4DH2CDqJgbsTfUITN24vEoPUUUiFfU7ei4KP7ki8sW
BBclT2FTrNDz+wvWzzvbOrIkgbmI84EGKcjXDjAvQWQ3vwchLk7y8FohaOhlUnqD
hVP9x6I/zUfRMlAGdkYlSAmRvv8ovOOf8HaU8lgHh+izp2W0DkslbW69gOK6XnbB
YSCHT4bpt7IQbctKZOTAE+xvPV67HkdElkJHmXaFebFFEHGGtfgszauM1c2FRiSX
CSXB8TWsZcm1aHg42kwgNsF3rlAWlJFcPvY3jgAKqszehVjVDxEfTQB+A7jfiGdQ
UQ7XFBXq70/S7tMfvAL/qF2O+o3aRcl1MGCseQ9BhFXr8g1ErS+xPBzvbkBlB8BC
33QGH6DC+RtFybsFHi12HuT+4EBcHsnd7OIFpJmRreqatxXVTMrjztLIS4WmGLsB
T9pNjB5oBKmPOCiKRjJAIZ5tou+7/qzi4YoTEZX7U9TjjQbDtRT7CccbW2sGtQj8
pAdNtGLtXzXH9tiQo+Clvegum4e3bJwSKP+iaNtTDXrZv5sfF2kOJkgQaRUnKqeX
xnoMu/xPivVsC/Gh9H82ZFAN919MuyVZSmX2927U/8ehTDtUNhucx1A3IyD57Ry1
Q4pZ0R83hyMSn3rhCsOk8cApzgJIkjilLoi4nTQ14qMv6m3qk72PvHkiiUmKpF5M
4NBcnqkRENbTXsCjGo8vcj93Iv5ubrj6R+MtszaL8LLxfsJi9lYuVTwZf4QGcf1F
mz9f0CODSx96uVn2g67P1PGU52U/Ded8bAr+T4osS6KULM6UKBoVGosutjW3fXz3
abTvyPy1e0WBnP0JiLzdi8WXN/zNcK5cElggx7umJvTjldEeYHJUHHXrMnWpsI+7
J+vxZ5Z+zg6bTyHKGwgHmmb9ls19nssYyV2MaBc8H9Q/S08yWjtJEMwqo3FSeOW+
EbpF0w1b4Xpv01m5AYhjBHbaS53A9gxIoMGkbLYrjbc/ndZUSYLfrt+y46ulAsgZ
BNSLl9auEEuGlO0+rHx5dH+F/aHJ+AAShllHUJWA3ervdXKqUDZW8COu7qYOMj6p
gb+tIWwcx6Acdjh6V4fHKHt6qG0os5T1bVY/1k6lTURRTy6qbZ/6wwHzpFAZt07O
55q1c+OwB+ll4jwSNvdwmySmkNJ6HAY/mzz3MOfAgX5kfkHOVnN/W8E4O7JtdMfc
PcJ09LddQo5C5ihkwQwuN1aWOSzw9fmvu7mwg8sj7bSP17CYmTGqqou4FMvcI5uM
xCoCBIRG7J3AVg2thrKbOFmsmqdLbZ/rJTmEs28g1d1lEdR597a19gDLq7397las
ASvaqVaohmSzARGc48deKnZGdj+Zj6Q8s5gZnuRQn/ODy0tGAkIbVtk9HGs4mp4I
9WOsrUH51DQStVoNbIea6MyJl8PyEX2EKMIElHGxYNG+I5nPQSO4ria4CE8XoXP/
1FdxNSY2nOvVLbKYIFndvn5bI1dBLkwu6KpOOyO2CKfq4cROJHjeNbUiXbZH2592
9em7/JKON0kvQYVdQlBvBMxZkyjW16x9d6sBd0NQVqoMqUMVkOMCC2c7pravbfGf
kgLuovRwiJYiNyFKnwTeDarBep2RQUh3xqwc001Lm+tuJqHzbOOhD6JERzYwdzb+
W4s+cZq1blBKdxPWNR1KozDoS2MKpV4xccLgd1UI0jr6174mU5kMcNcUhrgD+zWh
St5ordiGIuJcNeLKS7sjEJJifozMo5EMDDbRZ/nrVYmnT4qTs9TMzcsM6IxzOaq9
Xa+2i5q7QVcr4PTQjLklqbUdpKYfLI/+3o4MI4+Bj1rN3Fsynr8SMUZ0/B3uu3/3
ms759fUzv4KvWnCIGvS+UNZ1kPIPlifsgICEFEFLxcsFeilciBxz8s7+ouEqxdsX
OogABv8ROB1WXjMJFCSDsXzvefd/dg7tXvTD/U6wqydkp82DfvHFMU7ERX8myEVK
xnTrvBXDtvJqt9jvx719ykom3fQKs8hab5/pgurfcn4mvaVgJCxj3HCVbY4sUkej
+Fppnhy/2VbaAQokdiEmHMUzQ85nA4jz0RRsGniq1Pn+dFivbeFPpCTsASk2qSfr
9ZPVxEaExpHqxK0ooxfRtbQeF/YneTYPSaBneQtHOhMRCE0h3QOcWbS0kj+plwnm
kmK/sAO7+0Gf49G2Ah7U/Tn7mAhMxtRMv2I5OpwKqVE/kDUcv7IZF1ZhCS6TOHrx
u1p7FrCxp/WugIYHKwS0Cx/DMRDMdB/O2mgikFrVYJw0Qy/7WaIKHvjlrBQW0H3K
WcmpnDPCL+uH/IN0wZ23BhPQtpHRQfjf0gEoi17a8cTzGSAoooMsomYuaCJDtloT
byd0x/PlUzR1KHQv+3B/4eZi56hWhBr/mcIopnswCfhF6fLInhe4+WRFwmxu6gWF
St2xYiMenY9smQ/chsFDYNf0g1R9YILXVaJdDNp6ABIE5sd9qgwW6oiBxzxnSYOk
F/N216shlHCeurCmPLh7dcY/3VbcS2oNdMumE6epNOzOysQ1sYLZr7qtqy9m3P+D
GnNnfPJ3B4NpwqO26Jj1A7BTczBnqq+ZBONuh6jjhwxEFRpMUALlvKI0x8OSx1zn
YDDZpspWTNe4OEEXaQXGDqhDFSYtHI+IQY93PLC+5nd1c5Fbz3MrgVPNzHZYpycJ
lX0c3TR+3RUPl5hiCyXrBMhB+vSMwZDtIDtu2hTJUTru+qN5FyGixH8JLFiTsdrJ
mEjdNKfXsZ0uv6FwFo6W74biUtNtk/FHBzzDt9KslTnZljNOeAQTwhoxSKvhFwMb
VDus0U58R168y6Wec7NOflJ/Fqybj5vqTPhyv79slemCWctQR0odMEE8T/LK4Yyh
M2lWHoX59nZpX30DB9I1lJqgswSAz9Tfhp3w8ATPKVjJngERD+7dWHVEoeMAF827
HGsU3VITpvfOHtGJf8orBBbE4eFeCmVh6E8rDeGmua+AF+WV329mMi532SXXxyYT
98ir5rw0gDxla0CoWYVD6Bj2ZS7e+YcX6/lqRBFICNw465AEe67+Ifd/5LeCYmKf
AbihJa+zTWqm1zdDlV/D//2jl5/pIink3e75n1qLRKKtBf9ft0FRP8ZivNy/oGwY
pElOiEoBtW0iEI0ZhQRqKXgZhfaszKze3sBD/MgvYhiYjloLF9xA07J9SHs58Uhf
jgeKr3sUTYaQIWNyitiYVZV4aR9vVypobGcKaiALtm0VWdVq2opUX1yo22SoXIe4
9ftlgVf9F5nlB8/+9qsC8vat0sQdhYsk+z+JDZsT9mzLMLOr7+3T8jU/VcduhCN2
EfgSu+6O8yoxGL7KoQ+AQ+ODEf2FTwlSaCtrAZgxb5sg2HpeKyq3vuct8TpeMxww
08u+SygJGEMD62bZhsf8vPTOqO++Z+lbsXDFbNq30R1NgFpZoxmG5vUwRag9Wu4S
t9e+wKfdvIcOxmbrjIN0GrCy/zAm0/FQ7Ta5ya8v8d23dXhiLzKSZAccXUabRKV5
eeXVihC38/5+ihcAN8J1NXkkU7oGKiiYRk97MznZZ7HAaEW3lud9SP6iFSkcfxlx
WTzAB7hp5bE6Iy6b7ZJOOvNObGGHVg8kVLD8eQq4/mfgLka1qKGdobDUup99eJ23
wjJCBuvxNCJ5/WLG3hmFF54j4XhxOcG5D7UVnXu/fvL0rxq2wCyCADMu1OOcHYIV
KnY6RIYAOmgYcBfJcON+ufYQUyf+gFoVIZ2ClZEQFxolErbBRSNKvd4I3ERjTzQh
h9F9DcRGUTGjjICZEo6V1FVVqp90k8YSBVJV+JwEAug3GruM0MOsACmhsxj5Oiv0
fHIU0ie+JigeAASyBPr11QDxFWcsmxK8c8+Rac1xBwDw2FVHA/pJeVCim+xRgVOm
gsuiMvES7DDT1jMmPdVaukcRiZrp/vcmW2GIJD8oI+QV5Zsv128TjnIEFOhSKs0j
ZgeGizlfTh5ceBosgYm8vwtie2LkAPoyfhCDEo/9lvcm22JEpL9lgv6Xz4rYrkNR
36WDn8HBZ3CT0io+c7DPZJd+gTx5AwxM5MJ72CF+9IN/ObhxVCQ2wCGlEu5hEsTd
7OAacNx64QnOYtCVPp4/n/5GOEjQD1b3g+gTVBnPuUIJLYzgL1H5C6XZMK5m+ws6
Y59t3zL92LVK8RzMr+LB9u9TYf+ROVsdYXYesmXWMTVnl/ZiqKPqs8b3MYHrGeUK
iRncZeSF5LnKf4Pet+d3xCdc6UnAT/S2mx+YVyoERLiWdp//wyB05ffCOmCcQkO/
xhu6BkOvrJu/EhL+yiHopATzUQ7yT4K6FK4mdjjHWyPfp6VhDcV99nfM/Dgvg0C4
v9faa4pcMXE/8o3EnxwR2r99J1asr07iqsgQQJdJTnbkZRpVCvFv6hhIQ9zOrfN5
/EvD8MsKOjusb5JB44BaggOHmge2li/vKvOO7yoE9tAXRlDl5OXmCQbwxCbp9liK
+R+226e60+cqPqjZBdDnc4sPUkvju6OhcSpM+O43O+cLVbjpRWsiiILqOjztZOYW
R85XqtjW8Ozm4o5Ee/VitBznD7/DSUm1gQoQ/GZZtKdG6IdO1IEuAYMI6wfZdtO1
p/LPbYZ3eEeOx16FCQi0aqwjNbJ4ofqyxyMcqgrWs3XJ1qtW6o0S2cI7mOaXkmFA
2xGcgrUHJO8d4RyV3vXN8DtcefAHHBefIuz4A1EHUE9Ee+5k1sFmcML5bIVVcrSV
+j4kzp9v5Z8XhymPqfMXjcdHaGnY6+96/n9tXTB/qnM/BZ19scE8eclPci17rUYB
xcjJ6EKXp9++N45dzWdRJxs+JJ2VdulGAVbfTB2i0gxTo/mtFV4TrZX5JVLyTKUn
0UImf5vqdNkZoevHjobVLIyy7oKBJThnwykDBKa2v+PLaCoTV9kTW8xWRuHu5PjL
sLkN3qh5R/rBh/5KTnw3jA9Ll2x9MZBjFPgpp0ij0j0wlIb2QizdJC+ewllok5XP
/E35b1AVuE+B4YNbAs0hZSTzOfZckaP9KTfBAP3e8vjv/exoPNy8F8Gn9XtRjb9f
UOgVWSgsilpxc2RNnp28V57IAuKhvEtSAOr23wrSR/PcBmlLvfjhneSeyvUbi7II
3LHuP4T3lZwqMPWpfJYB8lqefmXxjGQLTc2MiFmLr9Q0PNJrdhmPu5k+K+R3oWrl
fdskIRIoexoMRoogDInYGP4qGb36MMMieml2/U4aYAUJXqrRKo5j1VLpOS4ZYW0K
Z+ZHsUju+PHQPOP1IDfPoZ7LcG4NfO1CRkLRgATjyIG9QNDQ+/CntVDvK5H5JmvL
vgI0zlTIG9J5aj8EJwx3UfNCFUjDKAM4oXN0kySRwr7q8Y/iH/Cz1LF0tK5b9oZB
5VrmrBdEXtM8qgREGIOusy0ZlNIjiv87utoOuUZ2p9QdDjyXaJRVNVUEaaYUDpfc
PhdkdvtLKL6/afgzgZMzLIXOoxxQSWuEqMCCK4ZCrtLqCl9ZJD5tC/OgSKdwHlqn
iBVnDmX1oNgU40Qwwk2WGi4rlZ6kxgNvvSmESqwwWfKnNyacrlk7DfxpUxS9u5Lq
8lBUQSHw0/cwIGJA7QGsbikH6m5u5xPg1bNveLRTzMoyjLZqr/zRcUzjF2KFv5j9
3AoXylzoRFy1pk8ZisGjY5+wjFNV+cYfZzwGmFsVVrGF8VoKxxPLXTO2213tCZfW
1YgXONVv80b65Jz3NuiRtmCNrnVYbAxuciJhHobRO1ynSH9hlHpapRmmqAWTWncg
sGmPckSVLaZBoOqFYq3hj+JcvdF5my/J7gV+jKslAnXulwe6NLPTKWHKyZc4CaUP
/9ilPKlkjt0YevDMo/2c7ubBHxfAZ/w0abG608AcA1qCD5cmPwaaN2tOtXuJblDP
3NnCRq+6UsQ34AiRiMwkuRwAuCPISovWz4CF2N3qc6/VXlHyF2mucBb02h47sRfG
QqYJe/m6Mjvq/PDR5/T/Oz7IeQ45NqzuXUTTvJqPqebGEK2klSk5Lr49n3EV1Ddw
XDnzHDw1oAU0z5/lw78ex2/TYG9reJ/pUBDje9I0ifOb9FZ5VcWTVYDMZbIW5bBP
r2nY+2exiz0OGKLE7Xhe9CvGankkS/JWrp028jI47A+rwZ2nKUsNRFMC2HxCwhJa
qwD3/eX7XkvS8gA8Lbwlhn/3Qa3o4onQ/9ElvM1zqPTeYB8gZzdgA7Ey0Xpkx9Wx
j894uf8u3/ufjjYF3E5Tfi0TCyRDrt2EDkgJFpupaYBn+h2ABNmanTEBmfAULYoD
hX/rwP70KLOEw6527M29U+3dxti3qgkt7IbzrB4ycc0pLCpi34z2D6wTXU3HOiUo
vkV92oEPkD9V09/C7DBUDWjensE8jh03FRIkdkI0smyo95X/s3pgj5Zf+5z3CTqA
tVS5aQEY9W1quJQTbTZJcJm/VaYKAiDHEc6ENt1Ka3sH6bvWlWnp4LF9Zxg9QKfr
ATeAGiRAKV/D8F6MMyN9rm/bl2lpOKCBUXt66Q9CMsZ9fQ/mFGXtfz0G/IGdnAQL
96+6wYVYLvDpyTRlze6r9wREAqb3I2HgfmrERPZ889I9w3TX347eCZjORht7AY8N
mmYzXw+HPD9FyrhUgyeDc3TVOCkTuFxjIB2bmC/nPL+wrEoP3+hav1Sqj9CNUVri
pIToDxaNsh+lLkd/LuqGCIAdorrvVzsLGAGe1vPMDzhAtQMN4UlrhWuseR+fS0V1
LJZRkAuK0D0mJGN9jTWqy0CM/w1Q96TvBHzZlxrwxYOuO3KrB6IcjUVhyFflC1N5
NYVGXpT42TYEFV8CDaRKXSK/xs40ntVEZxrXIIpNF0h6gTpRxCboZi6IfoSfV/La
KEHKgKOEQ4tTYGj39ql6V9tbK1T7wFCt7asQp/in4GhGV0ue5kyVSY2+AQFLXUpE
9qf2Qc7M3Id3MFy+bEnxM99MDVreQ1QznGfkv+Qw0RLfjF28mC0tvbDW7H6sJMts
SGZ1oaVFcQjU2EhoXfmPISnF5xye6x9QtncCHb3CVMWbVFOBpttPENNs0kN3Ttzw
l2cIK+cwlHrhUXezzP+54WG0pjYUdxDsF1Z4IL+Fz01tor+6kPFJwIHwlPOAx3BC
OpBV23Y5eF9QVGQQ1M6Q43UxOYZXMx9y0TIg195N9zxDqF3OKJB6EFSn2nbPEibh
PPgGlkIChdLcUuRtRCBXeIxC3jAD+QSDBsDrqQAVrErRbh5Ih1xpgWD2H1Ztdm+8
WcFbo9CgLz7mYUP2T1PZugs5zmZQnXSlbrarWWz8axbk0whjrBxQEXefbe9XgH1j
ydTwKe4mgc4a0C1YxctQipdR1O6ys2uIQ29JsPY/bSEeLkeAji4vghyqFK3zrZqU
C5Na1YP4G35vAgzLktyQPwCP6z1tShg0ShThoSAraYMA3S69rPMABTX+BEI+HLk0
MVVOmW+NeA6Cb9o/TjcUll9iycwXWMlZIXPLtoAPNBYRb2hHB2qGt1l9jKgKGGQl
5yYbgN6FpK6kIFmmgcFBs10tGLl7/QgGptWHPjsixVKDPhR/wcJ70pKB9yYyPLaA
nKNT/DsuXIKlQe+e+jUp039mxRq+AeeyDH53TU5xgOoq9BxjKL6vaOXj1Ed0vrJN
Bd2FQhUlCU9U8tmYmHXQ7/+uyYIhyQ81/iChSoIbwhD1WHptxSfzIfbFKHVPTzrf
kHrVC6HM1STxCR29DQYvBC8eyLTytV+YT9fjZ/pq/6r8Vs4runfptCYRA3p313lJ
RcvBwy4nIjjfY3bbZ1JS/xn8yq0mFviZSi+VY/WVNaM0GaeSNWBQASP5W4YJTxMr
frT80OHUkYbvkWiHqTQHes2MgFxJEtIGeiWItlUuw3XyM/8Xf/D3mQi4kTSjapbt
9DTowu1Y6ifZtpHX60A+aFn91HxSZKDwILVBLEFKNTXbal8WHM31H3RXIFoI+ZfQ
Pfj0Mbs10mJJjOcuzMq1E0sfqHlGwLI3YJynFiIL479hAdKjiHkSbx6Ksvfd5KoU
EBdJPVOlWxHi+uhXxOUGgxupNN+USsYRuJ0gl3Bw8NvEKR0A2x6E+spJAM1pSJWd
+d7IijTMrBF9j+sxiaSzqkAkvXlvEfmp+GnyDT4iKELzYca5Qau26Ss3aHnjIed7
DhxrbluX7UjwqnRHTsJtR4UCjEN5DeNKN36FaL827QXIhd2nElfrEkcu1awOBWvF
tcUj4+BX57xPwRY+RbCK0kLR121LElj5QiqtyJZaPeB/eT8/2+wh4OfIEzZc8LSi
HXhC5rLwSF+kaouSLW8pE3viYykeqXFxBhlPE15uYnFeTvPUyEMdiXKBrtWTIaqk
jznXZm8BLvTe9LJMe6dIMaOayZziBLQ2wTl9X9KTW5OGprU8uOel79NvwsC1G+bh
uuoaVBZQjafshudckzFFAxf0NWiPrw0MmKxHZhxxtuMXE2+5FWdmLz5zaVt7CklO
mcbYWZYuGBeAqFNdbArPVMtQ1ju1X+0m9Jo5llkPOiKJzd8CBtGsqz0REbi0X3HB
gSJFMORwsI6ViY7vuwM/FHnN5GHE3eE1DdDIVdWcyfUQx56oWudVa5mVLk/I2PGJ
APjzFVAOBgDcFs8jmBvoGOZ3qyO9AbK+wbiAj3b95gQROYNl8wpZCbQ8u3o72uwT
R2CdN4fYrzD1iAlqPcN1mFtWvBVtYJQp04xG++MEake7Yt687QAnAGdNuE0vkygh
JF0JNm4zo98sjmG9qw82QKpFcf74/EAWFWso3tl5Pi5Q7DgCsyoB3Gk6yGMy1xCm
WMQQ/FQaZF2zPAvJBIKBT2p5o4UqlquCZHlU7S1FqvXLKzKYeOPvRnrCxO80Z2QT
ywgBr5MTeyLumD7qP5fZT3/BPohKSHsyh4SnPOLJc+1026t+3T/SauMUduumiEy5
Vp66YFBjXo1QP6vJnbEsaGeRTbdIb2Sp6Gs/60OSUxxtDndnbRq5V/JXK13nyApZ
AeO5VSiV+h+BrCv8LQLM4hewLXzrQJYxJNtlPuLcqL31ek1BkhPwTuoq+vn52FkL
tM9UH3jKLJdkdmyaXX6nC5vi/NZ3LShO78jqe4LhwaP/M7BlheoV6ZgjCOLs5Pm0
AJiVSGRq2LKalwSzA8ujHnHFCL4U7A4F00PZ+e/sSgf26EGYOqqNcnbPeHMCg7Ya
6WZ8F6Z+xHy1+fy/8wemAGIgcm0s7iDegRTvSmyS55ivPy4NOQDsOqfy/6MytY//
GlReyH85lgIsJfjVe+onkh5J7jq1xHW66CKpvWDSEZhceOWN6fw0JZLiRfy0fEKc
XpYCMseeOorBJ782wLRkpqWc2BrXf3v99bvTLkuw2ALilxO5Fw2B/LmpdaLV/3R8
ozbn/JrF3+mturG4zTNH3FTEnhGvEogIJRexvkUlw7UE4gHQ6y2PuqECEpY2Xy68
HxV7cEOsyKBzXsYZzEsV65mu+NmHHXz65D3/FJQ68+wZzvwLBbbq6gW042GLtn3+
XJYCFfJtsjcadoMeJTm5+915gs+xm6eeA6Hux6qSVr0m73cybxpQOFwwhv3zH5TC
4oHqE8BKuZn/9ZfPmirIDw8aHzw6hFp4tnm8FoabdPEVEIKNXNsz4H3EI/ddtQr1
xncAtWmMoP15+QyJA2MGFlyWi8agCL75kpguOh7UVoUow1ry05jWGtxJgMrz3iZ1
KsaqZhsHA8awzfxaVUfstH7XDYuP3IguahlFBBnJ5VZ2mwbn0tnYkJmXUMVqM/aW
ipM+MGZuQu9KGeXBePaDZT/jg/FyO3vcgpY3xlFBmolVJQqVcEVJmpDG7CzVtGtd
oSaiuskeGRZ3qUt0GDoG5CY1+vruqKKDvG4WarEtYC9edvruywiKUjHuqzgNwwCF
5dIh+HyPkGt8kEImS+GY3mwXAguy4GciUPK6kLU+h+ywFOyDiksMewaIK65A0DVU
DyDkbxUPCzu4Puu1TpvBg1DgOIHSvmtOlXrzyDkBGLrLzY3eEBckgn2xiJHOQWI4
Va8EgfSkxiF0POitZ6zh8Op7vwLhXVM7jqw6b/Atz0rWYX157vxs7i7DxFgy/1tz
OzH+Q1CFEYH66mvpvKnIbOxjvNYkxDHCl4GwiARemU/2Te3J8Go1LmNWDng92tdu
f63mridX9ig+8naMs6AkS3iNdEoakHZZzjI7FReIrShO82oubuCpMcqfGg3O9Z0c
OjwzchvZKDqq86/Zf34lKiSR1P5wz3ZscGbn67uQhVdIT6UIDYuBY+T41+B8R3Cl
92Jg9amigDGkjfyc9UCppmqMmPfUUm6fEreMHBue+QRXZ5Rr8r4mGNz2iotry0fL
JPjYPCoJdZJKpuFpPPtTdm/1gwOp2Vk40ca4nNkVvQouw11JqbWPV8znQpauf6Ll
f3HtAfv58nbeRuwJoYRq+rHsxjR1ppBJY4/Rk09Srih4ETiAeCA/do+yvQcUkKYD
tM1y7ewrDoeoxHyrcibWXrq8qqAK06ejXON8nnRZdjIq9nk+Ua2joA6Hz92J8j9P
UHTui1/lsWrPPpSv7DJ5ILE8FBegEMZ1tcKYxBU2O1LexH176m1Ei4EDKGKUOro4
HC5XVuo0WwQmNGEjpX2to0sQaJhW+c0UoxAXY/Y09DsmFPh/UVrKCRHcdiDQHY4O
1teYFWzvUnJ4hEbuPLPt5q9pR2/2gkIVZl0mV0NYJzm+CgB9dB9Hg38ipN+REe7N
zebHiaqszOo4UhmrNmk1NjVdn1W8YU9pJ0whb19E3mq+RNVbP/xk069Eh40Qj55x
OORMXpUKrOaY3nsFMqIYCCnP21H1dNoGwW2PFJqUgtHIAIOx3O5t3XZ1jet/NM0K
vz0IV0674iMO0KvpG5Y2Z2fiSWI7NQ15kdaH38ffLR0Lwlkm6a+BnBJAqWwi6DB0
hBjJhmDhVnX9NADUNP2ioQpyIBWFdN2xK3ELue1pQx10gfhk0ILqr/oHSbXhtW/u
jj/jUtMssPPADPBYQoEMGdkH49eKeWEg5m1Cp8zagYndYa8uAh6B1itnLrCE/BYn
++u9dIakRTfGWoKvgXoULlMhqUe9t5vvk+VtadWLNQGIzkZiq1MFZWp0A3Ka7IN7
707DLW+mgg4lEJLX9kGmpCfeizuc2oxvA7PEofvWKVKAb4L+hMvhhVXwyjukbHD6
8HtBLMthF/Lt8pICam+GffOtUdvcEDbj8hnLMM0RWP6kV2fStC1ZrYOwd1XLKl8C
+cl/T1rHgAaUvTMa8imQ03L4jJRkNWofWSfgTZ1B3VwyTtCXObMc204ubWcqGJrI
Fn1csCPxmkNDst2bPtnYb/wXiArCI/bW49ntYsZFQJEQHLItVioOg2rJ7UlM3V6+
iqkF/6+KZritgUc7qBxH4kuMD6a2soL2okY4Nma6f5KP1zbPKMxZBPsK8IRO/L4J
AM3EH8B53eP7N8HlmWxHTPnoFcO6UBO0KZ4m1ApEvwZp2CWl8S2mVUz9271I2hmP
P/yt9mj52jLfcXAACLkdRWHxZfhtRoarOmMBX8EdjuviAw5KB3hSl7XzuTVdOGn6
KJrrBCw75higt5SLFF2oxZusJ7nWT4YVs94SGtzgDC37eh8QBnv2/FdUZjoXmJy7
4SAbsHcwSYrq8Y87s+5sj9hdvgX1lZ6KXWuARNuoi5xtK+plpABNQhKByA50iWca
BrDhDAtUGkt9RPJkUmBfqDAEo74w5mfUHzSfCKtbGvDf4YP3AG6S6Q2kpnBSB8FG
Wmu1xmTT6WCgqQpCyIyMFdrUNP5whfoLwbjtFE0DRL1xlz17aqu8INaf6HCtBPRy
dRiWkzN+puhuLwvEcAWZuFA4/q9d+/hM8565oAnLz0/RSsyeEGntz9Awxl1IJOgA
JJC0KSK18Qz/PrDKPLXLOYzoU8zPrajBFuLk96Z3RFnPMAuFfRxmwrBFhuwLFhUm
PTxu6dFmmS74BfC+Aexs0P0WljzyQqK1lMZUVQf3msTcAkvYY5ZviOjvkxbTXngw
QoI6WLzfN3DGqcWZsEezZjZ9IQaTg5pYmZHsj1RvD4qX+YY8yXF+UhDMOGA/ubMV
s5KCTcbkmb5DiiqTRkG+oKnHbXVZ1b4E912cLOWa0lN8QJbHNQ8DA39MwGpA7YB3
IRXOSFJVBvlA0RzBl+GsRXnyQFrAqkSvzaUwLasm72p5CeVzy1YA55GxRfeU1VZ1
CHq9aqe8oh23DVRzxtq3Z5OrYVYjeuWKpjTTrUhWbwBi8kkB6gtmncDH+yTpqn47
4GeM2Vk8OeJWxGFVJYgd8nucd4KBfj/yrCiRZbUmpw+3F8v4V0G5J+MRYcL9GRK/
gz8+V9uvVNHvp4eABlzwxmPnRwIOGvKBKD85SD67XRYqgSqZ5kIFNNwXF+sFbim1
RSJRN/jvHaB7x3m40BSGZt482lRWMaE4YrSpxrLXSZ/UG4ULC/fEYS6K0mRtFccj
Wy5Uf/qZmZimt+f259xzT2OddVaFqtdpEK7XcAFoxsP7Yc5v4ha+iBq5t4fZTmAm
W2t3IH/cTW2s0yTPiQntJhksZv8+u39N2RoB4yBgTUnQx+Y+fw6UTom94ucjGggr
xpqYt6O4VSoz2qX7SZzbs1qPlD2ogagPkU6Ug3wQ31kUavsQTy/wjukrZ5CUf89K
2KiKZU/Q0srbYJxFn6lx15WiWfXi+bAfPcjbKBowC7ui49XiAIvgWOdYf0MTbegk
B05oRz410MIFqjqaN2H96TPz2JCx51ROwsksjiHQr4ktglYZsVSjVcugsK741B3G
zhRAwmgXIkYMvAkCPo5T5ADGgSGP84CVHCwMjpl+u78KzAzfcxX6koF3UvkxQrEG
ZAnD7vnLeQcaeD+qPeHx8l8jRgEly1bgj790i/MuPrepH8KWMlxpSCH/LPBKYy8j
L49fLvdEXrsoIcstF0vOhcY1S4MLHYbqbKiK5lAF9TZfxebg85b0OdVb6XmX3fpf
CEAK3LClgja6qDyIUk4aNvzwyDIGbfTLNi5dGvzLwe4xzd7Qea6yFIkaSZRpwalQ
3WMtG6gwl0ozmXug9Iv2ih9nxeSjy+R+gutiZBm8yEFimBmZ0OH6mD1hi2SNkDo5
wQuulzcYFBU/6t5TIyaB8MOY4yDEITOByohnOGh+3wPdqZxPN6Bpl3bLJakm5jvw
eu8Y0MwdHwkp8CUANUFhFB3TlrA7am7lw4dyEhYSIUgXs/taXMMqyA0xA3i1BJfH
exeI4thcnWFcv1ZCW7jhEPcaXP7+n3vRtqMUP8IIGsI1/bpByhJyJzCIyqWmnfGQ
PBKmnUNWxfsXYAnbWrcSn9VipYDJV/wWpTuRPICEBEnO+4qjzdlxnJWbgFEuBaT0
yAPJH0PBDy9QsYVXmct9FifS5v7ksCzM/gFaZg66hYcKNpzC3QPOYJYRDHEYevgE
1leDfOeFWBokQObwkMxNWD+9rClEpUJpb9dKffUTzSg8CRJlz563CVi+8IGjXoBV
SnihAx8g26e9lri8F/SloX/bbqoFV+W/ahpUZBkfFR4mS4mbcqyCMkZyXHmsDUDS
B8ra2uVExompVmArh/rt+ymy8Iju3R+FhOuRFgR4/9N91RZ6zyGtWHIiUThULulL
QLWMapQlosBy+0RnUMA+yajM/8FvQJwn0XBNWSzH+ZoxFWle16bPQ37Qo9H+s/1r
IUN1DenlazsVODkwpOlH0iPc+Hr0I0sJVPL9ufkP11ICGHhwz0DasIdYrc+zTQ8k
g+Oszy+2WQNg/6rnRpN5VkW7KOW5E3RgAWJ6li6+CNCVk3VcMisgUoZkvW8KTr5m
UhZunUcGlsDUuCVwkwIYnDk/qkmxlOo2slphQkTWAX3gtAm3U6SphVk48VwAEFIV
ITnEKwL2vHWZobLlmuFDvckqxDoIG9/iYN8V3C+YYZc1bEq2LOAlSyPJZ/styjaS
CNl6IF0Tlb0G/EOb1PTINQung4FpxQF/flHMZGHFFA7EfYsgRhDhabwnfiFTARgK
s3Ez224e1aCpcMeNpRPD0reFVCd0ZLJiGar9HdlZdWYXVitCc1akH8rAPiyXmr+I
zvpFu+lgNzGFLlbr4VS7C1HBcIR+jPkanh1l+we8tezmI9qgZz/HbqVSJRT+xbB8
CqSMcUsGOayKB3jjxM+dwQA4NqKQbb2s/FbE/rew64E+eWw57WNPeAVp1bCtyrDn
pkgQzpbxsXri9v2MEBUahNN45Nf1psP/qZE/CwEJmqEkBIQ2f6NVgq1jVU/BA2sN
zCMOGPB6mpmL112oXRjwOOhWqiVIJWOVMV08caDcZhJnqvrnfY9BYMSb519C5gXZ
rICSu1sYaRgdYCGWIVuhZey9ZNOBFKsbD3oD7NSZrxRBucDpwfiEGJ307UYGrMWN
xfmqYf4pl4/zcA6OANhDU661gmXU2FUuHQC4lkssUaVDmY9uRugjUAszN3jZv9Oi
60j5BtsVdwkJK/a/DiSpoHzp7/HN5qndNGWrh2Dc32knEwOMi8dnY5Ufmk8SrHxH
0wEnIWtR03rGJCKTsiXr0Ud97uN8wNQyRMKInzCcE+jZjRHFTstRLunlVOj2gnpv
jZjdTepwCVin1FUSkvOwf87MqLcgu1xmp+sdMtbfK7SRDJL0mJa7KmrxrJF8E+Hi
vhQpnjDFFxaYHRSfQoBlyphwzr5CKMYhXFINTCG2eKH16XY2itGRdic3CaWvazzr
+H41Nx8mGNJbzVJ6TA2k6HTG6YnAfvV8G29kYWmptItb4CEJ/aZKYNXXuCF5wXul
n13ZiBNz94CaggL1xx9+CNMoWGrEoi/ulIY/+W7GYV8or8NiUK6vj6eRIltyQUsE
Y7RkGWIfcjKF3zcMAHF5sAPol5opA86sc6eKvE2dTZ1OzN/84hyAGOw78Tmu+u/J
XXEToJWrZipjxCiAwoFDBkPclXN9fZge3NS7NDMgpLJ/ZHwx4gETFeaQ+1CeddCL
FJ+TUCkW4rDnaen7uSKO1bzah9kNF73af45FqV7230SH+z/UdfkfQ8IPxOKrVu3j
mfroeJNPkHdkOjYeOgK5FoGg4Z7VYqK0n7b8LiUdVE91YZT9oot6820VXRjG2jC/
c8fr3mryqidg32u9D0zGvWrUvtw8AgJxiVyv5ww4Ta40pubBcCtA48qsxVSlaFxV
z0K4eJrtgAqZi3E7RjeAdC+DPEiSHiBeE31MkfOIoyVOuXAexRQb+RqyN79gtBkM
FEu8d0ti+6vjnEjE1Yu9dRamh4DdU7svpqbJqabRjnGmplcZCa/sIkpw6dbgU9P2
k5gwNMVJ4W10qCY48AI+lvrRgpd8Kn9o+TmeFAeYGm3y4n+gQG/x+aZyXUH9Pcgs
0Zkzkv3ZiuRQ3Idhj7XmxnKppz2tR+gQHd00FaR0Hora+AUI2/PrYA9WEEa0/9fv
IAMokKg8oEal5qysudX9nx6Hz9ppgKDMJg0lS9uNXhLAv+aA8pDoorTrO8NcVL7p
1WbM6YKX08ZjnvS82L6tCl/yRA6p8ah2+GLcnoPVsvv0nDISe1L5/E/e7CGKbwIf
prrN+WaXPb2RsXS+SsxLwPMKvelt2ov2pdejXTz3aHJhXntwPu9pXSYTzCDsIePs
C1aNtmPMwlnqQfMGxAjn70gyArGlegrz6cG9uPJ3d2FEe7YvlgP5AdwRWtD3tFOG
u66kuoTEdVDU4I8Yz9DddWiLRUpvZBBGQ3unYwdkgoeWXGlDOYaSW9GawC/+fzM/
EOzJMa7b6zYOOjLPKZE3gneWa1VhsQUOD8t3xSRMOlB6fdWY8j/WrYqjP8//kBS+
x7tTR9Nuk45WIN3Y7kAlvByU6nGNgSerV4UyVd45/c+qsVdKxMLWK082tzJzf7qk
99F7xtX3pGZKzybn5mgPQjbjzLbFJlkB/XkZbc6aiq/pFbS1N6mzst0p+ubIyF/o
PRQoHwZgGy4/enU/4rCTDOUnGKCkm6TOqJtiTm1fBaVzXnNHDoBms8vcKnwECKQJ
2RFfbAFrBOIqrRndVAxmNWMQ89HsyUPREdr9A14dgLscZpsZuavlo+nA2zh4YUy3
DnTZ97XIrTnxn6WBxY5ovRpDNnaSL8gTnN0UTSZrINFdsfqTgVFZjrwOYB7KVNSv
toYILXTIRQ5v8NJWDfFwIyvzPXvxA5H3JY4OHkdK8wlLXjBAd0dspWmV6OEHZtlM
nC0wN8URCdIsHl3Faz4Wb6+koQ4BIPw+Olbj2PyfxzQL5Qn0884VZPRYSydS4MnM
DIJ6YO3P4nKEOHJCZBld+fx4G1C/7rhEZaUguDgnFLEpXE32XXWEr0X6bqq0JjM1
dDc8YU3Nd1Byj8b4RhpFg+N7o+LxLlAC5F02YT/Wd/ywzsyAwL6AG4yluHPzTMyI
OhLLmXTIESNM842T+dwtRPy9oQZj0KOLbYUT7wQOEeWajOICaMzvkj/zlGp00s9v
XaD4pn2dszY98mLu+XCSBAcxsfa82L52IeCk7F+vxdYs+OG9DCf5+sm6Gp7nxlgL
VVyKJMfPEMs5w1qM2ZMzJUPWuqIGq63nrA2hXKaxwB6ibKWn4RMJhMF8Sm0wMdHv
X/aUyPQGbFyzGRcqH+gdzV6Ub44ZqRx81YWTVkyWAcstz/j56/mersnfTiZJP5d2
RSYLrFpKmipjTSZUwJknyXPapJ2zAQjEu/A2vZa9Gd2ONZ0DsoI++1Fv5mbCdI1F
8IvPYLU6DUth0/ngehsL2AMWSvwOFdO+X4EP1HiT+VonRoG08h/h92y1VVkOJMvh
Ti/wH7EHZVCHDHe0v1aAybqlyCTGWdr8Ph0gjqeEbXMr6qq7UXOLRKhBcIvMrRjj
vo0yPyar9DC3oGy2Z6Ar2SWFVTZU9PM6aO66fiowV5buIc+WSFVUYfuyGwhjzU8B
mr7DBpb3ayaT+1rZGrx+W6e7pagla1EP5Gkjm7xXiKmjWY/6yCBzCfqpSl/csltQ
rpUjM0vUVQrpl9yrluye0PeC9yAreoo9ZEfNxMo8GT8USoGeWQfSSurAhyiuXuTm
JD7XhmQooe6dYFs/KOgrv/YjBFQtrPkm3nbc1iz7YVypn8RxgQBUIiL+b9q7r1+7
pxACEx0xY8s6NmsXkfaLLkj7Q55JaS4ArKouURO50EIN1q3ay77H1EqUCsN1Criu
wTL0BIp8Y34n95jqsQ1hkfU4EKlWbGoPYe51Ji8Rq0ZkQnZnBIGctS1y5l/FFyIX
ah6ZX93+j8kZT8GuRaBiv+Xx2yiqbdYMg9a73+v2OiuTb5BU18ZWWFDCB+yiFscn
LMfHx9dEtLE17yZQ7Tgt58bO8uVTWz4LOMWzXEwxey2o7Jtu3ad0rA8Jee/hFIwE
7PdczNcBR5EKKIpv9qGJwCLr4lLquZ1TyvLj5W9K8zypQJJuAgKgGGwvE+ydi3+q
Gb4L+3lnmn6PV50XJhAtEa/UoQestNCODYiSWCRi4NDKO1WWfMGJk+N0wcud8F6s
+Zy06zfVOFwGYp9syhwKuW04Ure8I4+ctUs111hV3RHG7D0H3EhnT+i4WCkLvdqk
9C9LEZ/DCo0+zbC/I8PziWDB5iougsSKleUaktaa2J6BphvurXBoKN26CVwnIm1o
N6TYhnIAzBUGp7fLYBhFbfgddFg2kT1F9rh324PGBAmz8DsqaG2/Vr7g3x6kDC8r
IidejrRYouQ/Vy2VVl+wM8yWL7lC0VULS/5KA30xDnFaa0uT7AMCCxeAdfBNzx0/
pe6o7b1W7hTmmkGV4MD0TlVMGSpW8C/7Psp5D1C2/v0oNaiX+pkSCydmeDRDe9R2
rX0oxaCM23fyPNE2qagVS9mOI6VEaeoCFSzUtjD4cV2sM7jcELnrUkV44sJkOj9n
0210SFxCLNiAbifcL90sZMr2xUnSlRgHIUpGaFst6cyeX2CqvidimUbffhVkqeCs
XSt4KWSuEwN0cawd50UnW/oDlvuqN9oWQyOVrJ6LjPtzgFsHA1URiWbDGky1zG7G
AyFNkBABJruAExar6gxZ1HpeyAvg38d5GwB54+ib4ODccjWU70snCMrwklZTzIkE
rH6mZvoiCnvEjdp2jCMhscpeN9WCLLwv0m/SaUVB06xQeyupn3Fy/NrkLFq9SycN
hzWhPNZp5FOQ4lkslkyBdxvGzLBjIJjCs59g+qKfPcg/CaP68u2Heh8+h7aASdNR
zTqB21CLyxu8oEOPy78EQ+PLG612B3TreuwuDMIAPCVYfs67sF1zG0/KCPG6Qr8v
+hHKdKHzL/yS0ctEHZqkapMh9w6I0cLwoTb2jxQRVFaLAM7o1+R8KCfjSWVab3dA
acdINgbVtPgrZa1k4687v8K89bMycJ8JcyTb4R7YE8sRgQA/WZ1Jra73e1L8SsFx
RmWAZYTkLeRxqoZBhmAceQmVEtjVkqp0gONF4DkW+pnKgD06Tqoz+lOw/ogP7KpU
kVv7tPOl7T5ZJ7gG49Ju6kvoRO/hz5SJZu+MSkMjEMfDW7DrA1KEhk5YRj7VCv0x
9+r2/sM+gaC5BmPEXIC+5D2TE5GQy0lAGODUobB9/6sQpNBkm9rXGG7dBVZuKMVD
V+fA0FxcHOcHN01vgWnQL6aQjt8Y7eeeQhCbpUMt9UaBBVwveePaUHWR0NBAcUvY
UI+QVGRpBxsfgxVRnowiBYg+s2sfQefP2zQ+5TCNCuIrq/2bqoH5yhFupwESqbi+
H3vkDSSOPAp+WvTaPZe7HtF/y9trTQASbk3UoZ3Jl4ccNVl1+3qP3N9lJmgk5aJs
FIZpc4idT6NG3SrT8ibhrYvI5LrsETX9d3lxPutds67CoKZu1DGdKUPOCJ/YSovq
8+/czl8HaagX4+7OEhN3jUrLXcRStKGJXvMXtWUe7TGPVeJVExmIdRQIzGao+tNA
12mTHi5hkiEYUnPrtNZc/sAH5HqNMFf8KOtXHHFQe27/7X7ezmY4nWeoVixDD6jI
kDxPHybWquhAzYmCPuEQakLC9HnNt21RzDFTSQiCl+xxZ0Cp7OFIiB1Xn3FunSS3
nJ+DRfQf0C4D4MWf6CHdrIbAY1fTOwROKzVZQNHRuH7bpmVcvsb6PKlpukCS6qgm
lc72B14Ph73WnP1IiByACOgaSyJI34Dp6rFJcrhRDYKG0eDod1FeZAI3Fxl0czZU
ru8OhROKt6ZcyTO7cUwShFEQgieRthFR1GZ+ydNfLmaoQZUso/Kqrg6EoDEZbQ8T
UaonxEZU9y3NuiyZkF0SgwcTs4x1ANxSIf9EuLjRWIa6CU9+sBeDa+PEp6sOzVQF
le8r27DvaGKByLGLZwsVj/679rj9BgxliqFut0pPCZUcAv8W8gUvxshe2SVv4S5Z
fSYMValOiS4/Ym8VtrADdon9GmVUNTO9/DZnBeXjZtpyb387e5ewTZ294fi6FqZ7
lXsA5Ybr5f1pHlCvMZ5OrA3EP9ofjAP3tcZxfGBwKMe8pFm2WbXJvUOjs4XLxRYI
Ljv5NJljOUda3KTgjywtLyypo17uX2KTVQhU7/rvBboUHEfFnJk490FouL3cLG3u
JoskSsCoaCtxzVHQBzPsU9dJvkvEDIU+1botA8B6p2AxBMPbHXtexTTXGs3tY8NJ
ip2C7SU9QWCf6zKVHG91rXWs4qYnfF88cJLamYS1jjII4pIzFdr3yn1tpSO6aqou
0l8qPPzfMAyqCMfTZSBSTP7dC6IflClQzg+AM+sXEU4jixbrcxY5sKxIMMzmnRxg
vELpQoyyvw3FoiI4B71iVA8+64kKs98fEuRE+bkJu5Ga7UfyT4LMvCMAp0Ub05GP
k7Ixm+RqY0M0vUz3qLfAlL0sQMcb+yqZBmIJRCPBiAU27DTWT4kDQeTIc/1bVa0Z
Kq+6Jc5KSM61ycT+C2UWReAzKYxYV6FTF+oC/l3KERUSH6XZU5ZSCmKgzJO27QGJ
JD5ySCSQorOnuEwbraRdp3BRP7KEPYRrGlymk+woageZZyZeca1KBPujzZvUEFpM
U89fp4JTd1jetnpy9d17L9ERdHscHe+JHlyj+7AKUA0gTdHDsR3/CGpChLlkNWlJ
ZrIAR0ERw/sTEER7m8fUU5TDdg4sWy1gI3ytdF8w+Yz/UC+A/A3CnOlKhQKDrh0T
r7G7AlahurNbfuUJvltfeU82gp0yxBR0oWK1guJ5GPPHPvqYIHq0oRpO/2FMGxnV
v8dVxn/bkfUPt0YBWtu6GPXXY1xg1FdrGnf7ENCCTV4scdEtKjyVE/F2FQ+KIqdm
p7vy28vypv8XY8ctptTSQkJ2K9QM3W3sdWqHOjv6VCLCLdDkso5NlQ2eM688wfrM
Q6qB0lN7l0S3LHHszfkkXRWe/5nFxRKQWWK5ic8GUQK4oMA4N2vGA6JFQu/vsa8r
nJ0Yo8Cs5ILWkK0fmrqBRzlSNI3mfhcMXdOK0JPA1TTQfijyeNgpcDQqeZm1gXI7
Oc0R+Acw5ZcCpSES9nXU+AVCdchqLf2M17RrzFUagkhkfD3R3RQy79j6IuvyP2iq
e8MJVnp1ad9r1ugN25+Zg4ZdQD185AsaKMTnfYH0recQw/95g532VA/1a7cq0EBP
sHjnjCawupplUM3mcX41M998IuX5NRY8x2lt+6DuKEO6rST72RkqcbAt2wCOPSzd
vpmF//ieZOuF62SJ9wj1LFDFmSxWNQy0oMGZ5W+m8cSVNIotw7585GlnIc7tzuZx
2uWNlWsgc9vUUwZI0VIwbnwxDZepYJB0BoJt+c+MAEsoT/tsJKrN8O1YHWeieMuk
m3w+1SsnM2+R+S/1GiJNY9dvKH0qxkK4MG9OnUZTL3M+1sjyeZZ4hXF29x2lCla9
3sF9Cb++c6HaKZX2x8r0/R7yqpKdE1T73LBHXQEAzVLVT75yqQD5KpsE7TYjCvel
Jn2pK36oiS5znA5XQD+1ww/fWEbnmN2DyGU/lMGBExQrukJMO8Vb5RbSvh0KqE/7
quhuuZsyQ7X6NTQSBeqXwBaqbQozzJdl31vkw8YP/93kcnDz7t9jbgTLIkkt9Y3b
UMS42ahaKxGO29ShjCpRtQMkrC5KA+lBbJs86vMg/iPZwrxswkCZWiaxf/Iiw2PF
/Yu6JEDEe2h75xn/bPj0ttH9wY1yjZj237538JL2o2Zg+30s5CJLwRAh5zeLvvUp
UeIDE6h5DWlhius15xiSh61xyij3Fg/i1NQG3a8f7vrFDfCEftwI+Fct2KHRLprP
hn7e9ga5x35FO8/j2/F40BZv/iYsV8PtJtHehoK8RPNLUzBZObC2UtR8hR+BuYO3
Xp0c7VUICw0RgOuusd6EGqQ6zOfumI3BIO6L1GSr9AhlpsYTFB97MnyKv8XlMTgr
G5pHWrLEpypz43yjCKd7daoLDv/9/+J3i4OhvrANQh6u+NwTyL7B36MCK+1Ajmil
WeoU1hC9v+nzp4F1tk5DDbMhu69u4AVSfqKJx6b6mt6jNheq+MS7u62WkzeWQ0FV
p+9XLKKmhxpiJmpoiiI9Rm1k2JHOX83iPa1yuHbiaPMMPtd8Aum/kmrzPv4d85pu
CDXtd8Si0FpR4SHJEQKNDTbdAiM5lOAk/2Q46QbjlK1OWxS3LXrqhGM2P4oHYByn
gZyEaoY+hZeTXuiTYsZy4oWitvsxZV7sLFTPyo/q7JBVbYVS2iGI2KCUt7F9D9LG
1pvVgaj9msyimPXV1lqbL5vdOPssDA6RHNnTwGecMBxZBsveLFzPJxHTUDMxJUrR
NAn013i91N0MS+z4nmSuWKNeXYVJAAhIFNIkBeBpS7rBVUavwEgnCud3hNrT2wUg
OmCxhhpw0l4VIlTAcOmw60rh4dWoseX1DJz06rw0fgiNo2IRVluGUaiZCZ/hU6cB
nbL0wD1KJzPQvTWgddRCIDHH3gcuJLZhoE5P+PjpeYDjh16uRSZVMvnddp1nX7Ng
TuiL0LAhDzifeuxxTZptNtqTCAuchJ+IjFwm20u0yfGx03Xnhmogog0oJsKlJHmR
H91W0rV1VSpk6vUCHxYn9G7BcezyofU92IliXAkLDzfynPF7leBtlclZ3QgNzKmm
ixrDUtuMAjE7IsxP0Tqe3B09qkyjfoZ1lNRuDp4B1ExHd9wCorsg/46bRgmxdsaY
4xRIiCofaequ8Tl5Zv1ctMhUaQG5psqcZlC6n63rEGyZTlIJ+U+0DCU4brxDNEfp
8gnSwJudV8IPw9RsQnhPAw5SjHMifshNl3JWwmwrSdInxLP8npRIUvGjt88JZTFM
9PPMlFJ6viEZt4EjNqYfIr0bvRl1oSC1n8h31KOSctC4kS4QdpvBbN0AQJovb+zT
Wu/eVWg5uM9vHdCJmpgiBtaMlXrqjVCqgL8pySgInkzfCL4t2ytdKdvM0J73VtDH
/MOd1U3HpWddrxrEso94SdxWajAVKhqPBfCIzUZwSCmW6AxWppxITEOQKcAQ7L73
U08UuLSlWKvS7KxuAFpFm8fWkvS8h+nUjTXJE8JyHVNg2tlGuPW+0YWaq1ZkdYnq
vKAoMjl+9+F5Vj8ilwhoDGOAekr7ORs7aKsSaYv96uR36mKprAsStrXGjLAwbHn8
dnqQNkBrH1AT0La/fICcDkW/U9OgxQ9T35uRU+kIGsaT221DYfAXNI3gcnympXGz
EIW9wnWLi8hxaimsZYhXHW/dgrV3rV+Y+ftCOI7ig0fr/NktAyspmHL/Fyy7KT6p
lBRKzJ3OO0GpA1DooPUAHB1BkYqUdfvIU5YcAApQHzB8sSPjGA1x5Hs/NmzO+Ywd
atozlTB+izbgnl8KxBr2lxR2R5bWvL26euVI+sXrmaQMgguwHp4x6ch8EtFBY8ul
vEspaF1jZxTL5XY+Ozr0XRm646qM0R77+mx0qff63mt9kT0uqVF79ykrxytLsccd
SM8KJyqH9vYRI7u8eXj5BCxWZXMS3m45ap76K9PA4HKEpnLzH4nA2sBUevdNxtqJ
kWxh94hm/L4GBSYYQH3LoNFNNtxfpyUCjF2I7WCP+OpGEf6WL3tzpCHlubLC0gvJ
UkDaUfBhkkzg3T0RQX9bH0r7cCo3pSACEnwBKhiVplmenkMkGd1si8OmSiTzU5p8
VVRdMTNeZT6UsRYhco6AAj/tyZXP1exdGEi2+BQeOy5GFLCHrLeHJVS3xQzY2M6p
98qs+0pw0O25UGmrxx4cFSsyUiW3F1/j16rXmL/WuGsVRQ7yll1J2J9slRLTHFxf
vUoo5jLUxdtJyPx2/lsPHFBPPTaCnmwZmJRCbXRUsZiIK1E00OhFG9v8raQHdard
Xj/RjID9UeHjt7Uto7FiELf8qtAlrfzFMwsVYeJ5lmP8wJCZjvUlVs4OWU+5c5Eq
evdwLXNSCDtMmbhig6jAPK1qCs0bph9MOYEgANmq/E0OxZ/wJv3us+f8ifS8EBsj
kZ2LNUXaao7NCmrYZAu8Rx7umSmixegqsxiQDB+FVzViuaYT0i5h7e54+RG0QeJ7
DhV1/Pug3jCPLkgJwtfZmlhDuNcJQNJfXC+4UDM7IgiimhEWDFyc3kjqB1aPnFJ0
qw89dD3zN828XQOQQBlKsMewsKXBGgBD3lcU9a8XQL4Jz/FB1L8Jqc/lckaPS8w0
/Rbf0EmWF2L9iaDkBXCIlIycYNn+ts+6BzpsYMpXxhoU+OytYyWIF8h6Iqh8zxth
h26UjOPCIQBbSHnqN5bML8P6ptiH33nxE29vhH3JUgK1CccII7zVUhBUV6VabsUs
EngPL7iKtWeXxnA29qmlu4BYPP/nyzOYRS9mMQAYPlQ9Hc4rONzMkt9MQaXufQcP
B0+71goUW8xwIx+Fj59sv4OKbEMS9d8+Ni9PX94hMVu/hYnuJiKCEKTKe+FJYQ6E
bjRqLsqa1pSgA7SU6BpEh9ekNZOTdxZrk+9NfXw1orFRnhog5R1INY9zVcb54HJe
PKUUqvUGzfvjAT+fMeWOle6qOFHxwQBWDGMkRmWPmSwK9FtllXTmK7toPYj99cg4
bUElWDbHnzzqWqoFtXskaAL8YuOnDcwpZqzLNo7AzCTMx0TXSilEm2Y+rl0eFPjE
F4fvL1WFf8JUCgkl3ipMTLEIfz5tnS4QAd5Lu/8+BwrfrLMob4rkuOjZVADYMEfK
YCr0SuAZBEa0CDdm87s9wUVUdX/UMdY84d0AGyS7fva88cOsVPdLfvDOKOq8KwFG
LaajhkotDlUJlTwKdJRDLuR/+dYb7yjnGruwqhKdNGZW17zAjOOTZkU3zNQfjPV9
lrpk+Y1JTzp8wS8+ROo9v0la9sSXqFqojssNS/c5und0mK/B/8Ce10GH4nACbsO9
r5wzP4zQUWiN+vr/Ev4g4LeHGtuUGPKib+pZi15kQhAqZ1DA728TdGt++bglQ1Tg
Yelv1ipLIhjwZDLiNbtXrgmeX/Xlxy3ZZQdbh97rw7kryeVt1JNSiU6qPrzqgx92
fT99YKKxPoCu0PWQacoYqgujlypIUBLEwtOxd51wk+iYMAXh6vgBit1AxYC3ILED
gOWrFPYoRl+yVZ0TTwbA3kXLUWf1nS/D31jnR4I4Tz82LqrZZm8V+Y/R/VXnQHwC
8Y8kvcqPiq+6rOg8BS9g0zTJ4uugEMnktV/8FLp+hUfQ40/h+jzFZnetSs9tDd4s
KtDi7AVxhU51XftWKJuZLEYbtWrh2l3tl5jnNEGuHSEzbjRBXvkwxy3615HZSAGi
Wgw8N4eip8p/iF6PllLAK/LjCBu/hVy5/sqYG3hPmF3WZJiv1Oi5ksnfSX40QI8e
OK0fZMFWWBARSbsfn2qrf2KGudkauGrT1tIrOopJcBdkznV5Lq5wbezAhj/71YKF
rj6v/DFzI59a0A6aSd5zTJLuxROiAuJB8SIxNYK2tsl9abA1vWsbxoNwmrugf281
Rv3YnJ8Ta2rrvsAxYD+k4gQZK3m1zUtWsQi2pvBKnxsvfYOD0MEngInpaWhtLO3A
4QCJhh0Suz47qx1JaQVWCstHNChkvpe65XSUiVf0fKfg9TnTue/AaijdferG+GHM
I/zq4Gzntl5yhJbZz/UCCnXhluqRAe/66sPzx+YvsaHvvYxsqHLR2d8wPhG4jiLq
DnDoz8Lm/PzBTyc3MgvH4mlzB7GKYEFYgN7QqHVBRvgo/HL9xcDlopCWNtsZHHk0
HpV3/5ttH+wT1B9v9OJHfb8gQU+l3FNLVpkHBH2r8meREMztVWXhVIS+dTcD8yld
PXrQWvZ5FHJHDkPNW7G0huMKdjGVyRSIfYM6SEkohoOBnc2Xm85eAiEbQ9k08yxA
R431YnlG61lJi/TXPWJtxIAo+W9M6Mlh/KpFg4hXZw2w02fBWXJT+iOuzUMQhguz
8/noL1G+1OAwS1BoQ4I7G5rqDlcf7ojqzqprVLGgN+FKZWqOFnxHpgji8Xrsn7Ie
aT/UoefcsmLGweoXk+mYslKMLPObWaq+V/ozVTX/gPneINZ57z3xkoJuX8p+7/vh
ZmJw/dzkrQZAa7gcVbb9QCl9jLsI37PJ0ES7jsfoCkIXpoH1nBRXayWs1M4WAB+C
VV4o9ZA8DUqx0fkTPCZS2XfncxVqKyX7RLz5K75GC/o43ouyjEu9D3zedzXQO+J7
BIcHPc+XBbT0AbVHMwyqMqZdVNMfyl4Qv+pZHsXTqEug33Ma0guytklcnweQnyfl
RWDtRMKpfP0KttBiJo0JnvtB2B6O0KA7pPvsgvARNZpGCOVBEezlOx60/uysSUn3
GE+MH9Esq6AAR/vNzUYfFxCPycsMjy2Gl2UhoonWfOwSU+rA0M6sUoYPhsT3simi
e4CbmI4pztBBPRC3r9eTD4nJ8jQXlBYjaneRZnIM/B42ettI866PIh+rTZA7RfSJ
L7PhNNashtjaDd9ADPpcjTPq/qKL3Kk2hZdOWbK1BThsqHmK7PP71Dw17f9vuHgg
p1Pa6us+Sf5oJFizwGjWgnca9yUw3BeETQv3XnYzjaC64lI1YlWlTKw95NPIVUed
hWGf5BS0y0ALcJlnIzgmhcPsR5gUJp9PWNok6ZPuwuKig8NlWDwXYEnlWeN8bF9P
AUS3qiPrJvvdGKbBcFPGVhSkTE1YROhsOdOBlzDKMakuDFn5WsTe7b9tQfL3hIZN
Y3EDYPJbzvnK1dZlEHlTPM5LOUn9Fgylqd51mw6etwHWMhPOcUxkto7s+qGFPzYe
17nBhy2Js2tM0pvkTBh2yQCpgHYHSqvCE9cFSwDDK3azJ6xvCMg6hj06hKTJxwdB
9CpyzNj9VQ+XRbayU3WPC4nOi4oD9GlSnDKk3ibL5ZEXbcY/LyDg+ZT6Yn8/V8T/
gQvM3LA64BPqWFy8ZR9apXp+XUjPm/emCT1hVceV8jMcKxVLLyHegcZw/ZI3Vrfd
/TDzSw3+rML4tzrfSYGfBVnTn1cyRwz1TymhCeM5Js5Icm6SR+T4rFFGzpFBIU6u
pvDTa8bcpnuYPS0TmyUu4AgIfeQgO3rby7G6EUPuVqniE37jFKB3E+fNvdUmKhLy
MQFFFIaNGzCOuxp+jyksKcu+GIdympVP628SnZSMYbWovYbl0zUMnoucLL06KpxO
t/r3UJsjZG6efTpEh2FuVsCoGSjWPRr/U34abkMPDVCao1nLRCdBrruNz1+Z/mTI
GN2ubZkfbKtCWeF/FMUq757jsbe108/qkDTAs25tGLn+MlZ7MF4v3/Ix5iQsO0/9
hvliAorsQxcVllRIvcxqIf/F4xMcruq+yY0HCWkXiMWmI0uijwIV0kVB5iFD5jEi
MuhEakjgTp2XwlpbtcjWj3yAUtVJi1x+o7J08lJs+26lu+Hu8xbt3rdG//T5A4Ic
q+AiGlTi4pCck2g6D9D7Hpqv5dE2PcV7jp0uOL9THLV5Bks+sKpj3q0R1BEyjMwV
eloX5jmDoDCd7HsTX5alLLNEb2BbOb9t8uDDswX2Q5liOaWSQQa3+6UOxR/LXoPe
3DnxG2WIdJNjnDrGy5eIshY6I5KTA5Phzx/IK1QFh/3AaY7W6s4lWyTmCDZEa1dN
XizFMhwmrNR3HUuhPIX2In733tg2QUkERqeCfXt3G3mHS9UWZEZCaeEkqJP7ElYa
81X0ezhGIgy/s+cpOdh2jy9woQwosB4gXAy1BJDdTHDOBk3DI7axFNGT44SmLOPG
FG4sfYOV/oI8WC9UYxAKii/UmqeGjCpKOkz+geCGtHY68AJ/i+8sTx2IAp4BXUDw
wXBj8cGJkdrue6xXWhCIhmlJ/jToQNw3mNVs4qGnj8RaVPGtxsVeArU1pcEyrvDF
7Zla9qa4iv3lxF1M+I0M812N40EtzXE1djdVl05E5yl9PvT+OZyVIaoFsNzZEaQt
9VsG2PruLeWwbDXNHKXFr2+aacNB5WrRNYl7hfs4xu0UOTWgCn7pr0WAjS7DXate
rMHTJ0xSzrH47+8WQc4fbQMDOfV6IBxNsfQ5DHcBBOoQ8Jz02oD56kM9bNSUplvz
n1Jy0olqvkK7aXYBJXvQGq1R6bFG8XEpScrLp8V8bABzOotRjziARsHbRzkYF6KD
sS8BumbkIOu4YDGLLVldHvfc8PJQbji8Dh7cviJ8VJ6wkLp7PqFp4gYZLnJV6RKA
LYpzju70y2A6bYZ8dXDYtOT3+FhAKg1UhGr7ZpkFKSskdDmFndeeHnd8/tw59JmT
VgFaSqdpHyMZosuqh/0xG/MO50ATUq+zgHyRUW/naNCbm3OQB42qOIozj2kRzwlg
7TPuBhj5//7MkitmovOcpa7NhasFDzmHV3IFr+1Wli0p28Wc0apYZN8I49hsZcUt
0PqpSSp5qmYGNv9ZG5phFxHj03yA5i0p//h6AVHnAR9VXpUWUR2ARkG5SZX0bm3j
plIHLtd6dXXFk1O459nfED5wLZx1oyCvtllROpNAk+cxKkvYoS3r7SZG19X3WGHH
pqHgly2NJ8raWR3hE037nbDWHXJ7GBedWMQuDR/DzrZBC+rVtRanuWQ23FRfv0NK
poTpmscmNeCbVWV6BrEoka3n6hPEqxBYBUaGe6tNgMIcII89RawNvQITn7m+Qx5Y
j+qrBHk0qnA7Frcdo4XHF3RrQxpaQW6b6OHZkML/rkdLXuxmHxgmaoCwpuFiP1L6
4Jy4rrbb4kBTU++Od2utV1rWBCY1GE4/XvOcUNobBf4f8R0VG5IPfFqEcchlUwR2
DHTMZCYkOhs6O6rDTrCxZlgrJHNlnN0UhAQNGasCS6CP8wDqJx7VOtq+ODHVUfnS
rFUyhA4Qr46QQnbMUF0LkXznQf3+x+ID5Co52XU754W6cW6zcVB5sOZmzMtC+Dbp
YH1+l64gJCB1vNgfwvW45nDh9ZiJzYMHZwdM8onsdl6rqz0zJIiu9KUCd9Fv2nB7
0F1PsyPb5uIH2yJRjVUg5HYJP1RqMGe31Aq/5ykCzZjTbwIoisDxsJ30Sf7K6etO
W03bBPeWcSUZGdMhWFsI0EG/s8EXkjKX7ETKpX21GgL193fU9kPAI+VGSEbThnCL
0tFRnZjqQbBMiBoEPKzex5YRyaAe/ZJbcRIE6boX+eoJLwSnG8OCpZz/9GyHI7WX
9BY2yBvqNDluxMpnYP8Wu4Aqi1q5m74BF2U5sEdvMPPW2EDWV+eC7hj1SH67gO8n
TK6wDuQUFMZAhZ0+ccGJ6ZB6+p6+LtaQ2m6FIXciuUznP7Uli45uSM6a8mBbq9d1
HcI1WZo9dCD1BIzz6K1WmBdXc62KQtKolsPDioaGeaTjh30EApY/+6eWvG3DvS6y
+hjMZpiv7KE8yI0wa5K91s54tylXD0tPQ6mjVGeKKq4O+alFh/aLYt+Q2NHZVny4
xq66hCO8ky8vOmnV5rMjqlzmg+wpoX/AlYQSVMi4vdMplIFL2b1A+hg/m16FbrMC
4bWO2EvmQuqUGdmQp5rOPipkdOl0vyouDeTwZxqlGv/pF/EbxJgElHOvify42QN+
2T9JuUn0pdJ2LgfqJFCCsHRASDUqJWg81l4Z9E7vEg5z7a9SHIHcTLn3JDFY9iDE
7e1NMxw7+8kPA4lLFiXl5ibrwDyLeWNvw9XjdnUBZUvBrRqstbh3ZsJqp4yJS+Ua
m/Pmavk0Q0+eUuGAkyprH7kX1VqxRLaJxC21pwbcSf2rxI0Zac5yr6Li9prTCxWq
7rI3cgDf1QrEljC8BXkv0TEwSAEFc1WpGgIDZbXkQOlQAlQuLwd7fNQIWURiqkN5
KWA/Vd61Dliu/5Fx+hImLHFuNl6khIK/cby5OtVLWRAlv3Z1+kiNi52E9XCybX8O
2IkglGdD0i4SeWDWwxYJ55fihxDmkPrO4fBk0djI+mZASXaPZ6/c41sTD3G26LNX
7P4G2VyEERyjiD2J/mRwqbc4Ad7ePO9AVlfSdBqJDQbtYfYVETLOH5vQyz09j5j+
yq3abs9CM3Dt2AXWB1y/zaZXKcO2RsZyyTwFVK9aaB6hEVxjuQOKpt68Mfi4TtTF
pFWL5sX5uIEi7MUowJAzfX1NjKBsL/OnZHND/YL37eMzq6/38/khLtKahuFHRUm6
4VrX5riHagXUj0FlfcBYb3fISygfOLUQr/cASjkZStvMHDz/n1ClNNpoNXvxr4vP
y+zUwr71TUo75+9SxxpVQMljbJknPhGEo/TNG8oCf2/ZXKqwNwkVpLzyWTCOVmbG
/tYspYZflXXGTd8//kJIlfMtvqSkQYsoxXmMqwLwIRU1DdI7Ncf0UTWLORXXODVb
WJgvgUSDtnohepmP5r0xOHCaX49ry9TGryGGvaHyiUazjHVP6w5P0Tvk3XD4hixC
OmHeHd4C0113JU0ZpYFSB6P98V6GB0CJ0X4LWyHqk1toHIKOkMtSuTWibpHCf0Sa
3VMvKa926ZfcuIVQFBt6oKtmVBo9Yu4+FdayDLgtAGZ4G6dbSqF7kDAaDKJabGpL
KQ8FuFbD+qpDeITpruTOBaEy2Pv2d9BC5JhtT3zZNhwqv5UC5goVdCVv+JIYSTge
+82Rt+G8YtEoLYJ05YRynwGyqyKXzCVXkR2ceQ0J5botvKGnzulD5yw50uDAlkZX
EiozA01lNt6GsKyrMGyi9SYli5gZmq1qyi04L8zu7jQ8XZFsdXRMzok/oXkfbPyI
/v/xv/YrX4TRcbMiFw3ORgmvwsX5uWfhPFB1cgpw25zYmS3PPaGY/OiRwiV9E2Re
s4Zu3jC8Jb0ycWuPQn1ctA/0ZS03cgV+wKhk4CjK/sNfdMok5JoehTa4AaMCpZ2g
rJ2hjpYS07wgrP2Di9Nil/Bw9RV4MXvGc6g0GyRPngZ6NWf8L6Vh0dhLXtnMIUdS
+I2OUWNh4aeKIiyv4GJ0kf16+dWTf3eJ+lmx4oaBvcgbDbpUvqNEBaH0ZWyGmWNs
cm57PIcf56vEqMIrsU7eU/pmZIc+/SmxF77bCsBZbTxgx4bqrzzj1pd/BNP2Yfoi
9c0aL3R+1aJ3tPIWGhv66ISyrBTu2rP8PtF5HzrItv6WE7+TLTRFS3NJ6cZ5JUSQ
n5csLdhIuRxY47TDuoTtESGeTvCMBBDmZKVzSwTz2jpg5REd1DKyFwL951fmn0iT
F14WYz5vEvOn3ODCmtsHbqMuNrRRtlYfS/pwUH2pZstx8ZpGEIw7FcRUs4lxPSo7
TRGXEv0PrQJvWFDBAQ0diJQIEHj1NXQdostDXFBa93qxndHffN2qTkzV/ILX1XFX
gGu+DGEJieo4OfHHsL2u8+jDD3+zNh/IIWSKNtBtiarIDgCQ/6Ik6IjEbOey9MxB
+aZhf/g7EfZvq+aB1v91r04MF8Qz58Wjw0IctMcMVSmvE7n4lxiHogfI6UJt31Cg
bL6bfKPAFoUFGNxPsYgQ5OtzDnaqCoRJ6ToYMFSKvoExl5WEgTF4hgMIP9aVjbot
xdBs7PEVhjsHtyrURjmmoeFVjI2qhO+9i1mWaQg1jZfjRPEwPpwBIBN+LzOcsqb8
+U2u/bkl4HdZLNFu75IrGOKNi9DsVD9M9G30dnQMTeap0ObDcVMMmQQA92LEdNRU
5huMSU+73A4Z3+upleNGw4e46vTMbjywGgjqwgEageox/JtmJ3wmt7yODi4116mF
1HqQE2XtU8uoLtyds3+pqcoDsfdJZpIgSl6b3GNnFMOX8Qlxe8oKtRiX/4hJElij
lo7aqprZdM7ybHQqacDtDg2vxmlwj2AWGR3348YxnplUG37I0OUhfSJMiW6Gw5gf
AYIMsKa/6laACF0+wx6bPuPXnvk7mNyHoHeqp3ZsHxju7248PI/gXwiipPdDw313
kUcLLy7mCRsZ6EJAysVdLusC9Mz+mZ+RHvAXj1hfDcpz+FyoIXovOMhfU6l0NDrw
GckkyE7QKeiF6kMbufc++4atEXSOlsZLpCJ3dgS7SFe1kzEuttNuZJ1rxkAG4Al1
0CgjmOauNbnMghFZszzphGuUHzkMii7Hzc6MAPD8EGcNi9NtchRty21UAx126JQ7
oIhiPCm+C9pCtZzRjZceGAqaOidrcwWVqcftmkiApvcq3cZrEofLy+rMyKqeoh70
uyt0TExGT+vmi2vxy3B398omZ7EC/+zNd7zFdHUOikgmTe1ax55JyqsLseyIpeDo
hhGK1+D8XqMc0HtzKuueHMsnZfqUf9Fu+yzKsDFDt/F3UhRKoJnWMrS6hK0nZUHo
fAejo/mPPMHRE7lYRXzdCTIMvjDl7cMyU6Agk71SdXCi+eayRhrUEZYXHtoE94BI
TbuLTC6QbTmX9xJQAhOc6E01qXlTNG5pvbYBi9Jg3gHFw0CMN28ox3LD/kIKdAh1
ATzkPJNcR27LiaJpxAlzey9lPq/N7DiFad4QDdxXaT8c4F+JG7/bpYbGIdR+aL/C
Z/8AEwbykIBL2KHD1KkwhRJc/lufOfYn6BRAiOkC5IMmqNLSX9FEHkWiNVlb/E4U
8rM8h6+QnPvo6cKamomrwwXxNdbUOsVPNIEB1RgBmP7etx6T9De+bSD7984EHANi
A42jwi5HRf/Q5U1CBdi5/IE/BtJZ3zUaI5QROl/SvgZJdbm8nwPw58qPYz/h0xBm
NG+TF9q87AhvDWwk1TyKqF7sm1BJyDcUx27MX2T9Az42oxpksuoOQYeF7y9SslGp
4WsUD7hUTyClSpip8ANfk/qy37EpdYjYHw7Wl5qvXz3VhDjsqH7BvbrspLxqaxho
blaacIZS5AYG36ayQB+ckFJ5fKEpIaUbaErniqtEhHqrPDfxmfIlHgktu3MDYmMp
4pAqf11+WEPrRiIi7qttKV+PkmiMQFMlpKvq7mV0EfGjozqauBLIS/oHufeY2y0c
gsCt4oR9XAqWgyUwHn02PuoEWCK3dlEJBgkPFLx3NU5KT53KuD3IwQOqcmM9iyZJ
bHhR0olyz7BpO5OVqA2VtAkNmeakbZeHi7d+/M1nHqrEYGe12VPQgmPM542MKiWg
KL1s8vqHaRCrjXVpjDIAMhGYtqNv/MQhFz968QUhohp5ukpyjQHxkuB5zfCVdw01
qGyJLLEJIBxNzns+cA+Cb31BjxeLmVRgMYwqsqvr+S7pNOZcWN95u1UlowGA+CG+
ukmDZ42pqF7KB+h8nzcXc/yBkq2kmJdTa6+DutWTHgOKGfrs7Thi0KcvW18hG9DW
ZXxVObnQFHjSe6TNuFjxLFwA3RKdkTdz5yFe1SmQNQEEARVagKn/b8KbFkX/VxFQ
hzHeOVkzUGOvy12P2+zqxMyPeIKHkWmCk9y7rHcA9bRLK1FtLWQQQz863q+uR9nC
ALW4ixN3yRjxsp8ZGyK5pk0m7H2faZd4FaOZoOzypLfC4cH79xST94AUjfX+SJlv
SrSggpyZ1oR1Wq7TBpjy0E9aUuhUEHGwNjqy8wE+cMLOkqK4IMHmfB/LJ6Q/YfJN
ETKrQ1me4Kc0O8fqrcPOb84CAZisC+87cXr6INnkfZFuNPDUwGltznCjXEIMe3ME
mdn97O+To212KLDd+9cdUuFGPvnOrEHim19B2M4nJ+smtZtgG2s/azvfLv6G8n1L
19P+hpB1bepB98siXFQOrjt9b3JVYcOyU+SxvY/vz2X06UXxMwwzREAoKQBF0Hf7
weHYatrcCGKHH7w80mfiOxHqWNCfnBGql9APJxXRmO1AoKCXvAvIhoonjfPP1zaT
rREpp8IViW/Y9eadXYG66Z/v7mQBt/3UGRy/bbuz8gzERKuzVfZL1NPILergQlGc
YkZ+0ZrPgzEfAvpn4RJuRbaQzf/lOyYgLKHwx2p8esNOzjLbFvcJjsU6Fr39b4Hk
fUveev4zoBnhX6pY0Kuv0uvaT0vGxWvbTKpgspy0pC7JStVqP7QJejJpAUFDb0U+
MPMHp+raTcAOaSN3PznrIIpZD9WMwRFK2zQKX5sGEwAJv5WIm+tT0zaWQtpyvtMF
eiU99/8R3FwTL/J4d+7gFhlv3SiZaxxUTQW12JJJbx00l9YvCFkIkqza9RyflLmP
5ZxKFsaVfrPyBAM9nIcS9V0jZrAhRVycOW13o69eYdon1rlVSmpT09ppnngmLNfc
lHggfH1aYCe0c+KTW2ZCmU1SceH6iItRsPm+1/FG55YxRwrNTuLRNRuecyJTq9Db
XwSRM0/RaXYq2LnIaR/S5XeDooEmGEZJ31XucJVQoDghXQUo7FgNShgiQqusI3ul
AYod7kBktnapkrVdqiaLc364BzDwu3htFto533JZB7CnYgEGYOyAlYmmqcsHx+oT
dBBK484+27iYRwIPnF+wKCFAN/iY7k2zvKABBjW5D9UNacTFj2NjC16Ie52P5Edu
8UY++mYR6ALygt2Qh5JbsGsmwAz5st3QUkBHSnO/1jbqVDodSj3ZixIq/a3mYcLa
Bm9CT97qZtxdK3MTOysXSkc4QpaaMVqBXznxtWxtf7KtijUsZe1IEc5exz/k5Qs1
ptrvdO7QCu7NUvUQ8mOEQwmdjJ2uuN5xqR0px5gNmxicZsSfVcu4VHTfaiIY75Fy
BsvCPsIkLGb01wqQOaE+yO/yn4GXLAp1/9KJAgGj0YfrehnX0oX33cIzYnCDp3qt
B9cgjylAFtyACEbQOdEVQAUEpxAkT0lE9IcXBrzKy9otQClbARQsiyCJed5l0G78
rEykK89GVxxWvly19qW7eFlnvTi9MHs9u4xsA+hkCGh8qOoFM3gFkiPZXZpGxiSQ
OXVN9vwoXTPAA8AKwN5Oc+xbIhe1Vj8gwnDDsgL4w3pBH04Vg61LODZnc18HBctt
L6rp5iZieLEb5rAPZUsqkkeCnI1qAnepdaG0CLtJaEApm367P83Mt/twCsqLSlgj
lKC1XMF7Vaf4SoO0mi1WNqhhtIC7nhTh7J2MLinmaydDjuV2dgUCOgz6G6+MYR8U
3q0wgi37t/CnclZ965ek3K2YM0cyhvKnBvpFTqJ/9EtAl0ctq98o4kE0aUulgQtO
JVt90wG8z9+wyJ77D/aB2QdEW4CtTxodfa5yMTFJC7M9XJ/xTCKnY+OzSEc7+P8v
LvQkw/5LzjcyuwRk+v2UUjv+c1ik9mRVzAc7Vimx1L/UZkLOwe6sp2JNeJ3N9rdW
D57U3iT16Nzt9vBMOQ/I7FQvIY4iOp+6MHapvRAyTaVC08iKw0eEnVZZOxYuUinO
8uHCmvxZifuzxz4r7AiQruPeXrbyLjl9M3FFmN/CNpP5kItWcUtBNEnRFoQpzank
mVeqiLKHjICPCNdXWadKt9dc9rw3T/CNHT5o55R7jv6nnvfDhjzBJfCKCYOBayWk
H/psDc8pmyr4/PpaiWyRwoKm4lITgEFcg62yIQJQNmRNz1QjVLBlPAlbkpbf4mAG
WDoDKsT8UYMxjU4CDCiRf8jUNbw83Lhg+b1DRs3i7fimhd6s5rW9lfP+Z+qLOEHL
CQGtdGLw7o3EBX8anvBM/BGZr9LjZ7mo6U9aga6tVYXensc9QTwazBa6tkWZJrRk
IpzEJFMWrCBNKP5qOHcAq6sl/Fu3fck9JRRR1UQONvcoqTyphlkVtFlWlWx+u0Mx
oqEXqX/Y2EeDGfWCeTfCaBYSSo/Y94X23s+q9NfTwqn5LJM5ThjGAJGR7vzY7e6r
m9KNtiI4V0fSbtMBjf5xHNgc9tK+9z0w/spC/d7519dl7hBWQJPr8UsjORmCTXsx
GN8vyaf1BOLJ4ckZlKrqXGgx2ZeGe23u5eAQkwCu0VwgmY2ibzlhJMYQAqWrfbW7
vWoiMptz1VIrgwTqu7hREx1mFAR78YZj2e96cxcpoZ3R8XnaeXzWol2oMtU0WGtm
kRJ/K8yGW00lAdkP+Wp3wTfzL8Dza/KDLJcLBhFMiqfo/xqD4E35QG5pyEKJZBSn
lE/zvTydMq0Fdkp19sNLtwXIMevYIZhMaGuGivxtSwxqZ1IICCl+YwZh4z6zZQAi
RLkSFIygyzgOfR//nep6JLFX4JTKzxvMtPgZmzbcAVy1ryDI3oMmbn1KWRcmX8Us
j/de09nw7vil5pTEDs8mvUaP5TIjMu0sU2G+8VL9+MbJMfPtreshXDCBNEyhtCqv
PnZSNdHFaa2ikOQQgAhZQ8d1LgRpYAuV9OrJEJZTG+U/q6hQmI77LlzDdB0Lxax+
PuMB3AKZhsX0c0mqiO+4iFUTjQBWWEAZjqX6bkzSpoYMNUTRPGgvreYE/F2FiLo7
jTKA/lt72eZigSX5UeLGsSKZJ5xXJTbQip6wo6o+zJeg7H6vNvafKtxH4jvcJXZx
st3b6EvX458R5JAJ0Ol5YDE9bDgq3eDl/mEshM4iwy5nwpLWtiKjprEwAtJGEB/3
/wZyrtPAsj/I11s6jdA87coM3vz/IGYfgmhMVcS1o0cQqzDRYb1K8EnVYOEUrfg8
DYOZ1lXz1tTvfs5+vXk3WNqj8MMGC9Ff8S7HYl+g5vRInTmfr99QiydOlW44dTzh
Q8KPbK10tF0pcbUQj7Vaj7XT4lf6CEnKjCLHWuMzIyBNnzhTVdt1bbMDa7LFM2FU
UzJqQBUQLUNcBdPWAIk7rgvBuhib0lBFFag2q63nDPKtgLj9sBBRkdLhobCjdF6a
b/pZmH0AS6dGrH1xZZk2NZnvCfm1fP4gUD39m+sQsyJR2YzHCzuLRqxlWLvQVhD/
N8uM59IsrkD2PnEVnStnVINnpmffB6h3l61cLZVat1UKqQ+7gUL9vb8MKtOt6MPF
t7G7/0/6zSUGzppMASW2Gv75i0EfglfcHDPWNG6zKUr3Mxg/6g3EhPayUWKAQ3mA
7SE15seV/JZ6jY0gHNTkp2gTOmWxgdTEU6/mfJUbQ/uBp3n51MHsE8Uy+dT9Km4m
EGQVdcM4Uz9EbTKRvtt6bwPd/pEh10PDAUJm9Iv3I/6MDUPSXQrFrZ+/GV4Hy+zH
pEF9fOtQfKJwNOVO06E7pSdIysfIRygUpklgRxlnbH2q/6NJQCUOd3hUHnvpPGCx
hBhB4DxZO7WzVWGo2c75fZ/D8paFHrQPudPs9dmcroMkA0f8AHHGO1L3LikSPie0
FXxhj1J7ekqoN//shiRKkkQkmd8oDTdBf/zUdqqEh+FDaFwrFYdoHb4ySdtgXlJE
Qx9aN30eLmggLBsA29u/uy5lueJAxDmeBXxQ4+nHgVBGAj7EqlG5ff1VvLocQpiA
JLXUZYhdEQEvEZX86p/JZpbyxvKmbQeOhETG6jjZmZgEMWySuqpQ6s6w0uFKBxuO
F3jcubU63fiKX1Q3fhALDxq3rAtLhL1crWVj61sFwwLSyC9oGTbrlkuOwctEMbuI
CDla75HV7pefdDuVT5NDnGq+OGy9NK2/Dh+DESyC/+sesZHwr5AnGxEdhUB85oQj
uU+9mOTNak54kXQC03xTAUWlanc+Q0s5B50GLNujIjEmv2Xe6Gv0NMDh4uz6IHdh
auZYpmlLv3exOs14DKLN4o/P1NRokPZMYPkFfFaYYLWxD3Rhj84jfyaASzM/UsH7
MoNusMJEH4iRR6rqC0FB7fLB7JoM8hCm6RRh7aAw9sZFAtp4HV81qh93TFDqB1/j
V2N7qARZd39bPS1usVrEIRyP837o177k6/Ba1tl6qKqc+KrFARxoOPNv0LIRAm4N
sgqF7d775b0vfHFxwvNY97+u8DNRVW1kLqpeLHk9IASYZpjDMkQ44/xnwlcI206z
hRLa2sU31sF6Dsc9PtRZuN0wm7hSmzI2tT6nSo+NyheoxTqVE15Jla5a6Icu0C87
eG0ziEnRUVytMCUugv3e71jSFjP+MHkWsOZfsR28ajjYN6dHdErQGAj7L1fc+6gk
p+nAIZ4nvpe/o1va3/YdZY47ax09j5Kc4A7IIU+dvLHo/M+iB41xMDtz83MaJ//3
RxAXt9wvByjXAMtMFByIrk1VKzbgyYbcwvF4en/gmsjwpja1+wpmEYuolElj18Xi
BHv8Kmle4vJZyCZ7dmtSoz/wBgdDdb5991QA0RjYFlwjaxjFwDmXweDfr323TxVK
CQkBkSOZ9/pV3KfYn2Fr5l2GRWnWrHip4FdGYO5wfk3yndOTo5yS8wzfjoPay5iI
ZD8H6dr69uYwroe1H7fzvB4PAVimQhlURkRBo0FHLWPiAGtbd38UeRT5lTVgHufB
RNTqvbuz1Oo2DKajrtAJnldWDjo1Clj3/Sya3Pz35sIGf4BrvB+gQLu4yCGGIYzT
elpMz9/yXqiX+nm1VUeCIwy4vJHQhvApCDt7hri+n7le77Om6aKh3FZClWZYPgyI
2M6zPmq6reCam1fZ0nDL8++aXViowfi2OBLZvVbsN1IKQ+iK6ETauT3YYC6HEsjk
sZ7C6YWHU3/UDuYp8ezMXp2j+crTFX5erGNPrfz7HNXtmJYbnCqSKxITeMflgFAq
fs3Po0uLh90ZFqmzY4xRAHDsX8IQXMBYd4zxRS527gOFktSLTalezX80bp8+MyYb
Npdlu9vp8/v4BjAz/qP2CcCCJRxYqn0gaNuwb9tDBINiHt+Eee9KEEhmHgVoB/PK
CaqRLtoG2H26/wCNCz90gntipjAXlXBkHPppHpGrgdCzcB1mM06iL+FryeyRek04
bXO/daey0YYYjn66PhbWjBaWcJhd5qOxpnvGKkhJGWonacUnJUFtvNugvSe15ctr
5YCCiYk1qyO4f9bwjQXIq3s7aB5ZUZnzyzjRoo2vBuhIGynPX2M96cKzPnBs0Ph8
GlOfT6cEjok7Bgx9zTmz22QwiXA7MY9i+GX+O8w3KtQdpjyyeu8dF9cbZ9li51d7
+9TGOpv8c9PHUzh8kQM7u8tgk/6KLsUFSEgNTj+O3wdHLDjQtXsz2Ltz/pYN6YYS
aptn624dx424WQwlb3aZbDzrK1U/9e+m+FIKDXgz5pPCCVYYbNnISSFbqB0fAstY
7YK5VEPvIRXPJXzPoDgZlhUnGHwqRXPPXmQRXoJ7/aDgUmDhxKCwb55Adim+uHtp
Rdw3o4kL6Sv4/91ui9hy1Jk9hURoURTPwBf7fiOQZg/je/sJ2LK0j5sY9Nduv1TE
l61yRjzmj0EqUWfPcUjwZhkW8079+LQI87G4E+glztDLmcVlDof3wd44yvfW/EkX
jv49zTSmawiUM3bqwxKxr4myylyvyrDBOPXJKUcPwDecWOMogJ+IMKZvcrcgnMLP
5Kecd3l2Hyd5j3OGboOawQBkFi1w+OkIbKqTZ3LojP1kFswRSDysqbbdNYvql0gq
P+DOaGUPcpZFdeExfNGKrhQaVjbVyKQo3ubCGOyVjvyxRPJnBp3g4fQACxf+rwiC
zSBvo6/V7oz6awjmM+EnK3291Zt2AtS8gvKr7K+jTVIBOA0FMG9ffwl4OEtDuOAF
ryc8xuTNsrJqmXgR+SEm8M83o087ee1bb9HyUJblC7zc3qnmLoXNBUobUCCxDuYG
Wo2qtQ2B2a1bvOu6HkBdTe5rPhXzIzHYto3X0Y6zHtvF1hp47ZmwoOtQyr+dkNdn
K1tB4IVggsebHdGq7tbrQSxBWq7yl/LuyQY5oEmty+y0DjnTCcTI1g2W8u7LakOP
VD9/j+KwznpEFFUXvnSfTg+5418eSpXdqF7fHdmd2w4FWC9+I9MsQtDHZCSCbJ+x
ALc34dbvebUB6NfKTKf5XfG227tOUp7gKjrMLeCyxnWvCRwfoNYBU7EGpS3hwkmF
wsI8bf/FEgo8Ti/fc8WqjrxjBwUgQZ5ND9X49LB7M3LvFAnbe9iG6Vr4LeM9E0Hw
XyRxAzxEWmJ/Ye5RPiqLzQh9XdfeqANjFdeXlscOmjm2bOHa4e2JgwGW2pxkpozp
9+ZOg3bd0dLdVfaowp8rNiU/djD4RQlWjQgM76zARLoESlyYjHTDG53VFtuaL/X3
jEuGUd71WEUEx6QTqtoQ1Ukhi+MiAgAEliFT3PerUpB775rQ6QfKYGOM0Cu4U1gz
NeTr4i8h5RHi9UuwxTbsemujtGF9kFEiBgtzqlxtrrXK5XJUaAWiy/XRJaMHIbim
nj5hr1w/B2YIzKEP0fCZPRfaqcHQiVSnsAND7K/HNO6sLpSa9K92nMAjTd6dmB6H
5jjZkicH2x8lHobJHXBiJ8/Q0VIJJ1ItQxz2wfqt/032Cm6FfA4d+faHNTuEUq9s
B/SJNLBA5zXci/YQbLn5hDm3dTqkZNGBPj9k8ek1fYCJfhmxXtJ63BUwtn3A+lMF
29KsDqhYfkfa1nA9MPOVpNASkqg+1VQHxMaAOoH3wleJIly7uqT6JDGBnXRmHgpZ
Cj4tudqmJh4BBnbR9MB98RkEWReDoU+m5vaOF9ZxH9nYHKECnMMp2sE6NKiXiQIZ
3hB7iknZPWI1hGASIJBizOHkt8AMGu84bprEvYNOax82TqLjEadvMTcyuV4htU6t
czs0YzqzXI5FubrsnC8tn4hxCReylQKpe9bSluarw741hKvhk97Wzd6Ta1Y+Unsp
g/pUguWn/3BjoIMqXoYWYb1LSVmezUFs7a5rrBR+0UnVKbTJzYSI1H9+lJEbEqa9
ztQwlIvfaVchdcKX4v4DCm+H7Wh7+ruPCor0sTtcNykYlO59/oWXHWCa5O202bFK
YS/gvY8KOKqxP702S2wEkKwydh34qyDlpW3TJD/LHM9MYVW9PCiTPvz+EfslyN9K
x0sFr2JSmY3E9jQHYp2fT70LCpMzWBjz8nSnqK0mVaOLQebF1GMliooFCLqgHa1g
ELY+6c684WcQsmnlwcEQ8tbkFdk9ubHpOgYv7mxylCeQfdOId2Tumml1CDzeNal6
gjCmRpGKxoRXp3IZAE/zlmWD61k53/bGyXXX0icv3gx25qCNhHUHoquF+RdRFtd+
+JGpIl7f6yOfOkdEMaEE8ivWxmHwqtRcNDJYV16geaqT8Der4JfNG8zdmMl9DMj2
dxR9WujD1OXJp/FC7wOxnK1ZflMkRs/TcY5GDvs7VTu6GsYhpezn2f2wRw+lHJpb
++05Ok44aE0YjOe6p3URYRzpzNrMg56FjPQFpBPoOaeMnkG6uCc2t9y7t4Tqhwlq
Qi0wzs1Zf1N/oq2KrKV10HyW3kjESTLxSRjQZU03scP9e0hzf91iASCSlo4/7uyW
uBLGVs+5heCaycvdNpQvkZpvkz0tH+OmF+qlXTHHUuWf0upqITf2cNZPvPUJqIcu
uKKdum+snHRzHYoPuKk7v5gfr8ZlAzitUJtvkKicVTOAbo+IC76qIAnRKMDHBTiu
JwCThNZVrBeo27Wk+RvhHmaP3wPYn6sNvEQxtlWpNIRn3OiZ2ffsi2MCJfSGPBbP
iMk4siw6HbGSyc7Z01s1FKUa1TBkXoKanX0W+VzOoTeH7ZISFzChHB7pGtTJT/c4
Q7rlIQQV2dfNIVnfTRCZguRak6RJDvpdnD4VqSKE3UDhF6nGE4ndAcSQr15JUm0B
lN/CVDmfuKDb4Zbt8L6rWccjbo7uXTFv2smFj1mExPOJR9gCUITJMh4d0kep9Ye3
/GF9Yf5s2vOfY/KRBTpm6eLuyZA86M70RVhePmUdlZzmSt5Hw3H8xgnCTkk5lkcY
etSCIXFC+YPUy2IjPiTWWAPCHPRV4/cDHOi25zKTtz1+XuTJWYfIqKyA2qWv+SYT
RkOA0bxGpubvrFUNbTSUgyVeFFcrUB0LtFx51gY90gwulBqmkDGqlU33KwonGVTl
TY8XXIAImV8VokKxeVEZ0BuMpQvI+2fkFbkYS/Tsl6p61UhRANJpwmXBdfjnf7X0
mS2EbJ7Pu1KpMOIRyxzdfDWgU9tnh3z20mAqzsIlgqK5YfGFm/3XyqexqQLb1FET
ssxX7NVacoS8XRzk49+5/6wnVIKvRSoNNCVVSWAPOg6ZRPCKpH3ltJ2PqjPpDtn0
R66bO9HTIGA4ltOrc53gXOGZqjwGRZ1chTBhu1gHouwurXd9iPIXgsM1RSl13gay
RopG45njOEWrNwzg+irr/AnoqDr8sLkeVQAfk2wzuCaN1PjW1Rz68yRwFyLe6JjG
GMPnhABsHO7oMG9Ekt2RFl6yQ1cvuhYnXpn0IxC2gwP2fK8RdxTY20i/oGsxWaO8
KvyLZ3Y+qGdXJu5rRPe01Q4O1pu2d88DfyKAaIUUvRYlxZNcRqcXGiGyB8V72Q/g
96yPcM2Qj54X59ynado7R8CpQdz9zrIHlxWb+nlO21EREiiMZYXNp18h5GV+0pAG
dvF4xzcWzcRpkk8a6vInsJPIQYRv09NmNWL+B4AArmHEYy458fqy8/o1posLhw7w
zvTtA7I0WxZT4GZ6y0XVk0mYGJWZGJyLjeRl3p/zzW+QIMF1EjR+2UxK+Y8rnKbB
9fAmAsbk0uDvY0EjWvkRCb56OkdyJhJgyj1BQs20706wEVXgwpVUu8L0sZ/8qhGw
4K+Wdouwa0TOmXB5AwIduCKmaFS3UTvesYFB+G/8wHPggMUGtdkPmuaUBdz3iDxW
qEMtqXGTy1AkGbakw7P3Ugyml+bgDPlGuLuiUC5P7XiLmxnBEgAE1ZglGf6rQN7e
QTfdmavpdYUD4PgqQh93wvA2jWh00lhf6w7mY6OJ1KPi1fbWGV2ADUm1JRFrXoti
2vKgVudn6J20QGFIebKGgCl0CzIXD/4KjQHzrNaxt439M8ZI4PMPHgo2bwHtvFbE
jbc7PpEXomxbd7wDvMvL+dEflXyWIoLU2edLp33DwUBeVtDabUKyOiLzAItilL/G
fmJ+QIRwU3JfwzOOkUWqJcNoUzOUYjAWnqc+8OmRSwWd4gtWf/RVbj6RBoOdyALA
naA2PxM7tlvwTmmxsndNIOPimEw763togOYI3OHDzCU+cbX/qlshIUHWsYbTO4+R
8WRgabnwV2qKNS7goMMkgQAPN8XlvkO+DuzbkImcBFS32kRXvIXnowxuQwVGLeyR
CaSsx/f5IZDyVDBe4SszNwwQSvolkTfOFBVoDp5zQKMps8je45BcrixFP/NM3A6B
kAAbvQu5LW7NttV8IM/6mvmk+dGqKklWJXeLZmkRTOV0W9s9JqauSUN1NSM7ZuI0
gG83wD2LP48PyCQJlAi5z5sBDBqwdCPUdzfh5ZgTgJJS92fkzpzrbYY1F5I+CQkB
jH+ajs80kMPiMD5wlQQAVIOA1cbiEVtvUKYECmUKilPaokXJEOQqiy41xzWNgXm6
+doRUSDE32NIyJoxMYuM5VN0kkN45iJCT9bX0up43rofX2ZeHQmq37RlLGeuvrP2
HXI/kch0R3qYvMQ3NJrMMmXRfpY4WIM/NT3o1mQALFJV4A1ObJ9ZMK2YYxAJ1TAn
1Fsu8jpEkFot8xK/OSadtXDi+KwoFE0NlebPpZKFxoxlv6VK4tHxBe7flBuIXUNo
BpWMmIxI2z04gaijRJkOjU2e6fydm6iLhcdw0vUaXx0xWtTzYSBa22tzfYuEvxMU
brYaa6Acc2Ff4nAk8VpP/Szs4QQO8nSBQJBBUI1yAHH2gpbH+LjCJtm63t05uhTm
+V9dlFHz/IRGNqZSsgzDOIcaFLbzJmRRL6fvUMv9uxvq++pwWbp8R1nN6RLca93s
fY/vcFzjRWowqqMcaZKtZLbPU7bHuzuAhZGGHqCySs17Efs0BFl530hYn880il4H
Pb5otTvDdDQYMrYGY5doa77ViIR81cfEKdAJwg8OWIsdCh/G/Y2nuvZOBMUqTsIg
LldgBZtx/ZnzdHXEmEL033xeF0+NJjTYfPjHbmFm5I7TNuc3amIaeqYMjj8Y9Jdi
n3KkizQ7T4GSFkUG8IV8mWWjIqLNZio0GUVRRybCfof0ksHO8aPbRDJozt2rNPfG
KiWnuFgbrjBa6hNhCWK+58sLOijHawbf+t/KsXFMRZ1ifYmi62F/Uvxi9qvAXOTf
4Tigj2Fs1aPWKz5ccJFa/sAOyV5vJiBlSHKKZAXA5y+H9rSokjtZQefGrtuNXrL5
qgictdNrdEODoDb+UoVugY1ccgRDZhzpcXzM5/6/7JMHWRNv/igwGrI1faBnn0JK
B99mZcPINQq4YK9VeSPA3mXilP+g9PZugVQFX52doT40SONYa2ZKC0sf9xdL7bW5
ftYmpnG10+wDzDn2lZSsBlZ2iMyJb2YQaGzXMAPysoEDkh0bImG8oGwCVRynAdAp
ecc2VN3erBax7vSvqgsl8aIebY47KlTEk/ug8bvhoEbycB6363vfl6y9CsVElh/y
cJdlwbUzKaR0gfWN24+9x9yvNvhuxv29hqwreSpyciHgVAPVoQu5o5YzEJ2yK0xe
JcmDgsV0cuLLtoRze8U6Be9ZcFgcUkndio5WrlVywUrPKO8xVCcJlLd8a/Hdohoe
hU+d3FWutyYMTuI5E6u5oX1CAV+5B4C7AWmaTQkYt1/Ts1aCXvhVFasesSSPMpNj
BSb2yxbVfZvkgzHUW7li6PWlKQmYYkzw6eQhfGKFMpO9HCCw6qbCAIbFl9RQx4Rg
odxUhk5qsrDzHqVfzAnCtRANphqFUKf9Mys8YwzkDJWkbASnu34fPCMqIW7+BerQ
2WuaAcjgwBvP/0aMjok2lGaa1Jf8UE4LB8H+Vg4xfcNt2ZBcxMKApBzaLUdUnMSe
/DRoHiSW3LpJPOrAIzbzidmrfd0IwXpIrehj9w5hmRN0ljX9jbg1nHflMA4K+JdT
GGtUOsDFoe8ZcDjvXiu79tzd9fBhWl/3hygtZS+bFaWy/yWb7bFzW3ZXr18cw8ka
VZ8x9bcxWex1aZf0403vAeIo8MQi1PbocfPBoU2a7aR7Bu+PIj4xDzxUapF9hwjM
V7vk2HnPl8UmzXvmdDxhO4HXjoRiwUdaBHyKlXsLNZAP1WIkNP9cq/cLO9RBet4y
ZYXOW/aSOn15L9sgVjlYo5m/NJe8SCejY4GlIgUKM3Q6J+GsCddCuqiKjGi6FMIG
J1SS+S789yvpdlCjlehhyQLQNYa5lAc1ljm32gYfc3S9I2FPcv7PQIIYR0Vaz/Dn
Q4xllfGud7pPVwQzxV9HbOpYZ7C6Yd4MUayBTdWWfFQ+reVkBJhXrKRyuGbAoNjz
fC6bgVUDC1KZXKQvfec1V1odVtz6b6vXKujAFgqn1H4X7ReXQND1hM5veDYE6fq7
jGFqourUnBy0m8iMEfKwBfUkv5jyw3IyNmwOJQPgNxCQbMW5YPf1W13Ayy8H4pew
SsJ+GgPdNky4xn+ecsX/1DM1u8vdn2JT3qaVbf2C5SgGrMMWOd4VtD6X/NAY07rB
sryWWx+dFqEm6QgH4DrWKsfVwoDpoIindR8hn3TFLjiujweZ1yvzy/qhrHoYUX3M
40WpLWrgGMWEG+mLiuzX5zMk63jW9ug+G7HRUVqqUTgSLD9ZkWuSpDoXITK4pHv7
e3YTEXL7Ny2xk7RSMTFy1hLfD/NHNldJV88XFjlfE4qUAJycXBsQvvzTI2azRAp0
tzWDcK6JDjKGghLJOsnHEE28wbnb7fzcVOti1eztyk6N9hAdBcu7CvioFdBmgX96
hfkM0+1ETYDPgZYcXITJ1sM27erjJ9dfQ4UfAJWSB6em0s4CCRn8YGLZ4LmjeAb2
nLFPHIJNzhLEjF8531fXW1vUTwLzAgCKJQHmzM8q7oga3El25M7MFpF+H7duJsXW
TBneQ6tUfXm8QxZRbw+JGupyk0xKQJImBBXuRGWaBr3asGwXkWIJ1iad0PO+nACi
lY1tFe6yZJ3R8YpG70OsAosyzqVE/3FfpztO68rOT8nl7fHUwfwnldZjVLEcTZAW
qbrfdP6tkl7H/ZIdG1V6hc60fedUZ3F/2q4Wm+03FAckOiTt5mv/cy0rVokyO/Ks
18qDPpPO8TUZD6i2vsvZl8iUhXz+JAewTpbmi+7IhLTsLw0AtzGMumGDI/2yfScu
jys3rlRf4kY6CskhcZgvh8ESvB/7eUMnAlL9jUM0I1AQDSYHuwo+irohKwLNBIQZ
/KoWw9GQf54WARDEallvJ1/yy55gTVYCipcvDkDRL8Up/4tV7ImxhAACk5QZnJS/
pn1yhA8/D0AXDByaM0ykQh0sR/7PqI6Rr4yUwydGY1d/1HxigRzr86CMXWZlLUfo
81f4SaBy/Qw/lFGKUmDL73fD6P/V24rpsjm3v4VvTtEXeAieE7PcCRggP18ht0YK
AcLsexjaA92mcmUobclRKOHhVh9TzUZEgr/Socd/cDnebZRLJjmbwQ4YNdjsEzIW
NwYRp05eLmNX8Z6NrNRjRBLie8KXKx6sNlqpFjCYmrdrAAdeifJHBmxEjz2lG54T
ypJ9QGobLA6P0/ff8vuYL4Eis8V2lNBf+jQ2nbG7rz0jqCCbqO7neixp7HZoajBS
/3Wx1X7IZiF6WaUnhgguJA/IjlFgCKhEIZuAUqal8/KxkkL/kCrQirLGEXEPxQCT
pDhx1xd86rcrBcK/6cO4IzvJWj2g4TtDsdfdHQMkZQYSsy2t0cyJNbodI7cRuLeT
vyegjjrgqooeT+oiQwooRsxBsuV/4pyt8PYRXHlKyEHcFeaXmsd1Fz6RmMuVhh59
rhTMCrqMuVdfddbCu/X9b58XfduqmPhPQ/qnk2Rp92tT/gjFYcu0Tc6SbVz9b7cy
U9YofYHI3CEABw9b8nhM2n0xGeAaHY74CV/2W6P7qYwrW01tA+plhiVawX16mDSX
YKua6Zr+p+KWWMmVuktWmssxTHYqTgcT5Q1c/zkWshm/MeGT5s52hVwL244sU1JO
3Cnm3uzxTS5VYLSCFa6I4+roewl74OJ1Nfa3ufBKXZw2HITZlHGwQDUhLJw8z086
DoRx7uArG7KwQhfKBsT6frlSNUmgs4727NQqVbvvUlUkIV6skZ37MzvGCglVoSbF
RUaWPo7aQXdCAndwfb3HIdbvahIf5BtEvUE4Ua1UY/zqVXMJISar2Np+fUSR0Oyt
BYdJFnzpng9pgaXV8iqUcJDv5qKrSQozqSnRh+dZvmyPY7MRemi9U7hOX846AUnc
WIpfi1hmWwff3QOxskXwogQp1sN7BxwIpN/NHydP5czmpLY4rJHxJ438+mCojszt
S9JpYfdlSVvlnQgEtnwzCZH1hiVn67TlnSzty598MSBtACBiYTga+qFrslTULvI2
rS9TJ4u74IHcDPgTtNHzBUvcoyo/d7Kj2mb/yhqCvTVGtk/Doj5h60rT+nEWN2uF
oRTozZKHCP6P4K45KbxxpmYl1ozXMOzpALtgG29KAmy+VJBee8tDTBFpzjx0eEzg
VIVgs8Zqu1ZdXKbhAU7RhIxgextzXiok+GdJjzVjBe5sa7+AmHRgnLf9g6hQR7HO
Dq4F5ijqHEVVSx84Fx9s5aud/7wdEZUOBaDycsbrAhFa6ejEiz4Yp/7/jzp49QEO
zAcjHw4Xu2uAw7AW1w0uIg5Z2fTxOs15Af84+yFcGtdBQkclstCnxPmkNM23K0dn
fVXdygUFGSOJV/bWzhb1ciXGqO2OAvdpjglAcNqZNJL0JpUN+0xwQYqAYf8tMoAw
zfoysUZbDXv77AG96S3FGM/vjj3cUVVy4XuQJegGuWzyoErLjDvvbegyLPttqD1l
Tyrrb0clS6IOTmhZzhY9FkN9reWHrfec1uC7zatfslpPpBIXK+g76u7Ajf06mRgj
44gwOMimixrnrfSLq+xth3z8gIOSnMuZ9FI8hL6U8d6qz2WJSg8/Rf5gjDeH0q85
wYJoN6Gi+Qo/SrJsWxbHvNGUZkUF0bo3g9imbtlcHKY/TKwyhwqhIXTPB/ZV6eE9
DUCHl7AJbYUJhtawIXSeP7BzFJWSyXeMMzUGekdqX6C3VVBLmfP+j2JzqTp3zIbj
zcskWxF1NRfbdEKZS8uz6L1SmALkzUs+XRZHNlpCP/Gp/ju/42ru3Ss21PTWuQEf
rvTdES2CvzQSXciLCuAboAy2MMH/p9C0Z9hr4ikoT3+I8oYqkok7SSiaGKRiMfvp
4ri4+F9cae0Io8x+Qd1ZWUZPOMZSDSmUYqxj40FrjrbODMGRJTGWrAiL0ySV/klk
LgEytjomoDJREe7fuEGcglVeDtnKFWK660FqZKA56fmv9vRPvW6tq4kDoUzO7oXB
xGSV7N8pNkJ7kJ1oaVqiyWfx+kojKpz50bGweVyOgHhLP771mQUt/g/gs3uP71VB
DG4W7eal4wggtl4BuD4wRZ5MsHuRgxZsVylIhI3kVh/Z9qWafSVuKpQl3BLgB4nG
cBPiG2vcoAykVJJOU8Go1vgGjNoMsoOWXP9OS6F+xxmhehV1MxPSafCYrEkAB5GC
9rNMThNxSVSNsPEw7o1cUvlisNTf04bcotbA8HWDyJYOwHeB7W9VVJHO0nuqskfU
O2K+YriYB4x7Tjn3nA6h8vL/ivJirxBtw6wBAvfn7NFP5rRaEVlpbvoToJOk+dxJ
uRJqkvLSGB+YLyx2gtpsoepybDvyQ04R7pIEZ/MpaQ5V2z8UR7F34rHtpgmmdMsV
3kSI74HzJWvqhqm3z/qmZYRRQDIJj2WkrbbxTPXyBVWYvb6Z+2uJBtqGSnhNByMb
Nzp2CBTQwlce/9gqg81354OBwSFz10E8R/fbxNCXsw3Lvn7c/5f2otlgRUhx6NMW
sTtYqYqeucZMiXm8/XdJ1FjfChlbGkSEmFkwdsERGzOHrU+TJTV0MUWawNMjd8/B
qmC0QV+InM90Bugz+ZLJYLrzcdQhj2TQtZLbpKlQGbA9Jirq4+M27b3uZUzJzppM
PVSmTR9hhVQn7VDwbQ0XCR2bzldujwtEvk44UE+gU3nCNZ0hMTvBCJyugsSdLUlc
EtmCovhZiubkZSlpQi98n3RSy1/V4y6g+yn+Ee6LwGqcljufes35MyQq1QDPHinl
/XgPtPyarQhGfhaJU8X2S6g1XbAqq/2qg90Hvwpli3s5aCKrtQRm6ytx/oXJuXqp
dSEuvabAP4ZFULCJQkt8jLQRPVYTeknNaEBlnoglbPGNLYYTpWvgIMmJ6KzAI/cq
6Kp4iwY5o9DOg13SbVW5UZEab/Bf8OU6x4iscD1TLzc9iFy8oHHhPwtlSgnMu4kg
AOwq7xvG71ABBX7YCHVMhLQpK+QMrTBgVgJnd05J9pYb88vTAoaqb/9zYFgZotfQ
XgqnZy+LhBsR1Vfx12i9gLGOX4wCSnMnuC9aXND/HoETIeN37ztM1aG5Nx9XiEeq
xLeDgbZxvT06Xn9xKg+MjXQ+X0lwHoTR0FsWI7i+yQz7bOJU4U0jSvwm8lEEwBxE
2e5cCmE8tzQf/NCgnh1ckTNegyIXmblwMH6XHoRggnSWA1mqvCvl+sdq9U7H7Bzq
YJxKet99HRBsXAb3RcEpO6DrRlZG0y/kbqh3AFI9pbHaBaRPOb/FWZf+gNJJIWwS
x2v4EKJDF2EB/tgnym6JjDTDuvOHt/0550qCKcRe2azgT0VWb+Pq+VazquE8ScgE
dzdwHCflRZGaaMjOQzlt3m6fIMd8sa5kyqLdS1qWbMPI1S0ONLbiWOoxOnpTluT0
yMWzduODN//0wREl1h2SZgAZwJeBs01gdQXTvnIWnIsur26BeMv8QMX2QNB06dzA
2MnUr+rLJtOpJVx8DGxtusJANeu+LHfNdmBCj1Pe1ZXSs+0LNQvPeqpBSZl5kTNP
srGe1Z4ykhLBBs4xZNaH+B+Z9FDtlRg1HNnYc0ZEcZ7HlUgLGVbQIT0ilhl4kYh8
ubLqfBbVfGnq1TYCCKlc65ECNa5BSut+Orjxn8aNXpC2EPMFmlI2nqZCzDpldc6H
+6NHDsRQ0l0olnM9OSWrTxtVmGu2OvKbUPDUIXG/iGbr5YYhc+9HG9kC1Z9ndzrF
IdPDcPr0OrzWDFp5nPgjFIUGvuQGWsEgGpiWgxJ2sulqOddnOXDzDHvsQM+n1JMI
6mR19kmAEZjcvlFtm7uqv7SO5l3PHwLml6QY43JjNt8VvjFOTZGGLHKobpzoePNj
UFPU/rIRdzrPQ2zgFc6M/SBxAaMiKipLcTfvJAQPLdqNxCBg4VYnq8kbBXeKgFQi
mM3b5BbW58l9pdg42ONXkw4uw0w+rKQqXQ5dAoA5FThTI6RgyXVLq4ugvog7hf65
85hM5bfKm1pB3KqMFOir8xnKVYBlM0H2xDzfaDCaX8ivYl1SoMOPwGe+B1u+SY0x
Xi3sXc64gMp+aQjgkrNUsmN5vKSoujG24BINH/jxvFMMNeJLp+KnHE+un1UhTgBs
TW3fRjA9ZzZjga5UtdTaq4ZSMpDNJk/9rwtQRCwyLGzZuYpbM3apl7F6P3j0a8JO
T2QbT6/cSZ0g0ly/efCH1rrIstTbCai3jTwS4X/SbK4leWx1lOTjynf+NYF+oX2E
mZMc/hzw66d1+FTI0xvQqBmEgBOLXMP/2vhjsr7aZ6KjYmopX4PgxDCUXZiscUbH
XG+/ChrXjweAjd8FhILXg7x5mdx6w9Ufxbu40vC9rVrlLOKe3pQmUsBoVa3A+I+h
rfVZ6pwio1Ubq0CZu9VgRHOsHutJV9SQr2BaKgjiM0T01sLYKVLTL4ZZblyj5Sk7
Ox79s++L2FnUYTK9kyvPaXYy/K5I8dWHAngHDJ9avj2l4JvymVVlKyYc9idyXcKC
ZDMYHXIIbETF2Vm4tcydPzyw2IiUhpaoNUO7U+po+9woZW1ruf5Ln/tVUX4Z4xp9
gM/3+5lHXNUsbaB70bTGvgJ+97Qr04IdZKIP3dy1jWmgnz++Twl06uZ4AaC/b81J
Hjr24IEUw8ctLpBIDlLczAm0ewhvthc21Y2inHjwPVRGidXXInoCMHGFTtltDO+V
l54gGm84apeSTjv5gcZUFQrGexlU4Au4gG5Vwn+tTgY3cDK4pozpn+d61waa2HQD
WBC6VabS7aOAOj0ZTyyPPgriCx902aiaMhJEGC+MkJZVVTHphLoSWK5AQyhCkkBz
miLF4/rzuE25ZqsQl/jn6Xa9ytCUpwgpBhfxb/rBpdOQv+hDjUPhubXFJd6xmrn8
SM9ccN36DtvhphWfsgCpgluwRpjD3qsed5qqYtitSPLdCcV8kgUoSCUZYxJnRi0x
IrOX566R1N47i/Qs8VDwq752MAkDKmRzf66mnj1ECQNk+uR36spvUE8jgEnLOk2m
icHtLuwYncVWLXJalx5n3LBm1vOBGF96PN+XWg3jfl95i4MP4gW1JcFIobUQeCpj
sUaJyXVkMdYDBd2crKvrx6NxEvrpYmahv/OEusPCRiKbZyn2mvGSE9PvZWnjDhtP
Csuhq0o1E1GV3SPEpOoGQZRCVSTSEh0TVfzpc53SHi8EuOd55H2bfcz907ETdB99
Z3rg4B5wauUQCVJ/FeG4htQVbf3Qa+YwgDYA9piViK2m7Tpxrs878mWS3MkVbGDn
/I3yXqRtaK/+K1Ec4hcQuk2W5eCBXigZJvyxePx3MKF3F6u2iyxhmHceTO/NRvGV
VY63ls8sIHYK0kVaLJrXF3euQrUK7l2fzwIZxgfIGrfs2PZs9WHKiIBNSOzZI37A
KhHSQZPME7TpwGm2fTvpVbxoLGqPcJVvrQjeKzv3hz4b2vJ07VB37lKEp1j7JwlN
5+cRZmDPzc+JBAFvGb1Z+pZCGRjLKuXzK+gBQBqmY3QuTCiGOdCMXog+MRwYnnc7
FO0B+cxXPjrQ/NRFtg4awPumggRpNPOTB9J2z/997NVOZbNrVIFFWQ3W06iaCHKF
8xagxmADEs6gSO15whV/5q/MfN7fzgq8EPnMoz+W78g9t2jgxs1+oJBwJAQH31n7
NDugkUIfi0Ltyc3TEIGBwY8VxGJ1Zg8wdFdC89rH00bJvf5pzQuMbSODeU4hpIjC
5gPEimu0UaGzzbvt6nYj8nLUcVD2RRTpLF/kcpejXpEa3qxlMCxVuFUuzkJPK85a
Fz68dPS1mQxHFD19zO9nzKWo1s8EPf+4MObX1micLQ4XTgdx+giqyO6KLVeyDB0U
sIG5Qez4vieJA4ICIfSDuXBvyx45vUGqyXdbr+310+qFi4AluhuLdiJ7aawSfSDa
Vya+I8yOzp1XrAXUhWVjK4RawKChP7IMRhwaI49J7P2UPn4DiRWNZccMQNlHFw7T
2rEaDqtE3/hA4yIw7ny5CBip212izrkMbaizLpXktJ491SmAc0bWZGRGao3FrhWg
wMRghMT8FfP+LSMWv9/hwZOJiEFum/XdMINQ6qfYZ5if7xB7N5YYY6oXUyk28ytA
s/38ZI4ZC0vGI82vSQnjnxvJWwYROjWAo4UU/yQGJ8/p3jZL+uYqMwHcQFH5A6hO
sys/HUj9IUaqrIuc4uf9rsMd9MWuIZk7Nk93gnAu5gME3VPJy1Ud2JY83TfF+QHX
zHZQMFrtGIfhMhAOCLN6u/CCb9uCPT5hwNJaWych2/8cejOQP3sLhXnEQSJ0DRlo
CKeoSyEOY+SMWjTzH+TuQye0ylsAqFO6fAdazPZEwjhg7AbEwkhSZfMBpQGcwBC8
7kWVnZcwbiabAbnbiOLXS5abIS7BN8/zZiBzg/VPiupBUMC7Zeo3A+Oif4pQ4JeS
xSVS+cubSZMt0ID5A3JIN3I0FudjLRHZbvZiLZ/Y85fBpyKJz4o5SqoNRmYCb2DG
Zrv2CGEJpCUoyNn/YM9RDxMVZJ8MnCzdNAu4t/ZC+HIqkIYgrRZRFipB1mNOYH5D
itG+Vfv5U9D+gbXhQG6PP7kPupUDyxJSf8Cjdq6jDlMO5jEsdRaYJ09RZIo7y8nA
6JFBAZt28zoX7iwcot6G+tuJ3XuWP514gRIet9oQ18fpFHPwr+4owHPVA4TINdh3
sB0ixg49cm6+fjD97YEgQ0IN2Qq2iS8FdncAfTf9+WFd5VmwmXqpVxB9rIosskij
KAmiQe6yAAyfyFFNJyjHy+/O1eL5ju/6eL7JncT1aFlTc5Z4RsWUuEH4Ks4bITt8
AO8jXLrCCGN5cPHupbW5sye54sLtRtx5mBVSX0q3lIRDQ5oKpZT7EiUvzdw/kJ/z
t0iQtQ7q0Z34Z6dJwbu1ozm3HPpb+8XjySfOMFjghK7IONHCl/wG3vfHojXg1QF3
439sLVacQEqDl8iUBeHgeQYTE+jc078ZfJ2CRJMTVNmAWotFUTUFa2kenoOayAO+
X6pm2M0f5DpDDb6gxbgvlOKfQvENmbnLhFXVtTnmlORAD0hkDF61PH2c057nUjPG
/gaGFhYUtb6sUqxko7eOyEfUd3sYrabV5XbZuDZsQUtPn+alTlnUsEqq/MI5TUpU
Qiw/Adjoj7umP6rnyoFhAUuqL0RNdilEM+8i/KuBsx4sjB1/05g7iA4cZwbKJkRk
5vPI74SrcUohOvpt9RVYLZHyNRTOVHg2wnaK+XYNVaKslE/1RYsROmPBWiiScSdu
uc02liBb6z4EqSakqK3d18CW7KKR8Hk0dXXSO3QSfqA4tjw2QUjo2T/BzLLW+bgc
QR5vSxFSlFhaOmvctBg1HehUmFEmFHHgurEWCnb5aAtzYo0kykmWsypivu5SRCoj
12izOA0aDonkB413xHe5ki4fjkSyxM1cseJsAjUsPI8GUw3cgCb0QhEOi+Z/O1wa
0GfXIa9Njar7fuhUlkL85Cntb1XHJKVJ0dnbfZmQOuLQ99G6itR0QxqLPb7+x7Di
4272NYyUAduTIXC/SSixtFqZn2LImznRqlmfmdIRHkdGNY24mp4o7CHjRpR43QVp
u3LPru3sdgym5WTz36g2DeQ45Njlca5KLiSPcTg0NCYvrbh3xkJLFJMV1MeBxlpt
r2G/OfsnCIIsfZj8pPzroenSGCWJ41Diue0Ee38KxEk+YHj6wCwmhXDbTQeTiAIz
+Ra01cuBwAgB8qkbaXX74pX7FgsPd4JpUcfr0DaLD+vM+cNaf1aKTUHVg5BZRWZ5
7z9AnzFZX1GLXHvfxu7pVLWm58jX7AHyh0SbqBwcNT8kUHIrTEDdLEoJ3/gakl2I
KGUQpz7KDEur//wUWcF0I+kyUbzLYf6GXRbPniWORMbIYPEzUt4bP7DKh3nk1hxh
UAuivUlBeJfxwJGtGaewtlSxJx5SItYqXepEgT9f3h/2utsTOxSPQrusGm1/q+zS
tQ/8FDTX6aOSV0/DTh2A2ut0vnsbHRAhuc2kt8F3SH0fl7QZEmygGmt+oZPX9miz
/AalAjOO5JmZp/pqC6LPy/TV0xKZDq12IZ0GQo5MAfOh9sfz8N7JD824Y0LEg8Ti
1wUoLwzb3ywBfm40FeoNd79RjwboqQg2pujOICCK2CN5XCpK6gpiatxcGg3m9lj5
odgdiBmEX5Rxd/3yLnxyeR5NJTTMA0TE4t4OskzZVCE/5MEMJrs2/Yrhav72cqAW
P8LMcV6jIHi4Ld86biKaVw1qKgH/mwwTwpBFX4qiukIOcLXY/KphqXussG9Nfkt5
btN0JMHkGNwf54JSjTr0mhsqlR90CLiD3F523aVJmnZnjN4qvLh7kY6hYPspDPOQ
xww4GPeD078hOfFnKmj7C6YdP5v8WXuS8Th3ZI82UPGUsXJ5OjaSQTda1n6FX6PV
xtC7LL3bjOjVK03xVVfgS+y9hSJ7F3lDWmFE+CthW5vbbc/eJH558uf7iqfQO5SA
F8wtew5ZbjddZIxU2v0Hf5rF+k2+grDT6HqpT5xG/DyA6XyRmayJmN6DK4LlnaP7
+U81gc+XfM7NBxH1Bl1FncgSjKPQm75LJGi9WhHWSmnnBnp2dxXtCJYJwki5F/Cy
ItHHro1FZVnLNZaSefZRYQR5bx++q8trsP1mdT17aXZBXHw1GdjWOY998hX8nHe3
pNLRZE8J8eAkQrbtgBMuxsm9gALkIq+c12TRdN6jn6xF1NCFWTN5h9UEHBydodvP
6h/BXL9rk3aZzd0XWMHd7MpJS4EtGX+xjZPMMymX79sYVLjF+JCvqm8XGFQKVQOm
K7ZWhEKRn0cSqPgx91Gia1dzfqs5AdlvQlmyNnSK3+kyXcndZ/bCZHJzEjIMCK5s
12YYSivtJzj+5zJqG02yNB3Ghyt60yVMVheRDSYV+KQkP0CPYSa5a/0TP+TjSLUI
58X9D085Ffnv1zG/vyhm8qEYVM89rrc//x8L88YjwJi5alRJVilRM5TKW2NZCYpP
cFTGPZmzMK+tdczrO1swTt+eyEqJaAHCH0PzTGZ6bqYooJ5sSGOrxvZFzqLvSsAf
1/d+oOB8pgh6s5O45+52k6GUzKeOyMpFyjEwWHsCnhqGJHi2PbpKU7zE4f/LKiyx
vqHwsn/adtXoJA3TMxFgBnMlaWDZ2QUbgNzRfnl9lZ9cPd5edgfP8xaEoG4jpIJx
v7ZlKt00kd/RGT7izDLZy9MpoBhn5MIDVzbvGfX9ixS2wKyBURgM3EYUse30YxzT
g6y8+gIcoTK2nuGOoBN1ji+cxt/Cmx+3JWVdniIXi6VQyKKHvUbudgKqJYxvQCtY
dN6BUArnHQES6/pY+fden0JODrSXSA/hAgGmjd6VIh7+HEVs1ugL/Jz8MCXfNSV0
PUleZnYwDjdXJ94Ea1QW/oQ7Ks+coBgluGMoE4K12yysN1NAy9q2pzNtRMIo/3yh
iqrJzKL/BDOp4idqlaIFyUKSCae8uiKu/7fS7KfrvA7bhtalcID6zfR5OTd8Lu9v
FRUKOIaLZ6DXWHMSr3gmH06OYuVGnW8/OJzQxGvIgMYSLfvEkX6J7ZtInU2AUVRa
lwRf2ihAvMZvB14L5DLhHWQg1Yk+Z+dWXY1wYWTzXWZIc2mks9sb7R5f/Y4U0QvZ
Tvib4rOS9njjrbVeY9QmL68GBzsb45oZQeQiKHusbGy0okT+WCHymX7pl1B0u0qc
LiYR0+jo/XipxWtXfctSuv3Pi4OGWcXoUyHNGxVDeZ9u7ffcJIPw9+2N77WtQIMa
K1+0gb0YlkpEgJCZE91dCBKCO5ptB7xjcTD3illTEeIV5yfM7u6x0jcTDX1p5oRA
WIWOKkzvWU+hwT3MD5iUscYtZlagYf1ksGOQ/seCw0L+196XdvZIr27Pgg8w6Hca
m2Mn6lrEgijhHnvUEwGznu6SvtHcMEgCFUoOasEXWMj5zoTMXe3p8HR3PMn41YB/
WSPRJGCn2NBKJ68iZ3y9SLijJTV+MyOgL2gzkGDhgWyD+bXbCeNbYB+tWcCNGrgg
C1t9G+Mns3BfClbz0eO19cgMVM/fktEQSUMPRrdA4oQ6izMNvlIqjWNkVvGb6fEK
hIb3LQQH/X+2FQGT3EyL4qI5QcFvcDVECp5+Uuw7Fxxizh/eYCWCENde61b7i9dg
wUwXjOGjFNvjoi8PRjXnJHn/Y9ktrFyX80ymYr0g+gK4G6YwqN+ExQn3CxR7xIq2
kY1VT3oLF7kDgFaj+GJh0SDHKin2UtK4csk1SfCnuEErA2FoLuVff6wsV3YbcH8n
8G1ySHXK2B0OQZDJtXOusjnm8hiGHF7NB80b+YGueiWskkBvxKmQqYJxUETaaoSJ
uVKcwSSfEHAZkvwaid4vNNNArZxecVDNkun+2TBKy2dCqcxCZwxf2j8VAdjGtZ0/
DAV7+AruCqHXyOtgrJaSs8nMVNXw0SEklW+Ks74FzTYolKaLUFXXaTJVU0O8vT2L
vfcRY+kjvLPvDzk5DrKxAj04MAzCWBnMnLhOh5GT6tJG+usexZpz3cFZJEIznk0b
xMD34lR7D5uhUDlGM5HOO+FZSoRxpjVRGjvQfPnPITtKdouxVV1RYTSAJMTPiuW8
zpHCiIqC8ge1gGNblSMzmG3zcwKlru3dhahaREdXUKahOIOE0rmvMfD6XH2cks+2
7wpVdwGxrNqQFNL4XL2wwa09DdSap/FA9I1EJgf5I2e1seSBivCLRCV40JgfHteO
1rSg2plVGyn8nV8r0gAod8XafuIYRzTopuN+SZIAoz/2MPNLIvBWNRI7la4wdQ7Y
nF5sul0GXMUDsZkk0XYgxLH7aohuUWx7msPrfBZCgta4Xxu1fDS6Zi9umSy7A1sR
Kuu0K4XYIL4qv5ahlrFsRPidafMlhtrzOoqlRv2GykOR7AXjq7Ni8bzWEaQqtvA/
hzozbBt8kHkmV6vocbLOTO/xkGyRp9aRVosstQNkfOclVsvG3+f5EkYJMRT8ujVb
0+X2Bz3IGBOFJriFlClJBwumaUzxZe7ySoOmnt9+/EsaaMCl21Abi+KESgF6CpFT
3EROEPffDaRD+ZqKYF1hp9ndsSVYua8oPi2l9NdR4j/lSAVf6Dyl+oL5cFuXg3lg
DcSmu4TmfUI9ggZCNBnr+4tXaxyzdoIbyIoup74UsRvA2gNGnrRIVgpdkwe6KQwO
JCHvt2d/S209mH65T7EgSzFzDQOwEiehAhB7TJi2+gkvaUcwtb3vXb4R/hzL/aXA
tSWYUxNUOu13qIKeRpv3GgcIx5w7viYe7f/tDTusfizIJiIc2owBCBoZUDe6O50K
AFJtE/OS/ObxqzxXuhKJGb1qo5bQ/TO/F8rLQoFA/vgzin+3GEzyyka4O8mDmSp9
nBYm755FUJwjKvswyGvqtK6oDL6/LUAj4a5JkS8zUU3M8gTfcMLUVeOdyzQggO46
W1Lo6F7vj2+1vygzaACEeyzYFNzVSBbYnM/SgmD1jEME8n4V2Rc9WLZ2J5PTuDdt
xJnsVeVLSvKSwCwLYzTLdAxlrY2Du1YXRafn2xkrB7e+c2W/XMKUxzrAy6Nf9Wmf
ukHOWYI7CPrgQWk+nhPEGsCrPhha2QRRLzNwZFYO70+Sc7YQ6k3sEtq7iDRY7vOb
MNgq+hHW+HW5IvSt53P2J+LgUtRJy4SBTRDJS+lZKmRHih8TYMQZzrVvRzk3yxId
6rBspuHYDzwPdFzUuGpEM25majgAraqAVqJIJx17QqD0Y+2+xyYQjTZgi5YcA/05
TDBVI3nQwgE4PsnMjVRCAXLZakKK75agpM0f0nKQRGr7GQ8Mqz6m9DlBt0lk10Ty
Lfom+iXnoEFdJYXGg74gHIjDtvFxwMTFQ82GyV9nDTZ5sxYmiPEqIkmLs3AnBBas
LaZvZd5QT6r5qygIbkCSkCRr9fA1r0efTrqMV0NVnq7fpgQy31uS0kCxFe3yqZ2I
4/BnffL75bZI25cB/WmZGWvFNHrjmd1jdbaiBLHhyNZ//Edzv0EJLuSYwto92dAV
WpniGAUF56e3x0dvsncXsxjonABX0ESVRpFV/J4O8l4PgIXpOE7gV+PHP+Drc3TT
9zndKawSystyicQxTjsr2pxqopiHsiPCDykEsQ4WvAnmvmMuQroCfUq2rsHaZCM+
doaqz8V3YchM8DV+tQ+mHElW16cgo+9Uho3ikIWwTcgALTIf+cUqThSUc7sNBiYP
1RsQAA33x1nA7nO1KMrS+aHOLuDzCTtJEX2vyj7O3zr76mWdqRejw0iG9b+XM5V2
rZwOlaBMFfwqbnk0cpqKz6HTR8aijNmf/vafcGODVetelZ2HU9KmzrvKGYq/RA6/
6YAdyCf2QS2R/udHfPOZ2m4stuI80yzfgNXq1ueGW3VP6cF2YPv/q0hizzBrU/4C
Bf5I4jWypbbEp+fKNJ7r214JF/k8PTxV0cq8VyH1xGH6Z/q/DJnw9KO9DxNtZGxn
dLkCGZGkoi8/dLESaDne88NrV/GMGUG49Ax3TbA42wAxvt3iSkDkz5mMuiMfa4gI
C4XM7YbY4CVrPu/MFQmpDHpgAbrJgo8KPSkBA26fdFoF/ZTGkqOfeNIX84ZcXMlA
k5zftyrrn7o0WPciyuzCje5CxbtAUz6Z9jgMCY6NcXZMtQKRhqlxg+8MIxxTjlaB
Wul3X3u6HCAdef49xWWHqR1qupWRfwMhaEG/mSaZ2HHeWOGimgSdHMhEx+zFHTrI
6BHGPtdrCoDXgwYPwR8bnNxtl2Av+ZxupDHJsXG1cNgC9qjFhB379T4opAeC3TIv
yga/zz0JSOvAdo1AUDXyw6t1l5NumiyP9amr3Cgh4Sj8TrqMc0p0IKIIdPWgguP5
rkQqBkF61x7Epdb7vVkM/SunzWPj6PtqqINZ7iD9vCCpeCbk7Ygm0nfNo/ZUhZ3A
7m+nb+voB0WjYqLiPBFYTpnbliHSiF1i4GhIH7/wwVAXkAoo8HfiQKBjW95yBWCh
gAzD0qS3Sw2niCMB7wG3GcNfJO11+SaFumVj2+BP0JY4BWImhSWJuk9yAPzMGW5P
MvM3aS4G3iJ7+F3sdoGmxlOR24sr+XRX31LO3kEW1p75GwHIuUcwerHXulfVIhUz
8CVIRSHTLjyAtgZvNPau/uYulBEjaOmLT1CS7t0kd0fEazNNkgAPB73+YwPaVj8p
qdWxxs4L5ovZefB30cAODFcxyCkNe86CePceul1lEXurVsEaQQvQHqL7XH3bqcXl
AabswXShzUMW2l0aACOSJ55kbkFZnwoF7xbVA5d5AHb1WZ1fXUo8subpI71wXDjJ
Gpc/Z0lhSEboS8Q56UR+Hy74ceTw7rDnQkZ42rdchB5wvpkbKFlx39Z6zVr68/VO
WAjl319gf09D6tD2cwEBopVRDDYgGphkPuyWOVnroDiCocqdHNavVojw6rtJ+s80
60FZinkVVXlF7sZDgNyplUhALmZKZaWyNZICivFiB4KvxBMHxzvXKP0Gynkcraxm
HjIZi3e/15qvBdfSVq9U07g4enu9F4oH5O013PzPcm72018pn2uMChTp+5oMhv5e
WdxqMHD+UAaQXx5N8P3IEfMxEz4SbCdC8vVt3y+qHTXFOfjjVG2JZHnZtoFpyfu4
OdgIEM2dc82dC0AP1Azjq3yg3dRg/1OM5yUtCgDabktbnxbNzgG9vsSrvExH+hBc
Y8WjMCpIb0ScFTEtBDBhclWtzlOGsCmi8pwICBUyzzSYY9CSWWHvXiz05aCJv+lF
4M/Q/Gdw8KTpiM1c6ZW0wu+w2k/XK/Zm7DuhIFP2V3V0gp3WzzBHG0XMSIBdAkAD
+q2zW/l2LaPLxHr+AaglAdH+l6vTPl7kzanffOOQk502lJxsX5G9d7b9W4t7Akwo
LtT7+vUGkCPdK9VxM6jKC3zw5q0tvPsW9nLLpk2F+n3mEvW8K8awX2G3Iw/5b9Qk
DZQ8C8gXHghGOIb0kmywGcC5jrfFZhI2nln3VeBEk1tpm1Xn1CPPyX7J/bYmhZnj
6DpcWbQOx+nC4u9A4KaBdO6iDdRitNuVXmeorxpGCyf8fiOuiQowU2j5RNVK9c9g
/8kjpUzQhbZ6yC3WBlcixRApbXwxFObSFRjrd0YZlfVDPRGbVKWQqgFlin4cqb3v
KC0uVW3TTTPesJvJHoqQAZZjUCGd9wB43ZDyNqc3dWsufaVESQ8Y1wKn8MygucKY
63uzuQmWj8in9c1qWJLNL2ISZg6idaRYwQo+S0Wwm5j7eVSZTysSaDFIBQf5KTXO
gsOpo6gdZXXgndsvNf3X8mtRpGSr+7/nSq96/uZlZmFjr9D0/8Sy1ZcXbL+Joaf6
9IC/31GU3zlfaS9pj5CHUjE/4kHkM4V2OGT1xNfBGel2jU3Qx72MWC8GwaR1q8Hz
dwD3oDRTnLI3Yj648WcvJ8hgXKoAnjv+9ByiYX/eBiiHOsgqCR3FMQksKnnokEvi
DkXjWGvM2hdw1n2eEn0mW+6ZOPIS9FOKXFzyN0+Gvo0rqj+oDj4nOhfMtIbpR77D
siZ6nBzOSePCO0yM5s5rImhicv3Pb9ZmLyySZ9YkCHCzzTOrF/XovxIuuDoY5NEJ
/0mTxZuuOG6rkAUIIgWloYUZREiOpvrXb8wPRykuPFmHL3r+HVDwSVm/sAWGUZS6
6YLTrJNPm4Zu6IdU60tiQdMze2EnuUDeveqpFffaKTRtjzt1+OwlimpTaGiOsJgb
9zb3qxRE4wDkEF/RlFBVDXY0ctTrrJbrzVCqDM1ffGrqDVz04NasJINP2Xl1bNRH
QU5bthXCMxqaGTyhcZfTuZkxuoOvhthUel6MTM+ggjqHUlPfCYaWXU7M45Pl0wL/
5B7R+tCkymlkFA0q09kQMzYM9WCaBKZcjZ1oYMsgZjcvi9G6CNplRSNLRVnE/gn4
4IJ+HpvFzShkqjs78/SpKHLfokYktLLS4+j7hRVHKdue/EuZG4VGpGgOvt3qM9AQ
l1jEnbL02xQ1ldbfdkmtfDi15fs1mBo9iFlpifhBrmmspNs4NhzkXu53LwgFvXFz
7MTrdVAiJvByvEpecCn9+ZVNKskwM3nHAQTZIU+aRyzhysVQXrgHXSHjPRmLGij9
t98CwftgbX64RIWzC2LJW81yEUP/qttsZPa6hH6ONz+f86MKJspmLdiiUxcY+7xH
nTjTxijN5Cpfe7mYIZbT4tzSbS0dA8UcpBhYKh+VHTnDnuMtsTSEBzGuRyuF4Iu2
4mdK3g6aPd40mpNqskgqouWnCEuquFA41hU67C9FvlSG8f++VM9/VipMlOd9sDAn
mkxZG/YkRplfOhGoNyLsWFxYukoFofpvBs4etv62CvXncmNcxVAi21EsNfG5aUse
BXvVMrTn1SVBqwwvtp4IcKqty6uRiSPIs2BjhaZ2rXOCJOGpsFhct1TcwK24Enql
AMF9FX9/jg9mq2ssv5RPmxYTIwwy0jKUqSTfib2RGecctJu3d9tJhD93vMeSX6BQ
fjp8Z19hD9Y40j6kj2mUcAC3hH/b9OI9hazoJud1amk7wvX89lekVAmwo+BWvyDB
Zhs5seLng4wwmcAdIlk2zL0V01DaIt8CBuErZ7QOD8qCXRZav59MqSueKOyJ6wCD
vkSPVjCw1y67IGayuhQwc8RZI8EHB1Sji9PTiCaALf7VwcDcGjWPWNiJ/2UaQT6r
i0ua8AGl75ZF52PZT579o/H06zW2ccUeS91rWOY6H8V6Esm8zWfHFc2JXI6uHI2c
8Q73IyrcdBbpEBnSHClZxkJL+B+Y56hKKIbWh2ihtFYMJqLQlks4xQsSfD3Minz9
N6piFbb+n4cQvcqgRe+a9c4yuwnWJM0CxE5OcrKbFVsGlGD4lRCqORmDm7YEaDcx
5DE0E80dQDDXWHMucA4/rJWmtLxnne01uo2+e8ai6gBRy3Fk1ghlEP4V91reBPpo
LvZHjYMv3QRgjruociiljJCjEfcv1AwMRGOHPkNXUZsdf8jkRBdbSlfvWogaeCR3
3440bDBAdmNQb+BUqincFk4frwg6aczq2F2MalXAsZAXOVJRSGZYO369wSiLaszy
7yiq1rY9jVfWAm1PtCJ7WujA/HRT6v3Le3jdb9trDvfnsTa+lk99nzp/XBrKNv9D
cyqTuXyskaSj4QxsJyrE+XKyANbtUcDAB2xYlGNXT5QinMgFYMn3i05IrnggGPU8
vtw2GK/5Q1t++Oig6g2+XzqC334NUDEAp1TcKGF7ivQldiHIcNyWYUzJn+uNcjow
xyZ84JO2pbbGrW6yOdQju/Ba9I+M35VZgCsgsOZSOJkbbmik4ESMjB1C83rYw3Ne
+lKf+CLg4HUBLkW90oOWf2uUueRFbGgDRynbzkZveWRX4Tldt972ltmyKPqvfQNP
3P41Ur1ZwDzvTGynmAhe9S8o3cZhgItPRx8yNI/1sTv65XxiaaHXVFFBdtO3ngPa
rZnHZBNLERpdG/GmxDp0DCGcNVFIPwmXMuITfSxD4v9FbrHaxxz2Nzf+IIuw7wo2
h6AG6o2jxbHtUkH8+lYopy10AmpusyMol4nIq4GgGF9BKGxIBxJnr1cyPJECLMmh
Jy3VB/4emOtfC2004UZvxS9ughPEcoSdqW4HO201OVouumGfnZrog7iDnLvMYVmn
Br2UCkH9LgdCNP7NO/QJ9ZphDuVBhKrEdqUQSBv8UKQdLnDsp0BYYzJLHhiAclhR
1rO/Hp7VkUMPDKzstLzPX4q+E30RsrE0q/PvKBomc1gri6uD4iXN9SonFVLKTT98
xFjUxDGxQ05O0FHIu6kQNFZkiDwiEjXOnmpf6vLGnXc+cL5wUxrEQuieKkGNVO6X
3IYok8MTj19wfqJZ5eYyPI804cQSMkJSb7RT+yc33Bi342/IlVFyiPRAcw/qXVkK
SNhg0vGy6AZUtb12GtjZqS24fie6HVLuSBUbH4mzkfnPz6oCu4v3+sW6S9RKIjqJ
lZAdN1rID5ybUfF+3lJdBJMYHNVBwg5Fxbq0KgN5nB3Gz1gO94VmMK9Tm47HtYjW
g1UyLfrlDX7hWXDTKDYSfVBodZ8tr1S4PkABjEGty/I9xGjvC3DNkJYjiXra0THy
gFF+B8PJiieWB5bIrrUSrEY+gx77pZlG57JThOh4JosNkwgKQdac5aAZkcaAz4/U
79za+Zspe+y9ACaU39bf0eBJNOcHjOQH0tpzMq/QZdhFd1gCO3PDwE8fx61W6lue
kXUhHwIipLGlmzkK9vuHT4gn8SbEHfR/dJHwYF1Pk5MADZ4i+IvUYYbohZ0qeT9b
cOdRmC1Bp76IE3x+hcFpLlv8VCa0Ox/CdwsQ8lFo43yoq/HC+a+igBClbrkfHdyA
sAodantV197wG0MutHFIuaC5h3Xj68Btri79CicT1sMJapiBU8yrYDPNpkn47T3c
+YVWs5sf91qRvSXXhzEL+GkTNCAhcd2z5NIq/OH/796+X6ErdRAq5s0p/2Vuyw66
r1nd5CcM6Or+J6CU3mD0hQjtjsiKqUdEHTlK1F1s6NtFccpLBRcAiYRPQ+JFIPLA
kQpJ3TwuBoLyxQ/3VKbaxJHqZ5oP55eUypTDRjXLLy2WoWiDUOKCMRnFUYnYgGhA
2J56nOOjPQHItKRd6DwBND6LOrgZN5NVhG6CD9gzq8HIZ/7b9RugJQ1M0wrCwkt2
l2p2LL/OAszJ8a69FViTBtc+X1Gjo0rkN9x23uhmMnkY3vHQ3Hv4EqmixF1dO6u7
CDj3AjSb5S4QBPv+iNiqeTpJ9XqGyEiho7b0tRmiaOLA5nsnRYEoocI/2z4scJFx
sCbbNYvPfvSHfMJbfme5kLanowEOCEw51GOsRLEBrx50aWLcC+ilKankEHxPeKS1
R/0Yxv7KsS4RoWLn0c7EXSgQEuBYfRVUB7FoEUH9fIsjGsctOoKt9Wd5KRVMb3IX
OSNwoBWpqDrR9CM8YxDWXacQwK9t0ViwPcjJSoVQt9R4rm4UemmAXlOxRr39mXEr
oRBuw5ZMJtGZTanihr1XPhK82fPdHRn3u1/FWs6NnAzrEfayAOqA7CoKvQ+4R3KQ
Rj/1x6MyN27s5NwylTn13bitBILcUWYYv4QVV+zsg6x8TlivC9xlY059sMs1Bu7N
oRNto/ueRv0kcIxLsgj6Usp7lOXL+xqm7Dk7u4gXAcSaZQNHVJyRHOKLKlzpQyIb
GIozUg5/+FWK3E1kRrgoU7x4yuYQDFgZdquhl5BGB1MyApMu7/0ccztQXRltUNp1
psqUFdcZVxosg86uL1I6FvHUKglReXaoybpFS7luMTMuQO8HWdOx3oIp81J3Kf0O
lMRESrgRY3NSmR4GenvRRjueV+ZrwpVOCXsZh6CE5qxei6L6cFlg+oQrGbxuKC9w
i5mk9uNwV9W2uUGTPE9E+GtLYs3iwMiP83lNYmQnCiqfWtT4rT8Xxfn5d7OVjrL7
7rVjaYSJzR0FLa0odUJlVJfMCf5p9FH3LIu6+Oc9dJgUzBK4UVI0eIQY4Xefgc6k
JNLxHMak0/CVw/Q6MDQ/pWmELK0Hu48W399PXLMfow0+Mx6nXcXQpoxqzt+Nbtjh
torFIp1ovkW4La8JbsXBqQz3YpuvXCd8c/znOcbLgO/R4IG1Ics7UoZFe0f5MKay
ra4+qHI5YMpqIYtgLxZKzDd8O/GrH0FF+4WNTnIB86vC+y9Izaf0S2J6zdKB/nMN
bra2n2PWJQM8ylvwIjSynbETQxkibb8+fzT8tL+FgNp9v+VFiMxEZxhEjBBL54lT
DzQ1GEYLoipf9vHiTaiSZehGgHE3Hv7XgQh2MJ1edFEvo7CMsCTR5CuRHZiYjIqK
qIC1ja+MUHvaSMG2oosPF/R+Sm+UwsBeDFJsTS22Rbb2uwlLmZ3NTMtzh0UXX/DO
QZVf6bKEi0Bgjjy9eT7YAmZFj0c3qxGaA6pFS3LL4bZxTypaDhPeeWAsyAtGeEON
7Fv59ZDFWqB1tBVbCLfehWiRowiDQ/kknsP5oYClCH0JCuCbGYs1//+gieTnblq5
nGDcKEUJ3UWAMZcIYVPxcWHSv25+gmWCsl0iQ/pKy2nTp6Kc/i6v3GbhQsCxaaoM
otVTKw+0FJeXV57UYeZVXrXFtFXTwjEt48ztEZjoMQmNwGZok5ghjrYlt8tO6+6y
ltkk7SjHxCHYVU9Bc6C7q1xtUVRJUhrV8UM3HNOGdq3n5bODz1H+5+OavCZQd94b
JlgfSO3xWPdDFW7rPtG3JK1QTdrCLsA384mIePWXsdiNY397Mo1tmgeGMzo97mQG
/yyLBGtavJihGCz0+XJbyMY023yh6dj+15D8X7lMZQrnwZNY4NFec3/owheSR1Fk
sKOzkwv5Wmy/ChP3Ux3h0J3eG6PPqq9XS/JK+tiGBzdtrEoyIaF6eS/aQy36Mclb
M48qSoVyRSEsYv1UbuFJyN/eCEn36m7nEiYTs3P8xmKHrgYeYzmC0dx5a19yJwTW
wd+e8wk0Tx2P+GAjVzADFYzTCpTKrSd01gxQs8gHBvfCQIbjweLj3ZmOcDNjbLKH
ZpvRKQlm/kt1YwQc63wMYVtZ8xd8XQOWpZwJ29qaaUpInrnAT4s7d/yvpXeFvQSs
zaYohdvWacae9sY6p+iw702nNg/DkUEpTF9vUGny2TNyfQJNgQN7Mv1C7nMNnD5a
65097HMkYHBL4TXh9wGBTu35UvK8RxoP+bE9kzSGvl+OqfETHby1fUHsR9b+mHSN
GgVc/tdur6VJ/5vZyW8NEbayG7rosHZcki/IXIx6ZOwk3s9YpgIh4ZhwVkoLV9Iu
D+VbvizaakVEo0PCHWakcMg72AXMgBUbH8JlFuCNAkAdD+2bPnD6+POw1Kcy0RPH
+BfwsDCclDD1HxoovDB40Y6O7y3gg0Gd1UqJ16ESgNGSkKKTv3hB0shaKEFQ2UvJ
L+XaKdZTx6/N2ks5FbbNfpag6vAQTGo5CFxMc+24tHbQi+RQmGKSH6/RLdGprXRC
kBdldglnXsnIKn2h3UaL1x+pBYQfNzpMpXHLEsqH2WNkTEL2siJCD3cxjlxQ/B3B
VkHzTtc5PG5TblG7JjUrcFal7k7EsMpKRu0LgTL/QWCz2mVTdArV4T+BYXB657+P
nafOZ5sTdPun2vBzWViRX5RyamdYVIUlfr6XBf78RcrAUtneNkFG/OgbTdbTPgAo
Hj35SaNc4Qt4o14w0IdTHsziQO/vq8IhzvJ1Kx6BPRs7vEA5lLOWHjT3UYovaPLW
YJ/G84xP1bU1BdJgmfWqeXUdjFaeZYN1DfSV89OnE8vpKB8HKGywohW3SPA2WrFM
ZV/sbAs4EOrs10gDKYzBcixcXcNS0gJdcO4fQMeDIWdrAw4+wCE2d7IHUktkSkxW
bRyLnW3wv2Lj8909qgibWakxtAorAncWZ0xoqnZxq8c6hPNiQtmV7VsG8ATwMzQ9
eZmWMFGWThQNn5SWI6+vG3ykl0XxaRBXL4kv5NbpS/VIR0MGFpqTJUorYGVg2RoX
FkSBq9IQB+2G2AnWFmMoVys0nmCAv+JmGbMKjI4gKgtRtMSNDOuSNECPcCWfnqHz
b0d9CUcoMb1qyCS0rVnNu1RBuH+iTWyMdT2pqB1pk2jwG6mlUKL8uTwFR4fgQ0EY
hi8Id8+fnrMRYENUh4VI5+Kzd8hEW49IO/CxHYw2+WzkNX54qXYPYyP4u+SxSdiV
RYDKtgeQQ3Zcyi8LlKF54otymkR5c3VnHcn8PNva09kfs82HefBGXzIuFYO7n/0D
N85J2UVIPebbHgXpO2my3zYJFOHSS7KvRWAlCFA22aG/xRTtooPQf7q4EG5RbQgD
YA7fgv7avuDuKg3PUMLIYwo1CzITgI6mkjNNR71bPGJDzUqqQrR+jOrvpPJ6eAz0
0NVOk66zk27YLw62ho5wD0qs9kJIXvmlB9ywnvf+YgA9b9bgM9U0aNmSzv41jPzU
qAAyvkiwFzpYicEFqSj1+UaIPVrIhDGNTZucY89W+ISLJDm0C4+GOZ2QftQ6hHaW
NF5qAV4I3wIpYPARDdrbl9Bfkw/RAqITingfgmjeICYF6DLMnsEB2Cb4eg/uliSS
u9iztPiG0Q299UuTPmeHTpr7QvaNlaR6IdXPgWHoQVL4DJ0iwHhNhs7qz0aq8Q9G
AGHr2uwWrjxrtaeZxQQ688QFRKZqRLOE3XKgQoS122J4HSK7TBYqeokgRq6bfH5d
zl5wh+mAX90O1ayb3GFbCRu+9cRBUIBQUWZK9DYGZRWhe0UfrlJ9KSdgpmkDtIQ6
2dY4UBltqMYVR9VAEeRWprH+pjoNkNxZnu8WH7ptX2CkY8rQKhBB6G3gi9Ej0VaJ
YZtsjqBPo2e34tpATibgBKU6MPoAjKDW+8v3eGCYqP2A+iY3o2KWRSTtDPF06s4G
Xd8JnluxOm+7GvhNJkWrVv1EJYjP2E1Q3AxsdZNg11AlbokyceQqnj6TuK6GWCM3
W+REe/jFmpMN6MmDza1pktDUt8hb4tAIrv9iEpHfKOx6uawhaoeJ40JLb/mQ6PUV
O4NTpTkiYSJWqhnJbZpq6fBTc4HfDfR6UYjAeyetz81h/GYNuxi2OVOKtp05/bvQ
hk9NqD8/tF/vBHTkO/QfSbWM9V0C4ir4G9ihUGpLXpuNhteKsOGaLYsNieMLVozt
+9RPYfeZwzMOCZaq3iry/++laBJgXu7vnzIRYbLHL654osM1DppZZ+lkY9Azt4tV
9yKj+8YC7lJ3MSvSMQHH0axUHTSXJTexhM5WWbHGwV1je6lmq1KK38Gi54TMs+Nz
7d95MSfu8UD0U83dYmlBfUotN3rmaPhpJ3xuJHLBund1/qgs78VD5AYKcJFJVdVS
OLRCWdGk+heUTzAsveeyJaYqt9gQgtoaTpdZoode1vHiCbP/o047eSOQbuQ4HKqd
TiS5tdRMMQx4tmh8e2wrKeb77KGHdM1sp1vUTPsqqnKvgmIDHWTayv8g4vr6w/PS
yfboWrHKptUreBBSPZBsnup6/FFjpf2IZTbkDdIAi+I7RLZPaxD3l5lw91ZsUjbr
VCmc6pxV6DE49mZgpDHh3wi965/+2vBGvZnM8830pMVAI39yLjMONIToKz28PlVo
xYjiVo/F48y0/GS1JzMAGvTCBYcmmFmQFk9DzEl1ekV5DyQ/ctEwTrcSuZOXorUW
mzbVJ2E/+smJ9SbZVm+yAcobAQJ5Ys6sgmxDTlqVZu37muGzTE4jPzlStICU9ouY
h0CjcQw+6TDXNzUNGmkqIk38d7yVwlzygWgYXiyy6sqB4Om7RG5jpcfeNbZzOBFv
aoRryushSTO7jqxV7qLRGnKgiNXP4ZYsvYSLEOuMNxwzVqBFo8Bs4RiDh1jTT3In
rCqPVyb65x1GQ8PYDFr1R1sLroR3XrFGfZjFvQ6kjh2nKEtOJAO4EoM8F+E1dkDG
anv8sRErkb5n7Xch8E9vpkF4gYEtKclwWNEsHNk32o1Ool0LngZ2RXGCLuSPULTa
PCL8PDLlYrR6v2NLj5OVglV6oPNx0NFPOVPqSlvANFwC240juk8G+QV0co11J8FI
dEAoU9ZeFrIoEXdPc529zvXxlpkndXNRiGt91IbDeF9tTbcyzIQ2vcGDqgMnnu4d
thH180TGYBVP9DbgAMU9IQh/1YX0Hx9L6xyAuH9wG6y+920+uWr2j22s/bBqNwfr
QqCDUOM41liFTTKd7QhDKnbBzAxehAci8z7rChusl81+Tg+PwfbAZkiQcDYNpuBU
iTdx/rv/v8KOX910wejVbMX9gC/K56IskJ1CX7RxQSnq1wQqHKhSFVohoFb3Nezq
1owxwE6k4wmQMAvYv55eITOaUTiWc6d6pK53EiPFF2001d2MdQ6fM+3T08wdc956
D9GojLybEBcFAAOUGjrrAR9BOteXANiSDCkf4crvTCE/cLi28dHGO/Xwe7yeh+kS
kzzKeQPtk8weYHsxdwqmsnaIk4Cb4UyWBsxk/EJgATk8WzxQUqP4Ubs4UOnMZPqO
cvJ7IkwjZ2IAtSCu1spDJNElYzzPvHJRGStwDSvX0Z1cGO3O14BM9zxCvHntJlly
qmN7/nFFmXzlXM4wzp+eYpRceEPS0ptBtNsdVRAbRpVIO/AobOIAIzdMqWjCxnWp
yfmarhA39NRoI00T/kqDDnBsS5/MFmgDp0/25ibFpT2m09c76cknFOgPfW1iADN+
6k39KbtaThIS+ZgOFTmCJ7SvWgnMXWyJeWHQvTsvlIG57WAcTcjYPx/1PVASE4sC
mzXQgvGTem6Z5wEfkUSwzTvIEhnbxEdE7aMQ2THoDeECHyZ+8yq/ioltnfqHgqWa
us5R/daXEkoN03Dd/0q2MAtYe8bs8OMaD1i+lLM6mbgTIx2UKLk7h1htjkSm9xrs
+5etZyjolJoB6X3zWE+QNQB7h0MT/eCOoVd0UkpUtTPt44GWOt5R3SebbznmSoC/
1gl+HsW8X5Hmkeeqm4EF/NWaoSLmged7L+5s8zPRuF9+/TIqQz2uVZcs68IvMPRq
ooTQ78K5oscouyH7BvthUV2la0XXHsrP6MDac6p9DMwOVwP3bKJ//+n0MOsF+RfJ
0qA8r1/WnGtCm54XlSSUjmCh/p1qiOQnB0Zwr4Uls5xs6TJb85oU0qAxyDvgW16B
BbDHOFgiaBHk4emE6NyYvANkNzxosmLcz9IID4NI9drlLLf/VMLF6fLAloAdD76M
asl37b757CHfazmSQVH2TeVuM06FvJKk0qhABe15wixYyvxdHh5jnFm7TZcSKL3Q
kykPUmNxLnI4pUuVp4BH+Ewhbyg1SDQATVsJTi8CRCNBre703xprJjPQ1P0+d91T
E8KcD+/5X8bRQk8scHVR99j8iFiglaXT0bDUDajcSnRgx+CC5EolXmSUNt1mt2BC
UDhyjLfPvqM0ErG6/+3enkc06ye3c4wbOpzfW1WNqM5H76KoP6PGIP2sTUW8el0B
ZWHvIkkHJQ1pRJugUp8/yQdGkZfOYODCLjAkMhXxcfUL3NxSC+dzeyO/Q1NiT/a6
6EW6f2acYHi1IRY6D1X4q64jL3h7l4Sir02uC7PKQfPhBNDLX4I2ySukq8qLuhum
ZLLwWrOMs3xYgl0zpw0/elhic9AIuNd5UoOA9N7RLgNAcIEPYpRB1OkRAaLl9YPz
i7NE234C3TreX5pq63S8SKcJLoWElJMNXEvE95q6bDpSHHrJ/6PeXwpELeci0mih
I3kcBz0vfdf6gGSNWC6CuXM2g45gZ+rXus7dTXCzcmh7NC47LUo8N7gIvU4kpn33
tjOh2nNhEaDbLypXlwSe+gpjTS1935BgmEQBc8lkF7E/GMpXW0KjXWYtjQkqX9ZA
vWcZ8J4GMyS9ejIcITKSxYMKp22zArXk+53K4QfMKonXaeRYOGjyO/m7VRnyH4T+
elfarqGiDrGQTfCg5PlFimB2xOOzdNRYQwpid5Jqwrm4GpigVpbCLxQfsUgCNedQ
pqj4NEcyZMstrDg/CPoVzQE7Hf/RplxinaLT0vFxbIrA5clJmXYkNVUjXoX0EonR
tvkdTcbvuQPTJzXFoAiMsUzyFPE0X8eDgaALlC9OQ1pptXPgm6MRkKHwFDKYDSXt
ZRZLMx3fWJroGSTwAbWZTehr7Tx2Utx8hGcgphodXPqJpvA21QR+IQwU6AmDRQQ2
FszdUfy1uDk0lpve2r4ZH8u3txzGb+FD/EqTnhYlJOqVWap1kbFwJCalN33xda/2
LFtg7HW7QLtDQ2/p10EPxjczVO+CuS2F16+DKpAFrt7r+HuAa/dHZIU+V2JJInBu
CsOp/138ci3j+qOty9X+wPJpSjcIi5l1+KMFoU1nftU28GDrX3/vgmsJEz6u9Zrz
ZyUZCX5WGc08oiughxHKEon1CJ1sHyEcAl1EWJ2ujxWfvEZJ3U5l/bH9qF7UgoPq
iUt4vBROcvhye8q95q40K1Tcb2rnf8rtL25uaF9VmQ8OaM9DTm4nDim/Xo3ws1gp
fm+O2EpKMKcVqyiXyOiB9+RxyDttTfvMyjcyQBJIAgxn/dJNvykr8RRUiUjKxSuz
9o0TT+JOCwB98VsGcneWUeptbmvYjl+pnDwK9ZQLI2YCH7Fh4AIXueiMmKn0xLq5
2S116BhZmWD+U7xFDNDuQOxDo/hgVHmlec4bH5cCWSA7Z3Fyo39UG5OCqno8+5W7
5H91ha+qFxiemAPh3j5VnnDEEHLrySgL/ia0VC24E7yoNHMS96NhVjUWsGCEex7n
S4ttLSL5nKvjCIUdkBmISlLgK6lDZ0+wBR8gGOG/xVGN2yrVOhsB5+GAr49QX7tQ
1nVLWi3rHJEbtbatfCuQWVqi+PmYaFG10U6/H4VvC/cSrYHCGYxFZciq7zmW8ARl
2yKFZBoM/rVsXy8R5FmuTrZbFbQArR67RqPMEHEquKzrdYqnona7zQsK9JvagDjw
vAKhjdWJRNQo9mA3rjRua2LXBWzfDFCaH2tJXqPsV17gDp5C/XlfeP3cciMaqz2W
SlX52R9NzH9XWSneQuoLfK4OuwAXHfp6Fu/203PHEQa/0dsAwEBvmmNasav5KRlK
eMHcI2TFDV7M1IBW4OfuXZvzMsYbS7l0gcv5s6b72xWR065wLWaE5J2cH4Sr37+C
FF8oG4jp6ui629Wp0o3INaWMxfPlVoFJLsSMVxYqB8/j1N/sq088jymwkh0r85DJ
rVtirPy4z1YaEvhPUcMsdniFZvRcwXKqH8TStScer6eKV2Dqt8ATzVxMDISD6V5i
U7UJjRlJZfuvAH4xZI7QMtAGsCFM3xWk9JFZP9oMDDjpceEsjc2kG3JGU+vQEeLz
AHbys4T17pfJ8c6Brybna7gsuw0bidVOgcqwIrdud9J9xQlHKGwX9oFAesi3iTsB
vEoPOBvsOjTb2vrCSq9f+LzQB8sB4vzUqVpBLCxJPTGWg7BCBB/AXFGaATPbrewe
NSx/hMiRU1DXgwo3hkYOM9MSQqYpF6DnycU58xeXqLzAk7pE04+n1cSEeZa9J+Yf
WNnyD+uQv4IhRHjamhPl/JxlADKAY0DPbT6W/jRjNmXWV/dIoFbd2fX69lEsZ0Si
PeGtZToHfD7Ojr0r+Wggf+Z1zAUmEAab84aicjiZA2Q8ezAGJ9sTytRZdDq19e0z
oy8DFQFEKe7j2cpwdmRtiOSfUtQx44bISv5uZxCtnQ0SXYqDzudoYZ0r4ANkBsgM
58MPW4bKMrIcct7FtyEUpWwbxOY/Mz5OR4oXClPgqF/zgqk5xpr+Grd7d1BXlJRG
VTlYS6CXGfTD058C8M1w/O+pS6+hbokRi9wwQrEIuOidmnpRdtlKHrkKNlm9fTfq
zMXLbL2eySAG4BuMjc8Zgb0Bt0BseXooOm1/CxhLV+JK2wI5rbyCHCyPF1R4U/38
UI9S/4tH82TOI2rDqv3pyK5hmV49uoOtIsNBbPNt6VDaSB/ptTE5mJd8k+M/sCRt
Orht4XISoHc7eEv7mljhCbQsM9mBlDBIfmuRkEquqr7cIAxtK7Uo7EyFJB+hfwvm
1sYJIVmYpPgCdCxbqrkMFvybnTLfDH0I1e4BqRZZPgcAAekruDyQdhgZI99sj4DI
GByXDC2tpPZm+TVnWRqWw7n7PdaghdLbDt8dIa6yWWgtrgb8cIDUQoXwAyOtsufi
Vre1Q39FzkRQy64y8xjbK3r8xXapdn5ssz/1YgMMKfYt/ASZivQTGLJ1b7sx2s+F
I+zYuyE6ZqjW0+bIdx70VoawLGsPP+DWxxDgD81szNnfbIjB0UhQf0WUGZN91nJ9
hMXEValrqSJ8gWBeXqmd3q3nyTfzg3OWVHOjYbtbyUJZAH/rATLTmAwqksUSOzpM
Np2++BAoP4pLBsrcB+MCOtWx40KnPzxjG8W9BWaoBNv9L9mk82oVU5mcNJV+/BMS
TOfHQZBsGQDIBrQj6yhMUbJR+VDwe5uoP/svcci0fIFOeGCeU2yVGydBHTu5gQXG
S5Bzfyk2CdMPCgpKO/5BA7o2JzjPhH7Hn7KZZ/sCdnvqAYJJP9sgk+Olvom6LJ7r
Jzh53aSwlg7mqQPjHaJzaVVMwDIsXjxrYUqMPhkJez9jXEi1j66GfBw2WscKR2Qa
ENlFOVNVhOItzDzWiaYegDV+TKJc4hLvb4Lejct3QI/YElAFCPmy7gRIp+/EisFO
H4/F+pBYtirPYm1c91PZpNK/QxnCMid7OERBZM7TtKivLzrajIKukRfNxyhO3VFJ
gEiqB7EcQt1pV/Jb11B+HanyxgGYRiOfUbbne/YfFehJsSV8ccpeqsQOg1FKh4h5
c/cxEAIXBf4VKn64FGcGbNe1sh4lYc9531u9P5N6ZOFNJZwhd3ixsZU2HLfZ2+YW
OXsLz2nR7DmmquuWMjMrHuM5bj1IARX1VOP4oUKeQdogSVnnPrF06HQo1rHN77Bd
KatE3yBv1rTeXR3XHRYnnaolohxdccOdxKMXKT3aepHixsHRXqRhxR+Jnaz+ilyi
cqlFn2yaspq8Fxpw+EgwWcam4q2QASrXO8BKS/eLelp3uouNNFfT2lsY24NNQGsO
ZWs/vkzOZQ+oopzTIP315SOZN64bhwFLUJ/CFkJJ5EkIIlk+Nd2h7V7aPZgHlCn0
buAGch+UbaAimdt5pPqDHIupZ8VxaHIws2rACKlZ5GT2+EYL2MmImYWksMfiSfR2
rFmt8T2PCF9+fG30R2J0MW3kLeQWWnXy3n0odJWUmQR7gULWs/RNMAUnqUMbpR/n
QqrYPUT75JUwFtRUVdqSDcH1qEbWtf9PujeMtnuQPBM//sI+ydYyBvtw72BdTqoy
BR/65kBOdqAyDPTPw2UhYNYaWaAbXXE1CLivjWUge4iRr1xFNENm2Um3Aroy5hha
fRkZ9h0R63D4GT5/7UWHdxQH8npU8KxmLOkvTFEgjgBBiHxKihGObVGGy8NHRUfE
IgEh/n+6zyCJsMqTpjMwK8qOuAjBFJ1alfxachntxpV0YWoGaZqO+YpzJLRxbkN+
XU7AaeVF1DJhE40m4A6OcdQ1aDJtD+6jEISP5LFO4LpNw3h9+23pLSxNcZacZrFD
P2gdlQv7QnzqPOaxq1yHp0//9O7OeF38iiTxzRytprE1YhIJcw9zSUY4XSpnDsZb
CpyHel8j/770EeZpv9P0dy7ZwS27SdRkkyEm2d0JLgZJmcRHWTqWxENgLBl/+B10
LVRvMyXVszjIvgg9S96XeNXwWYzCPjGMLuO8oOFXbyxvK9+AkJX2UAq56XrpH+kL
IAgVNWQ3ZQLTM3X9ef7WEUY6axgfUZy2w1jbyswhlgV9UxwFDncZIhATNxNOkW3Y
HFkbRM2DR5mj8noT1DK7QCQQVrcA1InnUd4+la3BfDsKdQZArNTExTRwrADY+c67
VORZkxPP8vQ7g8sh7HwsbeEKD6dCiH4xgPcdlpyzLNQgdCFsB4a8DYUcYd2HpQYC
e79jCSD1KhiVZKPUSmMdj2cwfPnnpKiMPTsgYCDbeP28vWcLYyJ5dfxjNU5wKi0V
e45hOQR1iHe9uVIH5AwoQOt5Q/E9ya2m9/2u+5OxRhecEZHuhz9QXFktyk2H9CrC
oY7FfUskdbpLxZg0eKLEjI/oDPcK9jGxAz5SLzlbfNOLqn3z0QU3qBCnOzV+Sch2
6FZMHrXZHtXdk/WBihhtwiViraDbxebiH7dHIlM751ruh9CALf7zI2cRmATeLdj3
QltP97wGbsIOevpb0tzI3t+N2xX9kt+QJJrWJtIRS7nnzPt8hhBKJswQoc2hNCsS
Lu7skupOBsV5kgmHwPqIJ+PH5doC2KZj4K5c62fvAM/dytwfg1Gf/2/myJpKtgm1
W7+w1XPgFOjiVQoa3dSS9DTPCsDwmzHyFBWNB9ewuNh3HjJHE8GxJ8QGdeRpJnml
xC1uNMurxbAZmNzhF+6+2WCig9ASBSNKNsW9zMiJLQFZey6u5nPZ/gGPYNnofA8M
UYVPyy//WUQSVfXayLmms4gDtTV1oq5mEpzu3KrPN7DqW5CAAO8qkVdHjhYeir33
nHCib63QuOlR7KYRZ65u8+nZ7SyltFFN86p9tCpPHIwZ00DGWzL8uJw2Tarv/aMN
yaocfoBDEPBXtlqz177rJWdvLFgq5Ek9v/lHeDww9IZPPGA+FL0tVbdqKsjuntmH
9z5Je0UGVN0XNeqTAD4ZGNHSBagI0QIEEadY4zJl/W6/EXodkibYys1jeOTdMQIi
1LGgr08p6s3L3J+aKa5wgliOj9AvjiLiwDiE7YGMYTwBPLkS6BT1BisP/ByL2EBZ
0laRJMjc8p3Cciz9uQsTCkkqsx6/84q98mG9VNw4fR2ZhT8TfYEWB6adLDTgX2DK
Hx47ailej2pfD5S1Z1zQktKpQmKvXlhK4KimGfaKfEvjQTMEUka4JB/MMcVrA/UR
2UV3nGi3m5larjJTFThZBTuQvwmMy+vILrx1cgkHocJlWu+CkvMezyjM1PiojZOq
uicKsZDNNwXzYzpFVN30AqLBnETWUjd/GQGsSUc+4hLQEx3yeEzxTuoxmgTADC2U
AY2ENlFipHuBTgnQE5B/b+X5QPaBJNjWn3Hx/VF8p49sMqi/+kDQJbPnpIUMRoO1
uINBeFdtfnpLWWCfo9rlXJwM9b/VQ8H0Ww9y5TzLKJsxE/myrs9OjLKuIpLBCbJl
JVjUm2qD3xdbJ6dV3XoVP2vijPOl0K3vbSmMrYcmSg0PW+Slodoz5l6vZ/49kwhN
BM+me172bf2FhvcOQeMd7KgfjBISozmYcbK3Zr0HfpL4fHNjZ6Jocv/zSLQC7sEa
qG4LF8OCwD7yf558x8/2Tm52Vf4Yu0Td2cafwErBvVdahaJw1BP56bwpXlelVtf/
K0T4gLrjzlpZs2ixANwBkvElMmmPVUX+pka0sMNkes2MDbE0I2FWMr8bB+yVMrjZ
TvWoyj7Z4SaLblrLody/gG2humgoiC16i7iqUfnp4670fk/LsEJ64+Fy4NlzB0YT
hVc2eUo34rPHePa0CPW2I7CrZI6ButLnSNnVuF5MRyrPJZssKY6q9Jyz/z9cwcdz
nVQd2NF72mtQ1dYJl/3Bw0B24hP4SIKLCaEDNmC0GMC9PtIe937G+REKcOcl/2MF
z3NKOzZe3wobQzaDMHvzQDJZjz3Kz4wMqpDViFNNU8CkqqwSaIpO5fqRDMbBygGN
JYn17U8RzsYi6qL9RzoPBoH3kqsqAeB323c1fg4AwDCf/Nh70rYwBwFIwx7WuUNv
QkpXDf+JPpGvH9XUh/cUlK9fE3QkXAX5peaWOBmqOxCd0NS7JyeUJxuOYtFOUWQL
eQ+pDd34PwtzWXRj8EiCf+H/Tn1fpiUXN4A1D9QLMdLwEKeykbRgE2nQE3kUxKjN
1HMXnrWpwAOzT7989VeWC61GCgOh0nC0vy6rreSEJYtbYcJVS5t61H4nZCiFsl/9
ViiOodtQ+TjJyGzCzeiW19j1twZULNaqZj8oR5nnO9EKSxEvOPaBQcOHI0Le2A+r
ENc6XmWrIf0+Pf99sY13xU/wy+0X/9iu5YUgdNkVRtdQFuPK5Z5vt0vWLwrDwOgD
HOW/BpY4axTaRf+9r9GCAX4w3mBzUx5ZFeV04t1fBrjegPTeLlqpEPIiPaSC8fRD
Re3Dj8h0xoFb/tNXZQXuUFA3/hPljTVE0wZ0VTyubxjHd8IsTrEIgWbeqjmCH+or
d676NVTPiMQA3PlDyKRYTeq6bwdJfOn/5YTP4gReMRoHneDaLSFnDFvNV7nv9ypY
9XaHqWNCD8gprSlt6AVtrootlG9noGwmWgZu9kFRTKyjJGXSqc35SPy6GfNR2U5l
Md9aXcCvIEYvQ0lDpFw2ZjISmXzMG90bRYwniKrKYN51mi9UWGf02ly20HbdxMYQ
PuxhbCszUQm/ewW02gw/h8n9xXe/yKzgjBURO+OtRTQjyC+j2rJdaMB9so5PCcMD
gSdv8B+wPuRXKB6KpK4uQmBgClskL3D2fXhrLHKHiHPgayz+2rOY3oIIy98GppV3
IZ3eeWRoLh6LqjrW3S9TMLhLkjgIW6dDvJ4PVFTN1ojP+qETZku9kevp7rsKlGLV
/SASSJWxm3Dsyb0XqieUtzvRlYERYnM6qwXfdtqgHi5eQan0LR9Eyx7Xz8fpkX4R
m1TLKjLEYCfl9GpnmHOM+4yPcvqCZeTXXlarF9F+4ecP083SL/Yn28q/10iBGYZy
suiTxKjQ++mDRPPHjhcDStDZlKQDpmY5//86EjLYDyHtIIm7IR4W6bIOuZ5IfX9z
dAr2A4hoiWBkcRXMk7FdgAnBivSmavhn6vhZycgGopklnOImiPBQYzA6rzFGibi5
jeiNDcPeo6E83yuTK9Evi3r2HHSM1iwgaD56I8J2LvMbXBQ6dfitsunR/cz+hVGT
uftsnEIgApfvmCA1rHqUhG/cMeHIFy24v5pwDZGxVsQOEi6oz8BH6oQNpI7yjvbF
RDcSmpJ9GdE/9/JjnDELJpUZhd/eaNBxlEkxii/UzqwrXNWuSiA9vTJN5tLSRC0R
m8GV8/slIihwF2Fr3Asj25G9or/p03kq2mv8qU+6h3mcmJqQFpJ4aPbG9HAlX4TE
ULkQmYtS4ctg5+9PoOeY6wfwDyTSHF74NZDBgBen2gTPnLMmSOGYZgW9Vt5TwW1P
34TRu5Wuo7PkVrle1ZSM4DxA+YquAxN/SUHi0g0uEftPI/KjaUVNfopd0UQDt6EJ
sIWCXxV82squqO9Iu6G5GbnET65Rp5lpGRQjt5Otk+VTO7xayz8VFbuJq5DOSjoR
dvILcLUrqWwfxEcmeF2T4AHIBdgipgcChM59ilDO30zag+Lu/rt8w+s+Qxw86BxZ
Y4xWtTT5DHjIH4AEciq+NpxHwkHPaN+qjcXEePjhMf44B8IwrlpvX4k7C2e0AafA
PJIjvZgdpd8H15n2SJFGnhFIqhN3smafUN8PxhHofflyroexo2kkkT5i2sBEGJDG
TidMMPxW7YZbBMUiZZm28gMc+zpcdSoKJXcBDF0xA6XtMGWAw4bNzntKeeDCVZZo
Y6toBG+6qg9KEVLE2ZjStJvkUbvArg3+XhpJBlOziG1EjvqQdyO8J6aDsSuaXvSk
bf8YgWqH8Qz9ssXDxiv74PdDxaqafFW72vIWf1UZEBSbv971eWMs0vEwnnpnChaR
kGA26ioUgr/v38WRHGYqo7f8r/a1A9Dwm6TEjucGh7yNNQ0zECgzrQYe/7iJSpu4
cGFBycDd80rNIdIdp+ykr9JjKvHEJG8tWGfGcGuG/t4HHm/GfSMRnLr8jpPf0BqT
r/OXTxPOTHPRu5c2erX8uO2qkOhLnaaEV9avfhdLN7NKmX8VRCQxX62bx5t9kX5F
80/a8B1ly3gYoWJp6ijjeYdKDbzThX0GOyvMkSgT5IQQqmrcVOjUc0mXPtA67YqC
2SMR1ssDfjYuynSIy/2xWUNaYjFWPWqx762CZ/ujRfCbQdAkDuEwTQAt512ACaoV
YNccOidDTyXSRkAN8ZNAKgQImvgkgKX8GqLIE9Bpp26okNhaAOD8HTQblKrSPBfT
GWuKwZGm3+zGXo60G+Od0ExZHzIcDRYYBS30pZ39ChaAqQVST4d5+Xz8c4yL6JmE
DXB9ONIrRCsYPgTbHZJFuXbfKOg6uJA2AVNpBvIXOlWXrbouX0VKR0qTVV6vsaQt
pFqTx4CG1sxHcleShZxrg5+E+AGPLp9GMevoWtP9CdxzLKfAHnoubJ5H8CMQOJ1b
v/aDnYZrEb/d99Zh8jM72XzeZmGyrMU7Q6iP3J7303YrzlDdO8xLsGeDGfa7g52j
HwRjuToEvkUsI9xeBD8mr4nVWgoZ+sQhxirEQgpudlx4PrYLbNMiopWt1FQCJdCB
hhj5m+KYfDnfHTkEq9f4SKC+K6SUv4ZhGDoB9z/2AXtEAZ1M/H1EvIwJS78KBFXB
e/UKbfXzI8Yd6+pKw1NJbuGriSMnAnbJ/xREC4uOSAV8J6HR8hGeNnhbghajRVZW
wtuF0MU/qHjhvuhMCKR+I/3+ijXrPuY1FePpr/JLUUQaX8pEtBzJCpatjAkJ5uAQ
CwuC6sfxPhXWbFDIyN/XJVoL2yYAeB9H966KcI5ai4mUy6pAqcNm6y+8LhKlK+w6
AnZ3Y8q2ClKaLg0hYcyf6aXZ3xdrylIcLhmRyfllqmx4RFFvIT4+JbBF5vS57z+S
4SuLGDuRyEpm18jYc68GMppggRrPGyN7UNRrr2QQirY01c6rIsAcmIVx1VFuUD0/
iZ0Jtzw4KB2+Dx6R4pcdByeA8mh14RlSUqd0DB8T7ghBfN+RqW8FFNodeKiUjVHJ
P9kWluglLA6hKaR8XfSuTZ/N283UTtNZOTOHSpI2OJvcdncROLHX8DuVpjCzYVAo
PFFQvkg1LoRTc1wb/Cm9jSt/1SrbsxTHlsuhojcvfrt0haVWktGNSSfz4C1XUE5G
1etkzoNDsbmbt2uQyyX3vOoMbb2nWych5/8pEI+wqWUU4DbCf+ioX1hJlcFKLdHM
xrtOjZO0D7YABljuOrPo/SqwCng4Sfiy/ExTgTCeoaJXH1+kd6nf3ts76IMcZ6iU
Q8kxS7bligrgj7ZoZA+SN8PCxmWKFTuH4zLzUukyra15vH8Bi5AW2lDM9e6qw86T
aaTLZ/Y1Acp57pDzcr9OlxXbXwpj4dpv0PWlOZLpVO5VKE/d7iB10pX7Eh/TZCBB
QzceJ+Ad2X6xyoug3/kVM8Oe2U8VMZuGa8XSoxVC2uq+KULITqDjlnT5X5dyIpOH
8yJImo/VaE/hx3wMcPBW9/8zVcJE+QkxMRDQ32JXrq1m8vH0cs/9CDUpbUevjhTR
KwnKk3hCBS3lnmfqJovI4BXJElHZeOVRVWja0QgyIiz5kDtKDNZuQu80OZQBx/xu
vfIXLy4jTABbSk2Y/2Wlv/hxXnrw1mKnc4riqYG/Wifw+xfWPUM4TzMGjFASOPb5
x7jzOim9hwAtgMIlPcjDB82/iZ4W+U6CNWtl2bST8KLs+3JEhyS3hfKaIZM1e417
gw2ji6ZA8FGzyZOU8UnFLvQ+pROVZoFXuZkus03lJQ5HLeV2yZvbjlMARdV2XeEg
I1VQwi//3Tz5T06XQl8PtyehpT9dgzdlDDJfVErW+1GE5/lXRNdljBw7DscgbIAd
XfMaTgwKt16JbA5HwPOPmEetfhgkpLXMpQqAvCPHtKfyBkKX2zGbTkfMkXlFgATK
2ZTi0JiKh4wOujegqc3OKq4nL/ddwr9DemmV7fxaGFmDXYvldqMm/7NJLEvSAj1X
HRFETj1eeW4hjp24OPbcUYoDorrona1xu0fVXRMoTysCBZ+KnTdqlP5X4qA5dDt2
M68H5t1uxBnDbjNh2O5hbHg4XYH/KRQWui0cWjgW2P3msmBVoMB8rGKlIl3Mhj25
QJwzu/dKF0mZssPpgB9rouHUPmN/O8KZREIcHltVSHhIAbwNnxskFjOppiyJMhBJ
z3UdQOYkL1dsUv4/PZz2PjIOBZLG98Y1p/UGcDvfhVrfSxvdvAnmQhgLTZ2eKKcF
/TpXMiSbMOHCFO0iGNIPaoIIjw2vLb610+pUVXng/0oOb9jk9zAORqnKWkco8ISG
7dmtQfex3Oo4W8i43pKo/eAYjR67Kc/sUh0r1GDL4Vmxd4PEL87/2u8x5r9WRZPo
O3sdAiWTZrjYxQcVzFEq9biqr0VPerlu3EThoGBQ4P+9ssda4mW6QabmQ1m1SAsc
SsJMjwWlCyA7QOjcVkMCyzTFRk1gaRKn4q1lmG3bLfwTjRNV2L+VV5x1U+lJX+KT
DSiANzWIusbAdB8djnll6zJ9rLHEsW1hqebEfZ+BadtCp3VJ5BiqriIUisR97+0e
xSA6GZP69+UKctm5GkP9TgRV98YRKbnEeedNzFYtmnraBhnJ3vDgls3P4SqqRq9w
jxqENlxG90HkSe0xSvztel2Xxh1SzVtaWZfFc1BZOoGWxXdTKTd8xcb1Cq1Rpf6c
LhTGfsNCUYRv6ZG1bOVr9v9tY+YtJfzv3s1wMjEutbt/wk1BrWP4cNqdUn70jfVq
S0aG4FPgubU1OdJO/67sCoWK2hadleHaHne/F/oNDXKkg8nT5t9GToZYoB2KLPou
CgV81Qh6uQz+9/ExmnS67lVWRtUiLMHIdqdUn+trxOJYw4krlvxMuoRXvs8rwcMs
NcaQ1zBwLLzlgTxNtkD9EBvg/+/t04zgdOvloMR9HWIQEKVlovx2dVX0PmaPiGsP
AxvZ8uyjM7p2vDPSNDZjv3IarcVUlz+kDql2i7tq7A8krxC1PQNt+1s1rWKTglbs
gBHfu7deV8tX1JzdxhLfWztW/haQFizoWQxalEaclKaPqrH6EHHcskvZyZEU8tcR
xRQdff8z9SKFpOcfBt/nLuumAvbli4cM9/58XJahgfWGF60nrB9eC2dOKhJ7Ok40
P+rBgliVB89pGGpxRREq5YjaxOrl66vrd+2cj4EvjlPVMCBjQ1IJz1T5N8aGFl52
0kXAK+E4O6zgQ+KNWzWhh90CeZT4DUbo3wqAScSeYojiWrH60jm87tdMlFuyt6ga
RF03k5C0qsbZzqc8NgeE7BaN0b5TWQC8O4tEFQ+2VTUDWPi2a5PxrIM/CXUd1BkQ
jUQ9jX+/w5VOuVCRRxEyWniPMUs1gDgI/njGc/dddGitPUXXbgx/6ueV8AAOJVr6
j6MTIBppZUxJwBAUB4/PVKpPXxj9opIgwfUrAX2umWMvFjCFz64kEo4m1BXiS68K
ZxzWdI6mqZ8IsG6gLdGltY0aUT4eM6g98MtYVFx3wpQk0kSkIPARKHvUbW+We3fE
/liQDfV7EjaZ7uFSBumBTUhc0QlrEvlNKPhxp2Dkn6JttiMYuORrMqhvhMBOeIU9
LRVZMJgCO5dwj9p3qQwH4xbNCIKvipABjbmK1ngaG8BOtJSm1/yjuJdK4RY6b5S2
G28EvPqE0s9h59PTV2XytjUoP8UqQX7JVhT3AzeEHcTeoIyrecm9h27RBGRDIK3r
Yobhe5XlzvuwMx3KdAT7HAPyM/Nvc4rfuD813AVuyfyG89830g2eC5hmwYoV/ES6
Jtj4GfLksxCs+byKAFJw19BvapwqFXSSHKO4dfoW6e7Arj/YuLByEG2W3ZV4koe8
Qw+Vf+AHN/OSzyToGwD8cq/wQL3CznrG+U8kNHCJNnGVZyFoJyURTOu5+NkcNJ/V
nWFWPNLYZo5QXLsyKOY3SSIHQl6zVH5Q3/+jFO5fSGrjVhs7xRdhaDxFzeEmN+oP
fzIPd6eggShL/dBRME3tT7e1iImLiv+QFcy72rhlUm2KjXg6rsyHnj3KZ+yW/qao
N8GfHIFWtedO+9RtCeFxbDtMJsXRU2EbqRJxFkTXyfvyUghYiTzjYc1rrLG4i+oV
8m63nKSotNElSX9DZdSP9PWa185p+RvbDjwzZNpiRcKv4OtD2JfNeeI5UWq18nk8
FMdYAqwmOfsIPqu+B18TRejvF+p91woQz1WZR3+o7HwXUkmRPABTx39lTfh5AGr7
kPICEe3XJwmNoljcsXTT5oobeWi5rJPVfZuqrnzzD9OKYNqevFZzv48UXv+AWr5c
ZUW2toz0RIG601CDZ/EyRaFux8Vr0CKoJa8vOgwCrqiUzoFYWK+6LG/gu2GOu0E9
Z02hcSe22xpwIqpV00Cs3NeSfLCGIQKY3/4kLsSROCPWnO60+Ag2A3CM2AYho4Vs
mG0YPDMW6YfS1t/3uh132vq8+cficgc6s5xcWcay0EO2WtA2ZWs9qQ69lS1FC+FF
kTmtAWEGCwzBcv4JxPn+pFUmXV6PxYyXDopjCQTePcp11v81Ib+26cqyrGJA0Bzf
aRAFZZUI3sN6sez4b96JCIOLpIRaex+UpKPeYzYsKSswlwr0AB/x1g/FGyN3d1Em
ycbMD6olD00ULdp+WLKulbpaImqXY4302LBLFEbnwzNp54/4b+Hi/5MGhjR4pclg
w8mRBiW28L1c3SkhVqWCJA/lBzV9sMYlWoljBYEg/9jgxMYIJHh639Gn9cDr3Ke/
JsZbFn6TpV5R5gde4rBLxINrKQYrr+q524CXw2EoskfsABTnWyashsPL2YZnB/RA
nGTsMcTshH8GExb51/aIa5+I1GvHURpCjp/h6gLIR5p6I0I9Ck9U4ntilGCxMK6n
y18c0kMb+8VZdJ4PjPz+64UIuKaAZ/4JJXGAv9r5+p1eYCRcmT1FboFC1Mp6BCxU
1vW1yWpP0SLqxFTK7Nh2r9IAhYKLaohesTc2AtzTW15qhapgztozIw5wutZXkpuB
dqW/oGIx8OLGlXtVvuS7nqALCVRb1AqEXVo5Gtmt71Q/5egDVArz6F4Z1Tgo6pDD
d6AD/+WVUgZUlUUa6hDDo1xxgnPuhZNqLKuvhvR+7zp7k3mPDpzTO/DJl9eGGA9c
SJgdAsy+oapIbFb5laakxuyHxH7xW6wxuxzDBXi/un87BeKqG3J+Z6YuChHvV2Dn
V03BF5J1KTIy3v9p0IiI6c5MCQrJDk6Ag1xFzgJjSK6PPX1nA/V78X4mqSRmdYlo
MfkUvNgux30XHsVGemVi1vlG1vmaie+7d0Gj8ex7qvYdByLsklQAMrqFnK38XbY9
RB3US2Kity5EbpQBOLo6voiF6xBOY+dp1Godg5fmhVzuPz8m9nXKg5CTx72UdQnv
8fF3ll0l9MHGnRh6t3ENpDVCRzitSaKSVaw6Mnb2X//XgcSDpC5HRhNYPwpJLu1r
eGe7yqqNtNVIVXxiZ9ffB0hhD1OnNxePRy4hVp/Wt+Npgx8QavYCgsvNknoLSvQu
GfpHsZdQmefkh1DBg+Av118Jfpnmh7Pyp2GHughW/Bpqc+glhwEwvSVPpKchRWmM
wqe3FfO2m1/BpTuPr9OLbuTrVj659X5cBC60wSXOOVAT78ywPn7hP2u+EdbbQRgD
PBRzBUPlv2S0oej7/w/vrRdj+mqO4UgII2yC/gJWUUrKRMqakeTbPrRcUJ9rdlx/
17tXu6TtFpHxHSdx2MpwbMFZYqQYFI5cg+NWoNIfjNDdmeqtzCPUZaMOBD7ZdYZ8
ZQ8gH+0DXv1QQx6qXBIySodXfYYqjk89Wmgz5zGQL/rLdr3Q5Et3egiffZmGoX1U
80Kk+LwECd27gNR7tewE+8J82UQXpOC9JrhMJc9nNthsKtRrRFOtBb3csileb3U0
/kcjQPrSPDQphJn1tZpq0eMn5irMX9qf308Od9Jk3Z3JqeA2eJaL6070BM28uKh5
6cxvjfiwcyAx81VQgyQz2YGq/oyFN1DRkVe4tCVD9HrlXcxboxSHozUnwDKRT+JG
Hl6st+Vyz+t4AdJpqxEf9ReCviX63jKoZVWMMAbR12pzT+AXK+eW/vG5GIKFalD4
YvSOxx18psbA/wQIHNCjg78ZANgc37K74DpJWKHRs1E1KjSYfbIm1sTmsnpo7IZR
eae5Y5qWu6L50g87roAdIjIO9CVGJT00Jo88UvuUIoid3Ytc4Mkm6nKQ+tiKPmJm
LDu3v0k8XQM+lIGGWGFujisKdKL+37nHR3tu84PtZ43zL9RVEfj337feTwXNdb1F
EvWl1Si7kgQIOfH8RPnoEHwjerIKzdD9nTfoEXUyQO97sznCCFNxc6EDCx1B2Btt
59MgetkMYkolkwKQVn+2Sm3Sw8cdtBneAAOz27kJm1BUgZyqHki+X6oQn0F9EVpi
OrGaAguqyW1vKYot0cPwVAAkTNztPY+F/jWnloBZnGlpSWLX5aib31hMOTjSfCmj
kEVwW7+ssAwQXIqXc1mZJ22E+rn/m502BP9J0aflw7xjNe63TUYoawAeRaxDgoQg
Kt9YXeqlfRv+kyW1o/fJjxvzKe0sh1zo2BCyLZyCXE6b1EIx/4heHd1pPxJfvwMw
bShEwZHmSVjH1PF6mmRajjxk3rIWjCAHwHPBxq+imO5HGVZYscxOgm4Xbfmp1sgC
zg5YsIziv/Lx64m6s9B0iaGJWNP9zdCQNAskGi13DFIHXBC1vIjyEWhAeIp+jHGI
vJrg4Jx/aBLZQUV81L1NjXp4LVr+hXJ7xoAY4rxgNSu8uX6SxhKxFHXV71a7UHFj
4s3gxU0PLIp/XLWanagPJMqo7OwiD68hrePRVpL+XlBekpItXbKwn5PTnXVJs2kl
vnKGGxhFpscY/daGg9Po10o56L+hdQIY15VcZ/aXT5Q9iCv0RjAkyl5ExXpn2bF9
FDzlSvaoZr2Y5fuSSNZpqMIaILEDtHZ/U7143MQgRphnkaCdkye/BLyv5BAZpMqi
xjiaH891r7q78hsWycxte5qEgL2QoyUL6oODZj5GmP5L9H74ugVyjebyxDjZuMgH
f4ToOeoC/b4lBblFN/5tANSW/0cZx/23zhajQvabrK6CYb/9VW3DqhgtXgXTsCJP
AciIZbYGZ1+Aa8j+6XDw12kGmsp3DbE9YCjgsdbUb56p43+Jg4d3EHoXGZwjaXat
WezGPkTu9lnZSH06euucRfDYK+c0d1+tEYMk2lIMTMVCcU0RhKKA7T+Eyeasepjz
zNvYDUBR4RwxmHkLvES15pMLWOBpHulxsx0339yCCxYdLTbwjpcVSyv8sFBRt64p
/JA+G3pV6RmpSXv7EUWajwxqLH1ElJYgOHrcI2hhERTmq0OTSBVXcdzacVS153Q1
rt2af99dBwe9BXdfU2Un7gPdKx0mU5zKle/46KtReDyuXpuqZdpFQ8vGIkHYIrdl
/5MScvywIj2eHKCbfaHusCQBY+Dclz4xHuwOIZ0bmjcV8gF1zBFMtUG/94+wSe5X
zBSVOYg5etrPASfZi0wDZ05nNDzyvxHfgTLqauxhnNvAAZnOuR6GbkFyhEFUKiJ7
5FlJ8i/e6AbFPYXHoUK7wVmIfLYfQiWlPcOg2xIpfh3QyqCBlTkXCUNgOMVkbCdQ
CS9uQY6iMd0Ny24T67bJW7csp35uj6HAbLwXjx59nvS8mKClJkCxr7Y3j1Vy5ixF
XL4k0ACvN/e5mbK/biKKG7dpnsVH+QG2p+kDLCp39mCredXYUR9J/HVIvQbZTz2n
tLNpkpf37wLBxG7I1GerxJW4HYqyLwmc9U7i22fJGV5mE3IIOpPxTC4WPp4iwYY1
r7pdTv9xd98g1ktAz1jTijwAIVvAzm6JhTmmcdqgrF0GZUYEgIVFyme8K4G66SlF
T3jlDH8I5N8/dmCWZSHsyVuPWTYHa6nN+5nfKzId9rrqMvvptYvzxKiPoropjTgA
Sw8FZlaG6vTrRICQJTtiN5PuToX7co0rY+RYJeWn6sCZqBuR+XQUYfqkp6ON+Pcc
o1UuqNtTekqmonzYSzxFopvTHdtx5ykyO0qEiuqsBJeuUz5tbrORbIzSQ2/NT8q4
MDLk/3lsZeoadCdXvb6cvMEcqWCNzZfSrgvFJTYHHuMbzT/IStBeJ8Sn1G3jzche
6idsqUKTwWj4rNtn5cF9x+dQ1lDZsO/KcR3QeZXZ2muP0rOYlGwO++PjYd5m7pKB
K5fcAs/b4y7nF0ho/6eu1bVnfAQ160MTzvGdJgrK/uHWN48YyqOGjHk2+RB52EeK
lKTKhPtZwe1E6QcbbpHq6+jDaIW6FRpQ8T42K/FrbEj/uNPV4qiYHMc+iOKhuER1
gFuiqNueVtLlaet1PCYjeQoiorWpCmIK9+WXngsQafzweZ1uO3KvSvBNbQukRrzD
QnxyYNbrazKU42LYj33/PTtvspjM1JtDIFH1QGNzPraEqQuQSD7RCazp2wsjR4WV
Nn+1rxGzHQQfKAMiJsXbo2c1ntJDyWtKQ/qsZrIGIkC7u62DlqqVqOBDIa4GqL0b
8xwOmwIzSU7q0uLA2bN5sUag+sdcnA3CB0aeuDk+6kzrCQ50/DHToVuHMxZb1OnB
5U3uJ5Dkv/jbCwbLXKPV6LcOb7YpL4BozQCN7Gj8gdKUQubQpFqdnk5PBB0m4QDr
zbXW/dA05WI5UfkPtN6YCf7ihbDSI5PLz/kHyKqOj3jVXDwmGoOKZiJr+eNnVjkd
zEjeoRcIABk37TfkNCx+xiAz0fdLhMy7aHSOQXPjwia1iveaVz/T1i9XmiL8C3/c
jSy5s1MRneXs67xjr+eDFcjajWPFWX7CTeXAZgKVLkYUcrUOqxofqN7j8F8HQOQU
Y8tz1biu1JP0gXEDS4kUOLq929CM5ShxWcKN6QlJUieLwuFbxKhDxM/KT2RIIYcK
c6w5AmQ0tHAJhrlceTpSwwASqgca+ckM8r04/kViFJeNEqTh6MV4a8leZw7FYeXQ
9TJy2pDuWX1mMA3u5IHHcwU4eBA/R1yo0wxPnW73F2nKNte21T7zAT7iThJeO0eb
orYKM+Q/jS14OxKwb3EPRJ3CZXnND/bFOatSYlf1KEmWIcKvxkYm896zvZAL43xa
JUpTKOOsGdikcWdV6pB80LFg9Cv44fjUxgMNfgNMUtB7Xe4KPGeL9yHhizMCBXfI
MgXE5Or2Hi89Qoqh+8b/q6Qnd7B5tHrpTzG6AOwEBHY0Ga9T8eJqtbHStsLYEXoM
zMXHS05421+WDIdFoYBmnMzt/hr8L+98IfckrCkyGkNEFuKhcrrY6txaeFlYRMC2
lGoHTjs5mHB7nmywM72YqH4F5cmNFbVetvGMhYev4GtfnQbc+JRS9DdI+1H+McLR
9Io9yKLkvwGH0eFejoM1FoKCKIeXGHV5I+gR8EyximoJfHc05MQ+oNNkja7iAGaH
HtXkdfzziTXnYjAf321Y7xxt+JWSrPOjRjty15eLGj0LeUSyAdHvazXpaDjT/aGB
95cUiLEWOzPTAiacSl9Uc2s6dlOWv0YdI6UKYfcR4pDTb2xcNWROWMurePDeYikp
03lP70Uk+0Scb2RPOX6jdcw4z1I90cCkBCuNZ9+SqDDHbSOzwn9ZyYMzAURVm7Oo
6qksFGJSElF/MlN+6OaHBzrlgdYypjxMKGjy4jk0FakwE6bdvddqK9p4sHumuZ6L
YygLPCo5l6RpB7gLM2h91tVnt5jrRSsUBS3b+puN+aVHzZqw7ZpjqW3+m6VxpA3c
DQ56O3y5Ap+xiWlyo4tECB/jRt5GxKXCzKjV0DahM9mlEsgDuXKu1FNNQhRiETp6
1zIVc4uJmdS2BNnAkJLNMfeukPre7ackjzWoZ5m3k+/I1wvkP+oQ+ct8cCDA+HVj
h2DsW6sglA+xr0PA0eRTXa6W/MpkFc1ZnarVH1pRHoA0xhiYF/ysCEDCtZoKQJ7m
Xui8eUNun7qJk7F+Nq4AfQifBTeKuV2Ap55lK61Bdbf65lEYMhaTR62JzPWwvemr
tUUVobmccr4Pj18eZCqP+iPLK9iFJL7388jJ6Xxjm+NZWifNeOXueREwMKrT+G/Z
n6RmVxeu+xJmV+9jb1DmlSl9SYKrwFgGpAdGSwKcgfJQiosBOaZVodwyXfLl+oub
b1fHflwS/G89Z9EcGm3omY/jQxM00e2/1p/mu9i4ii4QJqGg6ANDPT3Dj7yDyRD+
LyLqzTROOnxhzqhPEfp73pfSUAvdpJ3RRf7Z7QxCJSWylSRu6jXCMtvGKI1UKGMI
P7R3OOhpoo+IqB8XSxFP/TsyqJke1lGHHwM9RcTgVpz73LgXAvuB8OlTJG29BQoa
91k45HuRfrPeQ0hP/Rg10AzB/yqgNbdx8eaJbbd2A4vmVrJOD0Xf636iYXr3gcuc
HVrqtOg1fkrT1jl7x+R5XTtZjwjiMkKpwjyFNVO2fmVzryUfurVJ6vjK7ygwVMMo
ZThjv6sFUECbwOrFLvSGICThNIeecUSX34J2fgZCS7y08xSr0QgNgJdse9nn/X2Q
P0RdhofM9bGx0ljawPIjTXzvmm7lqbfuJlCvvR5qVXO+PADiInnnS9IXltHY7ueZ
zohSw7JXdKpZdk9HZ0X4wK8whxWXi6zkt6xl07uDCrNsTnaEkBExIL/P9UasZMuw
QxpzRXNwvs8TjmHnpQoNHfMeUOdQvUI53LAm0dGko6Lgcj44k6mUW/8zuva3womr
u4caoraPlLFOFvqoGsse05p/smFohph0HqtV0EPJlFITNbPqAQgOIPQGxQUAisTu
eanBaeVp73kI+uRLiJICI6usNvgh0Qx7q3Hlt+/nI0AdRtYLk3DUtasEyOCuOTJF
0bwK5xj28RbFmhDGgrt9BT3br6QeLAL6qgYJE1/6fjdozyAdaHe0bguPImiQGGNP
VM1o0r3uhYQx5xtpweNWw+S4tKzXScs++kYOXsqVtg09KEU/eHdfPpaEBg6oQQOR
aYAOYSs8mYCBI0DUcVU5sZGOc552Gh4nkE4ZFwe6Tc7ojdyHO422AyR53yRUqa+h
4KQ1hpGW8dVvD2S2l2+2wOtTV2QlAlSJud5mC09Q3rvXB/QkgjBNZtKTcw0jFqLb
vDg7kwql7+E1w0Zrofw8rTupsr0CYVMUh3GQ5T2PhSors1srlXxJZiM/pcXa0KwH
sVunZCMyzhTgvCXmm7sNham2tTkGowDwIViUp4SwhstOudtLemQ1IrMUdlN+loiA
kSXKz5EsKXogKwAOLj/aracljMmRQlFnWUgxLvvBrVhCckEKj3NLSUIVY6bQiFZk
wugca7VRPkxMsZ918vcUE4z9dx7FNhJE4yazxnswj4dQ2HfbTQVroN3zE0O/IhG1
g5QKSowz37k350i5wwCH6rszOs7MNs9SsmDOw+MXS8Ga4ooZ1mXO2p81hqHvNRR2
cEZ6IA/tv70psdwFWeD6nq+jHPLeBjCDx0V9Co37ON6NMBbpztB8oYpjo0YQWKMD
FUUu/cRSlLFRG7lWn/LMKPUfbkm8JNBbptFUzF2mm6O9cxfGBj6ssnJIhHXiyJ73
vvL8QYHLZwSxM04tbE1oOzPVB/FNEZEmzwnccau4tdpnZlX5w7plMBru1Pci+xwd
JJjMIG9nmGE0W409ZyT96qtBt09Lqn8/PjuSyb8HQXLPKc2EEpuGKHRvQG6LIgNl
4ecpecO2Al873vFAHxoI3kZB0Ac00/4p1eyda88RIbuhemAuONd04h1LzcqgP8bM
3FZeiJ7tZYZgAx7/LgpuxvEbARwpUIkyPkadl+FkY9nVoJzO6FA1M3PqqUXVonVj
lyw8/Gknafoz76wCx2FzQIR2+VqFOkgyMhUFV9AVp8OpmmhrSDsdJ3Gfds3mYuE6
XQDPyaaL7zXfnJCWqMhJKB7gtvyaCtToqZIev10JwvXB6O/mxhxPw9me7FbB8UvN
6HJ0jKrIr7nWiByFDz9hOgnMCv6AO8R3ZjJSsxvS4VHvZ2+zt9B6MZNB/Az9VE+J
HJJPGfOWQN/+ONulDYMGCeIrnfwJ/earCXK/Cx1Q/Sg2tZtnBZSTCrFPFgBgP5Hj
B16BZYizpBIv7EdW3cydpQxsgfF1cNMA5BiYQKqmn0litjk7yVy9W5KDWd5kTzOh
pY0vAfoc98TX7tbxKRsJri96wa9bQj+/E1MF/JKcChfs1X1RsqsWu3Id8jGzg1jy
2QrNlOr2/6/BzqxcQWxCd1tsWv0pSUzC+uV1g4oWXZ/PgredeDXpdXsHMFAHBsdv
UgGGafeSFz+XzPm1gXqRkfxJI/bKyoShBMqA6HR02UFF80GYmCBBoElsvLTa7VbH
+x2x4NTSCD80ktPafyEgDh0tpTnM30NeymsCBOI4RFiaT5xEsmQ43YOMCM4Me1I4
Ug/PXZQzPtGqaL3XYqnrIxAvnRVeDabfo84dxX+Yno9TVUmDh/HkDJ9Bfu9H3rbt
RIVeboJ3R5Rw6krCfuD91WqyaTuWRQBrnzpCE2XEBCZiHQVVDGQ5Vy7HraMXdmZZ
q1HLANFNniiRgFgKwHUxKISEUrpc8z3A4MdoqM3irHbIFTnw8rLOHxMb8V+BbFPc
CBDM8HFrngFiQfyiAnsDb6tIk+UrmjFQLv9DbeJ+wsf+mbTmwLTCc4S1DFhLSEzm
AQEzqxIkwzs0XqehizuRKhkRW5g39ECfjbos+qJdl0bHRNG+D+AtqzVgV4DzkQLa
7xrGqa3m5DqqQp7f5OaAU8WjSdG0Fi6GXOZuEOo1B2e765dm8bGfyh8nRiDVkpNN
I3ASnqvsaf0HX4GyPtZesUQ29ALVV3wf95r78GAqN8sgn+utOv793g9/O0OYy7Y5
qcXLgAEFp7u9NzSSywrNjd9ypqJhAcaAZfi/XfbEjXFYcJaylhwGj7PbE8qmDG3M
SvuJd1tYDbTus3lGyIm2s1/mr6GMFgT46vMxyf15k9v7Mz+qDSA6WHBodB2jjqCm
9I6rNFExTemu6jmN2m2Nx7YYxdorFgiATNED1sf9MyG4ymg1nzB45xdjeBJkPGZo
XiKnzFb3KSR0e3Is9tycxvxx/veWgwR0EZ2hp5C9P9WSjUaZ3kbu4FEtpqRHDaj5
r2/Rje7t2gYF8wdw2pTuHmOlJMJm37L7EK93o7TAtJlEA169qCiYt1f1BmgRvwGT
GqkYGOEmcUyEE3cJlF3lk0IkYx6ojS0nf5KVYjhsxbFjIBbQF1Om6+G2FoWxUWq+
BWOy1nRdSjwUbDnBr8BWN+N/mSEMNi8rShMXMbciPiIhrEuMI1l12eMxRf7xo7rf
xMO5RkaK7d2KraYwjlwXt9jZbLTJmSjDhRYaxzPHeJUq+zOqEKdf3YW4V0V7TQGI
vHRclsBM8p7Ua2PKnsDd1ds63rZCtopnVC3Bl0Uxz8ah1HVS+Lb70HEiMwkgKjh1
SygQWULgNPQnDC6XtExbLIwVYaKMPyEfxVelDaWg2GjI/lcac5vt95mYaSHzO14J
SRmaySivdNf5MRwwWZfJDIHxb9qXgsAAAmdlQvlRci+Q4j6NuJjW87W7thUzmKbv
/4R6QEVNtLaHiM0pJpX+a4SXwwoqGE+y+1r/rcLyfxtF4ClWMswIs1gLodyfTic+
QpWKuqPUv7oko4E6UqPkFEjaN+Jjc8b+zmQJI4iW+DSMhJNldxJB4ygjDk94iHyl
Y21+iPPOzpnErZQXTsa97T4Vlw3vZdI+ClYgD0CRuv/AU5br1oLtjLsajOzEfepu
rsxRuBeSRd1mNVySTFXuliqZkGdeTg6+mRDp75y59O7qVxzU/t541JYtPSh9e/sz
EQv+H+fJ4RmoVD4cZ9V27AzbBJN/rZXN/aUOG++vaa4k+47CFpkeZ35u7omu+VUZ
bPKnNkrKmF+CtKPPqoLCuS6DQZfReP6HgpEzTq24Z+6NbVF49xxoMGvitQU/hRo4
cb948P+wGm1BHn3dcVWIWMYsg2I+tzOZ2dxAuyn1d7V0c9ur6lcxPJA3fH4aMTSN
qZLbml/B4VU83hVq2kgs6uW3R37l5qySACiFIbrhNf6RCKigYRi51rQYLCeqRYcc
QHdqK+zjxyM3pAUZ51Y3LK1g78i5HctPpconwEx2PK6Bs7gtftTIpnXx9DbWF7D8
gQNz/IvYUD3vef6fMahgjntkI10ruf3mwBZMjjb25ysgPZ5NkK2OLItpauJnaa0p
FkIp/bOUTR40ltgW5N5cT7NnEcyQZyJEUKRWCm43QJGTrWoG4CqiT7gLpwKoOWmA
lXyqej3ylyEDWzoA8ou9SqV9CAkcciG8Xv4fyroaW7rn0rz+CnIpc4CGDfk6oJGW
x9BjiYCx9LSMEw+wcENgyHDwKaQqvsYIYNjZroT6cfXsGEIEzBQMepIjOcj1jBgK
ACykpQSFcHIDdURl4NrFPii5JjyiFmOKgHjZcayoxAwn+lOPbsj0buznSrm/Fapm
IBw+plux6LHak9eC5LbBU8Uxnrv2M/EmqQbuIGVtQfyBVZlXtQ5UgbzW66TsHfPD
9lUnwY+xn82XkLdJtezWxWYagtK+ctgmko5o4UMD2Ksy/RwSfgt0cJ23DDX+3+Q/
EhA/dOSNf5WejOGkJ/Z/yQ3rLWNLMVbVr4d3KD6NX3gUPnxefOtyCdnU3FY2IHhl
wBis92rAxI/T7IaiaohfMw91voK3SoU2IfH2EaCeFU8WOFLG85q0MIIXDFKyKxet
Rfxm58zxlNopnrMvw07zTKdch2XHiThcITF7ZRt+ROEAezK98yuynP36XAPDBXrg
fpdxoVAQPsUjl7By1bWJuz84SSFZO+FhpQgSm8FcngdRjcCETYqJIBQCTonqhxaD
+dfXyJ1k5yhgoOt7Vbq1wn1fX4may2GOygHajiQzq4rXEY74OxVhw2VWfTBgFS7T
ghZLeJ9Y0D+s1Rm8bxaNM5o/9OfJRF9WN+DAqFvfwrHpXPoDDw6RXbIZUFfMvNmn
f2czHwo7Z8C3SlXy0lrH73HNN8siodR2YqgISFCgdSPGmhDxsBJ5Mxch6Ke4HuS5
YFHoJpuBvRZspBf8gjfSkUL6F99GvFvvyj2uBEyZZB64BAtrK3ccXcQvJjvLJt77
Ffge/g5ZcLBCwjThuyPGL/K8Fnlxxl6QweR29zbU3sa/O8vSguFFRxakrPUPaXor
ZDPLRGwHfF59We4napLbw00ZIP16rbca8sh/HLPKx0+b/tGmvI/RfISNSM806nZU
Gbpm1q2bxrCGsPeviE4T4kEFbLYlGcH+/MXPhckMy+nSi/ZK3ngbcjlq71QFgjUo
jidvtd8dRK/g2D4SDGfs2ZgjTVry/CDsIPLjfQkwr5x3TeGLp1agDSadNeh0IgLY
euVYv2IjRZLmQw019ishIPVEQw0qFvbRu6LOa9JlVorxO5Ve9i8oVPSIf2d/SypN
DtO2Ro4vOy/UF/dAsBL8gM/XSM27nD4yHP6yR3IryLi1casJPpe5+jsGhIM8/rVW
lKtT2EU9Vh5xUUIeCi7zLMSnnNKeFcizEREaq5l3b3vUwu3SApsMLQ3rKzr5OfmF
AMIXDv1gLQDYYnfhaKhoIsNXcWZVHgLKRKDQgIMMBRq0lUwaX6OcITjqbpKPbkXG
LHVxe8EDMfoGaRd844fezZ9DWQelzCwQQRZpDE4LwaWj5KjwGHCjKKobk8tPe2Sw
K7E0wP8t1Qb7ztLsheVk9VzDk4B+2W46yslx2XkXVPnvM3zjnhbPXJX3vikZxYGo
ofirXZaKYFvi/pOi61SIAVYQzCKfZCPXxvGVQ1NdaCJur6uy63JL0zAALDc2i8fj
ViqEExx7+u0REdQIBDo6QvmnBgCERThfr6wYvjj8hF9l06G7xLTOsniuzW2/TN7X
Ltkc01X02kTMlKfRQ2cW8AdK28tj6IvOn1NKgAfkT9J1K9HV0xYS7oZH2Kh6EYzZ
cfq3wuYdmFLBh5pfMIhY/+DRsB4zHzGmOKHURG+wi8PJu+fPbZqaZRbl5dehmCn5
wjMpgscVijR+1DBAJzieLWQm3IUKH405izM36cl4JuChdRDY2mjWgdfLn+rfy4WH
tssWwyniiegkE/GwWTXdDRoJKA/3vPdTS7z+HKIkUdSMj1PUnaT486vcxRtE4eeW
oUL3F7BnZFpe0xJ5/7dOpUqDpv1fWreIvOWy+xKuRkn2BZrTmMnG5eojK2iCZI9a
sy87fm1ep1W4+BmLIdL7GPdd7Ziw88LlO/vg7yk9mr4UKHU1Bw9+xRdsXEYEj7Zf
NOVTuGdSo8RR/qzkrtalhb2ri0bE0VPeufBRMjm6o0xb4B8MkhJ5s7zDacp5Pau1
jPE50d6zIVDbFkH7ZrxtzYdfxYXU+4FS+avFzi7xX4vWur0pmYLxvTEFPcla44r0
9K2Wit7Y/0DEOkZ+bwzO21DDTlFUPEXoSbkacaQTkBI/d0gHTUdQ+tpSDpqWKQnr
Hpu4copdaXbwzWXMQO8OqcRfMao4t2yAQZzqdnmHNItVMMy9HWA0XVIGoXZtJThv
9MB9iYNiOZOUT6qXfcoHjeGRdG9nZv6gPJAtu5XksWMSzLLA940FpKGFP601+rWD
IalnnLR5mnU8A/7OG1LFsahWGHGnkcchRxJiYip44NkzLjzwWeYMsmg3IcpE5ouP
vU2xx3Uhp9BH2l5rZw4iabpzmA3DLIKeawpHryhcv7kOhsL4gXNA6n9JwCF0Lm/N
Ew1geym/wBNMNj1PE314QcziAixKQmPAB606wxod+rUkBKPWM03sonHGKq29BR8a
/afg3tMXeq+LYx1SzDb9AOe4kH2o6NcASy6bJBLd0FWZh0xJrXHlXReKNMuZYTFu
ABVXtKFzA7gZz447DQsCkmORuMay7RacU/xuGplgxZGsmFjD/Yln9pl3mkQqzLcI
6pPLvAw0Hr0vn3kzr0IEmsCs/gXiSBysFpLAzTNQ2X5iKeuyraStNw+eo0X4RQ2A
/IICPzHfPf8MgKz+rZoQ0qsGwHrNkmzJDUlSOxYRwgJQJ3Uzd210ZiJCe/9ky5Nt
nZ5obszcOJCs+DNVYW6wseoX2wpFwlQMaHuvyz733By2zPoVXwZGdaqI3UkAtokG
TaqdxiLglJv+Rw9l2rkurw3MC5qz0SrQyHtSACkBMRYDcBbNtw1c72w5w1O3HiA4
5YosSEbuwPoNMt1OncLfSsDsfIiQzRnfap57kP+7v4ZS2s5cYtAr8gGF+ceb3sXX
7zJJgiuRZoiLmEV6B6X2lR0uGlvv2eyr9/3/L2bkxxE4+cnmjcBkITmnNbXegZjC
XZhtjS6OS8Dn4QGMUKOR2Io8lWt2qUCYre9apS6kdQdXqIGNSPNCmjcS8GmtbQ8/
Sn4jELoTrPkLGqoYr1kyj3LsKD6Uzy6ZD04LmtFQqliEuMNLHjlfOHHWM38c2BE1
iXbl37XLa/PY7sO8I7nijoFWokVnWH8BjJRSR9EsyWFR2/AUXUXIZxvsK1bCTFs0
OGc3gfUjciohbPr++wFVExdbqIPPJDAY2NPB6b5eiQJrPV/OoKzfY36AP+NyCmpy
byfAopyo314ozbrsfl/PkiZnDE6LWfxMIPrPGJq0yJSZLvLCc3RxfGkILqkireuD
qVACmdy3TrV8rHH9kHaJbXgYo4vHEYTkGMNqzQlqssjtZzmzPm30NtKSH78YAcPR
v1RTNsWID+sHjKu9wO7Ew6XMTAvPg+7itgV+1tmJl6sooUaVAmLDgov734ploarl
602yc+M3OvqOZjvKiwcF6feEYhRhd35R71kil3ha2UCuA/SI3Xn0xL+A117wpUyk
i897HVncaMOEx0oZGV8M6vHXmWohNW9VLAhjAIkN55qSP1VvRqb06pjvv4Ju0tBj
K7uKC+8tmsEY1gZkbYhiqSdQ3JQfn2oR3jvAwygp4oarJzK/l6OMYhbC1plYe75e
quSADBQnwxo3nsUSO7J2+M0ciu9WdwG3/kaOpaLOh8pgbL0O/q1FYOZ3v2B4/FSj
I//lu2uPUQMNnsjjnCvWeyhI1n2/dbN6bfkACym4BI5WDzRwMdkzUUeEFsJTdtY+
u33GqQW+YdU+zU9kuzncRhnZzVVqZz4x0jw0et43IYAFKTdke8do0VIH1UwUKhsx
PVUk3ZAwtcOhtnjXotnvctywis5GymimLuR3cdC9YFbltlMVnVPu66Ro8Ng8SIV0
rvBSBtHG6duyNSuyRQYclJrkwOvVgAroqxUFIqve6ZKLK6MD5on5Vwsfy2AkYz0x
E5RC/Isb1+guaT3AjrESvKf0dZBYNzNQqarM20k6VfeRxUtroVutIWE1h3+JZszb
+KvHDHIOj7HjBy4ZMKGX3EszHtU9+Y6eT2DvUini1L2j6/0Y7AmCFj6o5OY/dr+H
94PpKESdqLQrISWX9JOGQbthjz2slYcrtsUG/O5Wfmx1+MH2hGzZP6xuBp4PHB2e
HwXrJzdxyX3cLVf8IrJNeFCLjEEULipNIBJWfqRi4QTw/3L9rObo3KQREm744UHJ
Sgw0aPwy0K8cbrISNnz0qnVjzG7hFSxH6bec+rkOnXClXM8UAlnBs7BtRHoY94Ql
aIY9OaAIY3x32WeLbhCjPM4xwE4zQqUNudEaZp7WqFRsa6Yo9xuzMp50667yEQK5
QlBquzkPaYh1p7na2dgCH5KqvOgj9lSdO9JIyXF7VzYjNZA3X2ryOWnA0PpDyl1X
uPPbB8RJ4aTYShcNfIYku2y0F7e2ZmGklwZY2l4Ca5oJzCWNkLhrdx4G/oo+6xyH
Jk5BwqM1kVYsDgt3NdxvcB9PSFOEuFhBepye044vYq85322WOIdXt0hcxSVdXLRb
/32hPAKJqF1SggVIUh3Upvb0ReIprbLJeQfvPJ/QJGjTFvt6XfWw86Sk+2xP8yPm
SIH5VNP3Is0L3nAxiphvc8ZllxHxzarIkpWWqjLpTNgsijqu647EUO4ZliAMtcGN
1AFRDTgQFYfgi9sTF6B8yT4aeQ29NeXUKDT2pT5VPh+9gMqxx7KQQCqRpDP02sCa
8xVxlhoXOBNnkpAaeNKbwTkWBFfwv7cvVf2+Q6b7c4ersZdoK/RTIapYkTbu32Uu
roL69v1efKYj/zLYUIKzx1i1lMC75/8vHjxqwGrjHzHjAexrL9wx4C0bDw1HZn4r
nddsvFuqN+igRIk/p8wDOwN4kNEbX6EmYbLAZUz9irIbNGEHddc2Swk9/9hlQbV7
1VzmN6CFmkwNmoMXbUkxNd1zTO2wv9iyek34avGRoV0KG4YMs4TzFmX5Mssj25lx
oreWgeYyWn+8SEPC0VnfcdyNH5Eh8TW25sO13ipsMRbQRsrm8nmulgfcTUxAApAo
9qcaK+bGI7MqeMxnld9DtEA0vXhd3nNUeRBGyM+HN3xDoOuiseY5yC9z+08WQ2Ln
c89SPPKI6pIRqhUZN+h0CnhkUXTAIH0xoU+aEvJRNXWFI2DXOPjEYBHSQHAlrQXa
PwcPix44hxKB9kCMd8p8FQ7C6j4iU8YPrHONz5aR/CxD3xVG18KWrXtGmbRL4OB8
xZ9Z12yj2UfJv46AAOCKG6Yb95KmJVtVWqhjwMAC0eYJZ7kwS9qfMxPtbn7ovqAV
V+vGo64xbfHcsqQNSLXVpRikMO6Ko8uD8WgtR4Zyh+TO5ADE5Vw6flqBwVplppcu
JKZBcysEIhYHZr0MymTXDbnPRRptOEQt30xSpbtX/TkF5hzf3adgmvvDDMZZKuKb
azl82LhKbhYxqiZXNK4kU7ei8bakVBL79gl9JhTd5D/LRHuHGBObkMz0vmys+7+d
auPsItm0eznFzko8KJxNhaKBvIFvoHOEAmhTmxFwzzg0NWGVLuqg87le7sq0kGyi
rxWdRZ7RIImcXWAa5NXcrbXUsOvCPuVKUQA7UeT9ZAYYM4m5MkswsybYOVpGni7j
0ZqFIekyUtOi1kxVDK6BtT9wyDy6o79pra5WoatZt2nL/uDtER11tTpq4z2EVfc/
dUGUvmqkpElm8gMBRluH/I3Npj0rzPRHSaqm9BY2owqmbB0aHZto5Da54PnXaHQO
zXePE60ewPA5HbRgY5EPm9ckbPAkMv+74NacFu5nwY3fDJRgu4PRVrdQviZuCvKU
8TVtWHLXVFnLMgFMjRgvnxfGMAfeMM6HOKUO5ABcDVrLZdVlzWrfJqyg4mXJdX62
paSgxPl6xrU/hHOYUjJMydqiRzxiPD5CZHvolAi0sEe5XpB5bXnxxTzr7qagDaeV
uO9tV5eoFIzKWQBZ7MA2jf6pGVuvkRE69gHmcOJZbvYeKWLD0QoGqW8AswQtkJuH
TjXv4KiStDW9J6l9t/g/ugymYBKalxqHNjnzS0tiSzVRLKEDu4/yOvEQ3Sp7qY33
TlemhP6202kXfcfoLLrP51Hy9H72RM651v09caeZXA592Vuw24fKdRHGE8rsS3nO
xWYAXosqnomqFA81KXIIAOR0udpKjF+6qK8SS3aa6tFykleViyjNqi4iGYNkdtiF
8iqDuZpu/d5aBAmWSzyzyuQ+vwptbDfc2CIRmMDrWSzYuLL00htQVUxGb7TuqSOT
o+d8sV3kSQ7IQuD5ylUkzHIRSG7lamuexPdqSdMpbXBMn1as8RDnVMMuWf2kasBD
b5xIbJnZjk+O7hc0veWULsggArUXFtYc/h2qkt+QpjwqEpMOC1Rv3s6yxfCxUwPB
qmkGMO1Spyolw6Nk9wHV/ixP41xRoZEyg4q259I3C3SnZmwDjpTrYRmqCOMI1qsZ
lFmz0+yyOjXyGx5nSYm0zZly5D6ju/snyUpvMkAGTTwR/xVbkwAFYshu6v81oCXt
e0XgYLUIfVuBqaMON/7hW7mCIUed6FSBNkZkpimpT23M4R6Zk2nnNf6mnWy59MPY
E1uefiaZNb5DOSof2WTFt7S+v3xj8eOyUOo086jCrxcX8DM/WmY+ZifNK4r9olSa
DF2tr82Oe5ds0rOxGDa2wJDKfpE/MWPIXAVapqiseWPgoQJ/n/oCy/W8tDvlNsi7
C9/aLMy0Tk8TusGIcAaxnJm4Sz6L4pmJGAA14I88RTkzTohyg0EWGzrmjhuMk10a
NnDy1WIBcKyhxaQvcz9gQX5gQENsQcWMwlNRD2ahQ3jDg4MqjfkLsqwS5NzRXLp9
+8xNQcXdtJEubDCtZJrr/HFN/0pHdzqe0KMwObRlwmtK0t0jOB1rpAXloguEYwif
GeZJJlVT92UUuXID1uhNOeVztVj0hOFSxB+RfMfxJhVvy8QzzlBvez91QwuZath2
NeE36XhPTrwn6R4xSuLUNp1HgYurbJ8n0Vo68dFW11fstsWiDutO31sVgD5fddL+
GFQipTRhw2+cugSFQFT8frrpq9gE+WLSYMtluetahnSqYJJeMz+Wac+DAI0s4nbS
jnnIHThyt4G5a4Wh7kIUtoCEADNja+daXeQM3sbUrluP6CXJAQKbtglxBgRmyaDR
MM63C6NyIOz50pgpX3DiX3uf6lE1+kj+uqQx4XaHvTdSxSC1yHT2jzA2YC4cJt5+
Si1RZrU2IA6SgC5zlqKgrjiYoIg8CFMky44Jhl529mRhszGbVdq9+axxhiHplr0D
Qvy0RabUj6RLa14SLJDm+q6ssQ3XFuc8JDZbMqI9Mpz2vzFPt4b3tQCPV7+jQwAx
eoPqYwah4rI8WPi2/ebO8yS+GnQMaGDTUkksacqKgBrxNOuypDDrpyBYATdZf7+D
+dP8S0NRzPQCVORbY7WZDsThF0Zdzlmc1oEq41wZ5oTT7Y5KA21Pd/5cGbe2c7Dl
zBRgFWDXBxyIBSfrdGapzBS9srS4UwpvVy8fn38pnltBLc6mTvkkrn7qUyQjg1u2
gPypLaBhxwZKdeloiq7Jc4dtkIRTGdgAzTyBuZhrwlqM1gFOehYpwOife8Lsnd/3
nygZqUhmj+3hPE26iivD0voxmgCa/+bRr9UZ9nl9nY9LGZ6N7tbf1RLZzt6EFqfH
+7rJsFExata0oZKpKcCCBArTr/6zTDXHjFCtFEIiuy4odcdkVl2VjKkLpy5/EyQ1
ZyVBxKnx5jEbCG2fyP13YJ/DWdgO6t7XZP2X35gNBcn1KHBuFTwDAwKdVplE7Y2Q
vPLkh6QYl329WTNjA8WMInFk6RYw41+uA1JjWlyONFfZNW7MwRHHtZx4AdN6K5V0
FdGf5iNxIwWKhrmhk8F5av3a2zRFk5ONQImmpl1rr+34Z9xWwGXs37oY+kOHEOAY
7uqRIYrzPy3wTESbTTfYZTimd6xEMPfWKMfurk5Bqgw+CEtZP5E9hzEK1G6+sl2i
LlDq7YB9l773dc+CoHcRzjaTUtSQDWXxofQQq8dIo/nVwKfnSy7LnPBW4kB9j8UK
Pi9Lxj2rAb+rqawUU7/+E0Ei5dR3P9QJ3HthC8hkE+fr85ruwCeHBMS7hYfwfsxJ
absuXcaH3TwUD5qMcOXFKCukAguqGXtduDIjOhjIxGS8hd76e+za6nK/Mas/hP5D
DBhCjXD3ilfD6pIm8ETBIa6NkIkkMy5WN1ksF7hH779vhDdb65jQ9NaVXLc78EH3
Grjwfo+53uN6wvDqY+rncpzLagJl0LePX4iRc5Gtsu7zsYLIL/eisoZ3zbcKo4k+
6wWBei1lptv38sxiHCvXLTPPgF5Wf6qCU6Cs0lvOVN95HZFAWH0Nw9+sMk9W3Jga
UClXr/bv/GDd2ZQmnMGarmWWtokxik+/Vy69EIv3HHHWiEZZpfW+zKz9bQIxV0Jh
TBXesJRyjHXhk6Qho5zZl4YtLjq+q1yimP8WX/SPURoYPZGVqRbrJgHl65VgVI34
HjvyNR/bNA9sziN4hEQsL3uEMaY5u12r9AkPj8c2+xncEOXMSKHahWQk91TgNSCh
y9kLMH4TYvU0HexnTLNTMvgpN4PR6he+xXsB0jVasPDU8klvFBEvH5fUqJZO+mai
6LkgBZM5XTLf8htT3bWJMuxH2gf+pc6O+fvKd3QhVtiuLj5yf7uvy6lPtVIVi7LN
j1CRsiEmRgGnnLbK9qLr6qNp0/RQINSNxNTBalEPNNDrs7pmkMhpjy0sOXrrj+4V
wlDxQ/k/9798qXWDI7vZHH+gOJoAeJElahpC9GC+0rBxLCjjAGmuchX5k4blnl48
5RIDr1ewqvz8Qvt9/nKIGSoTHfbBmJ0lo57+ihThSFYY0XtI6Z4jEW+0Fo+cM7qE
7IZtMiNSPz7IElVU9EcjsJAdISV5lRjiShoZz4oObHovVazk8B30zXqlczV6ZGLP
sy/MVKkbn6Xsq1RmYXY5I4AHQbBDWaOZZVWy7ZejkfAzZYcrg1WtuabCflicsNiJ
bj7xV1QWb9qZeAxzS+omUR+5s2o6SkhJQ6Xf+jSkYZ6YHudSxTNeNuYmGdjwYJfT
P3+PHXlxG5e0zY9wp81n+chI3F73h+8U3iDfA419pRBtUI0ZFskhhjGvnoCSwNK4
0Ie74XkO/SImQg/kYCDSlK5cpvQhR37y//2vU+RKw7NA+NB0OV4FGB+tP4HbK3/n
pEl9eOoO+v0+5oSL6AKa0jSsbvAgNOBwA1xjo0rqIyxRS7pKyIoeitn8AGlJAceH
+cUYbwmoXNhZuvva3SjEQQ+Tme+jufEXrb59VJOrtMHryPr9Miy8aNdOTHovTptR
22z4ErGVGlkU3CKxh9awzZ9/Gb00Zd0cf11q1l/p5JiWVwKBdSa6x1uDM/pDp3xo
YGyPxjlk7yvkXnN+j3FaQApTz7DQytg4nuUDFfcQWz/vQMQ3hCGSPR7dkul6kXp/
s13LBpMXUX5+SHJwNWnU0NvLMDZcab/wVnqGs5vyoU5hmNnp2pihgvqHUub48pCb
qNsxIImfMohp7Rc4m88PZUZT1kOpm4vvjczZVqE+ZySUmIr1NiuumwQupblzHMRg
ductzigPqR17Ak27ORFdQT519a4wkh94ZZYb3vsq2XtlhkjNaNq0hN2WcaI5WFtL
nOVnDMTy5fAKVhA6jF8ycE0l18yDaGw7ZvQ9fnOk2YGZjw0GCthnYkNo6WUP3xNp
OhZSPgCI0HaM9itIWFi0Dcl8SnOeeW1DNQkE/IpJpAvSGc3QNLDFp0ea3bCQ2Acf
HwSUd5pTBlpoS5VZPkZ/lhJkXZP+RWJrTKUwa5yMsWpY0thI/Ne6WHGUZLpA6dtm
wkvTD9m0IhceRNEmMZuJdiGycF6vaKvLFrraGdA2gvjPJ1bXpF0gCZAKhsYhn62h
j8wg1pHILs8YYu1kYaoXMi/Gaubo4dSKeEMtbx87f8p8DpWaA1Y/N6oscDYnNPGa
3CP7rmAOmizLFRseVMlO70/VwnH/bQGcFlZFgs9kHynrSIcgEaOit1Ggnb1MgCcC
2A6ljO2qimRSEjA5PL/GeRnogQDn4Jg8P1oKAhzpQqrCJatSC8Oc5nPsYDE8ZyyH
gqagQ7jcTO9wNv5Z+T/Vnu7CsE7J6eGmLI/lFJ/5Obvn36MO/oiDPehO6XxUT0au
vR2u2yzJrkOZu+pqeFg+FYl7EPEhwSZR6iu+AESyZm+CmpakAc0k6NG9+D8++JJt
waaL0zZPBJypTacgV16RYQxZMBaEYq7p2v5vo9DAQStZ9i+UXfLhYRueLXdH+rui
s2vto+NBK0tuCJHbGiF7rNjQhPX6+9r/Auk0sFpbOtGfEQeelvxi9ZiYFTxtVhMD
4M0p4r4+UzNxNPN6jZq7ynd46SWwqtW1QLvc/o34wDzbqXvJ0aM8tvTVSTAsTF05
hwnBT3mGKz0LE+/zto2+PsKlucGHamtMaqoh9+5RDb0X3W+G4X+b67aPJv/ci40d
QecuQ+dTbInfCNnY+bXulvd1wlQWa3r1Qg0+1eHUybypvORuUHCILJ7b6aSD2PiN
uydiUQkdcL49FV00rLgHlUjjDbtVM8xLKhPspeFgM3HbiwKdjk/WMQZdZaErlCNx
FwOv8Senu9R53urH0DTAl5XYnxmoJmXrorPW7WZ/mHTZ6QTm4v5M6vGYAg+En3TE
3S8NnnenfO2BiLvA/iVuzXJlfHGTqxgh9gpJp3Pn8XxjOti3Lrys9n7vW+XpEMjf
Sq8SygapmzBsEhmHwanLdgC2eQsxHXVHqa65ZlC3KoWt9REkWKH9ZY92jTniaTEd
itxtYbjg29LIwgMnZQAZB0bUxYVgIgl/h4ZdnkRYSplpF2G+R27+Cg0zbAR2ZiKr
Wzo9DDFTwa4kaONyfKzSMGctQul/eDWd+8Xa366iil/eLiloKDtB+Njn9q6P2eJi
hoQne9dJprsy9ZuXwRspPmAOisGWCNYfKxELTspFkyoCfiB893TKx4HqDc6fYYan
vG8pFbS4YR+8VH3HgTfZ057l+EAcHvRfX5aIZBvKy3d3Yvv6lQdKHU8e+J8NIunx
zFFkl4sbb8UxOb/xmgWuJDvkYWMAGj6A8L/cYOJTw5mX1xOVJJi0WIYR+SIMH9GB
48LVuOsyTctFFDyM4pZHwjRIBaDRHqS6g926XT71Ceqtka0IxpF6T39Us9O97kA+
vOhskF4RfrdJyq9yMEQjyKy0+twuSy+M4NLFKbUCHtinGzvih5ynu03v5AejEd37
DummCbF+lSGuTtjT05MfxgkxDAq+0zcrMhLo2XBWByLyRpTz52kdBPZejbhJxlWd
AGEEhB6d0P1fM5QhVK65Q0rYgEYB4h4FuDNK4p7v/266ponLo3vLRLAYsAqVZcsh
dRTpjk0Jpnn0mFG+49+/Db3bIUpjr0HhP+uWEK0KZeM7RpOV3wUT+TDdcb7r8lWw
6jnoHvATpY5Z1wir7XoZiDlkOjdnGonc38UtiQJHCAVX/Qd25Us2oJDytSOBraKZ
6+sMHHSWfSjhMP1ncyDQg7s9rH/TtjMICrNUuPqGRX0YRL/xJl4IB5N//LwIZFA6
XdTAFJj/t8YSfPbCK+wcFl/eVNOmRO66Ex/mC28ILotR5bcqivnzXOqvOXYeqkOy
s9j6bma2NQq5OV1KmvCc76fauNL8KSxX4Rs0E4Y5mOIx6Fcf8SGrA5HE6mpfySR2
n6gJIHctVxSQCVyq66vgAHEycjpsG6Hrf6z8nUXQSuRpG7ivJSrOCdEz6QEtaGd7
9WQHASIWgPORgagoV8mP2hfU43MHySnujpZiEgty18AEicJ9l4eaVtEmT6/U8kGJ
TyRtKcai/NQQx3IzlzKmibMpn6WkY9VoLlIWcH3WeyTjyLPWhbhy4xRM942JnC+y
DDMS6bCRPxHKm1fxsh9EqVORfvlLg4grXWPoEgw3HlK3gaHKNSEDes+R3S0GBpLu
2gw7pDdsEwLuOwt+QtnKrxNfMnkm61xoLc1t/h/K0jXipA+5+MFpgzBu++W/MzVj
QPl1MXHVmTKf5lI9IfYFQWI4xarNEcbvnOq3O3bszdWsGOEloMct6HSJd37QaGM3
ow3oBOXTZZB4RnE9eGrMMIYFBVRGPKViozZQPBMxYze+O3jW90L6EA9gQIm8th48
LE2jNMYl1UWS0XkzzF0MFBIyRJMzhPFaCSQduSDriysd4RCk0VF02K6HSAcdGwxw
b5JRFyEtFNrn6ioMOVp55ANe+Nkq6A1hRALRohgEv4PSfNWJzksCKxWRb1q65E6g
alvh3jOuARDoE8joj5+QnMLeckDAV6mriPhoEbbv7P69AkB2IsE29gptPOH09X9V
Ws9wKeEl6fowUr59CbHIOu8k/EEg+xotxFTOohuSD84yO43Qcw/XRjpHBBsLzbbu
WyaIzFZX+J5itW8Ei+C5cu3x+/HuDfTCNm3EIG5VSYccrJLxFbdjsMEHG16vEIhd
pppaXuiz2WngUJ5FdtQGWYVpURTLHYwovDx7p6Sq8ZvDcPlBRIT1z3D56NjDbVUz
3bCsYyri7lQegmrMcgZvz6X5hHkW5/U8irPMRELwX3HmALkSt1bL/MnO5McSeHCx
ubo8F6vm2Es2upEgl2W1KTLKBCytG2etWhTqGxBjYUc5Zeebrr3p1gGfAgpKxTuu
XhPApaurhvc+fyggRAHjnrrNhQHUrCfXCFF9VRTcDV6Yd0wKNxx/KMHjMTCdj/vE
MQuI/0RJyXnSK5w+oXiui+sxAvYUr+TF3iuxUvTvXPZW3QVsTjyXeBxldoMHsBEc
Twi7VIesNP5EsPq0unB3bsLRuXQlQXyF9knsMiKK3yF/OKnG7RDaSpn5YgTLKF/6
LUxv1OMrnScOBw2sFXeEKXrX5bwvCDzAuUJ5221/PIXpKFqioEUEuNzu7LitkSfV
Tko/4y9FvvdFo13UXFzmgR4gBO4lq3x/6sGqtTpUcrFUCo3pP2/bHKhJUdIzFqSS
a8JOusZcg7rn6F334RIulf3NS7jEQMZUjMZ28EL0LtwN3YuYSSWc/l9j7rDwbINZ
B0cIV+T6OMZo8drNLu3U211SRL1EyJz2jgFQFR7AsUi4Sc+2O3TnDnkqA+R5d4SC
CMT2/BOw1g7y0JEJ6lV1NJWlinwUU8V9CpiK+mQ9gxVRLJBvs3xdl9+q5gZBSsOv
c1JIGnKLYIZ3NeqSd7k28WSIDzm80hHiwdvzCdmbAEOFClnWGedb8TBwbbssuoXv
CIwEGiKc6FM5RBjTh/xjLeR43auu98SDqXDdrl7NhRnXVDul6ClIZPgMCrTnjfeD
LnfdaV4Vsenhnf34a9l/5R9owhwqJALHyGMiLGEiVaC+Bu7LCcE2SsmPvQrwYplp
0w3LVAP3EZngrkMShWxWUXTL6zvRrD3HuhB6tFLAHYPYVcw1iI93uoam+nmy9LBf
u5blJEV+u2Ex6RcoGi5kW4wVlGi9lKKaehzTp3y3Na0n9lIEcMTRvjRJjx0ynk94
2oDw1HSnwWk22nGZzine7zVPR1HIdG16A57srnUn/a6ABZ0g783PjjBXwXZ1rOyt
34Qff85lC+qI4p9t2ymBchrgUD0USw7s1JwuPC6zB07OdkaOZQcHHXkpdWpLHJTX
mNtoh8qoIbK0ssNTUOudiDNiEPVhRp/HOljdXAlRTKw+awUvRAa6YHRGbgDFEnf3
7pmLn4jX3u/+bSlOpt14xDgLsMks0y6IQV4gjUlIdYG5EUa7XPafGElM02ljj2At
w6fz6mU6f/zH786fTd2H6xaHou6+QzHUMR77mawhcDYVSe7xgPIwJCnXvPTkUVBd
FJB7F7ZM/AuXSn5s60Qgnu5+n95hO0XoNjuf3/0nH0ySxQdSqxZsZ4EyFTVd3GS9
pdV3kXJbZYn5mbxRCKVjpo6wfMmnL9f0SnQ0NrdpjwyVEDajf5LdrPfcM2n+4W8q
S1mBaU+PyE2CBv4a8xWzrN+5DZrBEQXkWshSps0AJfw8VMxcXnriQqjJ2PuhH0Nd
uqoCsQmpbLLDof5azlA/fc/IeahxUSE4qwGdym6Niw1xkaEXSwSF1f6dXrg7AiOt
aMzrPHz/t7eduAzpp6W8wZ3T7XD5D58heatQ6SrTKS39paJ/oWV1bKdHCJKzJOB5
AvJhEQMtGlENvZyvFU3ldjTCBVMLLPPVE41zxwddPI55enC1Qz6fKBh+pVsSH25t
EG3K2qXjOedX/xzH9W4tS7ih2DrJh5nKSq/suizbD3kc7dyqneT/8o+IJ9R38jf5
bdnom82ORZ/AoPZ5WMRWHxP/EB6af3AKZVa0DLr/04mVRw9j1WeXxn8QggBr+YKw
hZEiULv4NiDNHsS6M9CaPv1cZB4NuWOJ9A1R+wE3tuhIVWcOVzzAFGLF+H+nCLp8
HH33y85VMK3nu/rnejhD7n/oPE6di18BALO8thZf3e5ZRzmEQn4tfUgTHFmXNqoW
0stMr+T2xwOAcpf13uPtIyoRFL389pbOysC1Oav4fm8/8MqcCeSGIe7m9ONheT5G
A44W5vbMTsK8W5mPRLcP2ObdOD64ls0Tk5Y5k05rFOMfbThr5EAGUd4RjYimNymM
KF+qPTRJuv+F3CVTstCyb5jcC3+37wUEatAUdwxh+eLBdvr8pFk+dHJFnZ/GAGoj
Kj01PcNAEePf0rP3OcFpyPjGcW/uTcxZzpA4t+WNTB3OxkAdJsaoZ0fJPaMJA+Fm
9pO14PLzeNNHhe61bOC2yY00nsuEtGFOlTolX5OSzhp352WO2wt9AcDBXAglm2Fc
mOPgW9ai65R9UnuDvhiY7KZKf/BvL55l0BjhaPtR5PcJUOcc/mBisLPUuJ4Md0ON
ZaMPXLmE4aF2AY5KGZDTPzEdhfJPoMehB1SKa8cPPjkoA/fGHabWOj1sH+r29Ure
ql7vbahSzqGSQaAr/1l7Pm0ohRLQZl3dZx1r0oblCYkqioQbk2qb6hkAlaUjIsiY
/uIKoZFtqvrtYW3BoZGd12K/Jy9pQZAm7jpasz7whEErLyMJuKAkb9sCsAH+SWMx
ZzvKv56HqUJPXmqIV6sK9LQWwBJYc2Yi2brh27hNmC0eK4AsQZnqGreeAcEiHKVR
TRmhcSnJUEM3XJX9pm/wALGlh9V8YBwY9L0BjBAEZo2ltDL+uTQbVxVPPBTfBnXg
uG69fG3gP37IX5gTPpcjM3cb5Hxj/2i1Qyg7z01dTpoXiKXC3iMGd9lN2NSR8exz
YvFi/Yc7ShrJrzuyheckg83UjZ/FO3N8xKvf748TaY1sDKtPrXOmloSNC+jEjkfG
V/eV0Vj+oITJ5tj9wmANcMX1sghM3hKSgxmjnyGWBdit70lJi1AGg92ZoYAKAIAe
aL/4D8WhcP//B9qr84W2+VTgclyxdrykdZKxGqbE2ainP562nkj875ShwZ99jbtG
m2+J9BH4xQt2zN8bkAFJw7CK4oIb0RSVYTjrq1VmGZ5SMNQriIdkqKxZNeNsdZKy
krTpIq1cLUz6njXUhXL5q6fOB/P0g0zP5NOlGLEYIr5vM6vBksCAHKi0U+4L2wQx
KVOtPVKqJU3/OrwdMqTCQ6BYrzA6l0EUg7SnA961gDOuw/KDTSTxllrW8NPNeh/q
nXJYEfV7w4f5amNikj9V848SxchTRHoLUP+5Jgk7WVyUGsrzXp31H0aM2Iqd5/m/
ElUDEUnF2a1I1p9wF1jHA8cQ6u1KiAhyw5ofOTHesqMJQyBZvKjkvv60Z1ZF+uZI
A+BMZO68wfE7VRp9uWa8/doyZ+Rn7suwlKv4DOohI+JeMvGKdSL7eiTnjzYq+Kjt
0S3UnMYPho493phOHRr5CT7lP8hgFZQGcFbc5zyEc3KDT5heE8DZbrgZafmfakON
StMMK0JOWx1v/LWOBL8BfwdLYwfBHiEvA+Nu04JQRjjvg3vhU3D/5IXqMaBwVg9D
Axkw5JnFLtUwTQNc6o1eV3pVUczRSciI+DgZqR+Ua9JDyfydQ8wQj9MH+WRngQ8L
2KyepaK+JxD4NG6zBVk2LPjzABe+pC4dunfhqPVMP2Bp7+9Po5Pdwiu1QGXZzXM7
ghiesPfpXcT6oDD4T1jli++JMmv3Gadpbirhchi8cCANrU5DgOfbAIYyyrtYOMw4
5L1ckwDZy4mHZ/iWAPsnpKg+wPucT3+CLvfLIwqJT5gZrIX/irBIxyJMZH+kBdx/
oDylbro7T3BQ/YvEEKj+v7FizKpwHqhmJ4aFT6xw7XQV9FTqK3U5SZZzci+X+JJp
KNxS1hhMUJRWlNvKEOObaW9eTSoyUQAOuD7SJQO8q+KWD2puCtrEjDhhMhOdWFIR
AtvcKOoBDWavZlDZY+aUa0MyhDXWfZJ5ZsYcZd3aB92Qlj8ta1SsSf9t0+FeQUrQ
kvSv9iBbEudyOnfIEsMqa6fuYiCIMqbWLeRxLIOsxtRXQm+AGhFQU8kDkWkPXBSu
eUQPdQHtK2PWlKqusvDwxMhL9TYSDWGrB7Q23zwVo49P3lFdla/f4pqLSvDgfg2B
BdWQkL5mGNCBmrOrX26h4BlYRxWjJfu7+Fdl+HCFSdWApwqnfwl0AAjhLCHh4tUk
ZahOGud0boIyN7DxQIQKyRqK/CP8W2vAJ+ncv3hSL/nNhhU7SDftNOnMtvPHxWjP
+GhIBHQHCuvsn//+24WAR+kZW+8IRh75vhh9RkLjM7GmHNtz7jQ+ZK0VguTrOqrk
yapEiyHVWjWKLwNIy2xUPqFuscPysrSyfs4Pc1XmARC4CD10EDinlQ/iO+y4Sx2j
jrIZChruBQdoLYBcfkYJGn1GfZlJP0eyjpZn80JlpZUsoDoGigLzDu+mHgdrWtOp
oALbI0Ao0b3bWL8RA0iCmSuJL0RPEiyVzCUrW0bk6mE2KFWcrUnJarfdgCI3Fr0p
xMYHrhoBgx7fps0Y2V7h/TQ96dVNrSYgA8/x4GefxuHbl11v34gv58UscC+UcXNg
vRZSdLMI5iAtMs9XyplVGlwaZ6Kpu0/AWjxY+cH8MOnYyY/ixXSflVd4A+/YUPLr
QsE6xIv/NTqecK+kroZQHl7qcwm1wbfWXDZkvMu7dGWCreXtPDtuDvCgzrA8B4et
7ufKF08PHh4OTQ26VA0oj6D3+1gETnUn/m+zDE35AgKAy9ufconAzUnnjEKh2KVD
MeqzDhIC/kdqaDxCTWymXwonnnBDepSwxUccdFp7fpxSSvnmzEcTpnwd7ttBCPO8
7VmExrAEnkbipqTGS/DeXns9Br637KcYqVhJCR9cHna8jK7xxnvqq08HwnRPvc/U
KGHIMWOhJqHd+IpzKSHcQHE/kCoCyR+RESuEa4TLjWt3pvp1HmIxGocaesuVhvRz
YZvQM3sBT7yNJn4HELruoiTFYh02Qql7P3TI581DeQ2GUhnbBpV2CQL3gC5zeC7d
XjDuMzl5/Dq8ZcqL/YMCydT/aJeCWJE5sdq7H44di2b740i3LUw/yeEjIYYENIly
KaEce65VfUhgOk1xKuNJsQZ8A00RdcXN31YIs9SBsUiswCU7TzrSQcLtkc/qq+vo
2trxFM/6420yMrk+jqXAav416mDkqayIhnU35srt7quPZpkqcOiEOOziz4I5xPel
a0bbxTNhL16YBOy5ZdgZN8wdeLL5jEifRxsvFqEHo34zLtHEowMCvdJZdXkA5MFU
FIbpEgyU66tyVNBT9ePTf3hXezYsmXM6vZF5ESl/bbdNISLuSxElffrmWzS5VePm
WouyY5+dDq6ZB+3krwabqiLr4Pey5DcWzPis7wGBM8YodMujv2C+RChTcg5XOgp/
1w6Ado6tgzDKjCqG2zKBmThvlYzgRGhEU07xcyg+tKMnZ2hihuy8FX6Fhn5QWrUX
Yfx5noEel9QOtVWOT1F1AVKif5tjmAcnbLKezTWo07/7gyrjpxXqXA1OsW/XQHaN
a5VegFqVUdQmloLI0tBi/ssyJjqEEMSiSmYCVoSkSxCCp02x7T6DMxdSNSYePA+Q
LrlxbQLkEL0G2p9RJzb19ogn3crDNwUOsUvpJ5cfuUxCt4dV9MGcGGbTJPlnldc1
JCISPJa0uBjL67sHmSxwOLFyd2Vv/UHBS/V7FT0BxHyOLjdkXaQ241ptCf2GJ5+N
gwCpvEe4HZIV1qhxQ2W5ZAt1R1oGc5tMfy9VpU6x46JtLYzXsWactt2ryoA5s0Ce
SVETEJEZvnYWvd7j+di8e5BjpC9eTIYoeCHvvl76hcwoNy891/GBuAtDU43Rka0+
v98JAXXsc7k1rJS1obG567Uiounwf3NqIjrZmopN1M3QFa8nqEsZ6iEN9NcZVeV9
F5Df7rfvHvs4E07QeKgxkW+u+4+2v4KyPwJV0GeTaJWve8MV8NU1VG26wO+qS9cU
XYAM4qaJkupzKhPjjNZLegBxBKSuK/0rBi6wrG2iwrl+u7aWTT7qttL8oA9x9nHX
MhFkPkpYi1mR1WxDXQsPnhdCkUME9fqqjrUt/aCHFeH+mwOxmPbW1Toy/U25xCV+
FtYG2rFkjme6Mw9Ma5rl2WZt9w/NTkhjT6zfxEeIY8JF9Rymm8NrlvBNvYpVbsxF
TxxD7kH2sH4XmIfKqEh/E2H+enPBCE9aWzyKcR0RR2k4vmiWemT+KCJy6V9dY9TF
QDz6Lo3BgYSvYpwXsg63EkGi4liiyN2Rf7h/dvkUF02ytNajAjpzF8wevec2wpzG
1pW0q8wrQQMv4Q6dPCIMNcvy5e/6ph6IgbxqnJxHRJ39aeg0DX3E3oGCdvrymckC
K+i6+RvWiX8JSkk/bEULvxEQv2Vw10dnlyp/TLbrMvCk3mGImhyTw4RLjU9Ix/Kw
xPZ0eZHLOm6DzfuezuqQYK1agnSdqRNSRepm0fFGseAswJx3bJSwC70/Re7c3yxq
8MU65qVAXIsUzFxdPYJStBD3OQQil66R0Pt8xI9CEyqb1/Fp73o4Z2I8gsbcY5xU
KqNMDJ5vrxU61ZwPg8J7gAMoUgOaPRfF/Vqt3mugapVFsP7dQbo91rF1OEDVl0Cp
GKiSO/113ZMrO1jJpdtdgbQy3qmPtraCS8dhG/8SiyoO8reetkFRUv8KqfOoe7Kk
4fQDDISp4hNX70vHHzU+7WztpvPV/hKfjGojgIuv+Bafwsym/xrfiA+AatHmyh0R
KhhVh9yEJA5Lg5aFu7kRHXyuLfaLbtP6smGK001Eb5KKgn/1BeY1MtqRYKJVnPwo
qyshIFNFEr/C8UgXO7RdYzYl6SjAepTaHhN590cySdpMDHfKtg5SXF6AS0Gg+SO+
PjF1DXOCaq+EOHDt5rYuwYmwRCfQo02/ziS58tZpDXZ0oD2F+qBWZURR3HAYt/iD
f+HvFk6F4RqG1pVDzhNOtP7w4PvKhHucrv8nuu9O4HwZkScBVHC0Z3Qpv3J1N79R
+lCNlV2pO6s67NQHR0EjvKr9lANETXPJevzVmJgmChue16KA3inakGhmhos0REz0
klhbBRfGePHSTZwExrVVM2KPi6YNe1/R4xRQdbnrTgo0CG+tXZ3OTMpyaQo0rIai
0ZWEx+Zk71/wQ942ABaxedQVug5d5zE8a9q9vlemsE2HJw7YY3bWaNXobbUHTMul
Y/Ym8UJftCn4JRqGXYAk4f3k4cl8dWnZb8s9ifyr1WSP9Q8u1C9BQUcKx3XMsvHg
nXQW43yObuDvLwWIrKRWgif/UH9/vQbAiIcrmGDZ1KJYocvyadL2FpbNVikWrCYZ
BTQ3hi4ZiDsP71uPDIwny6RYjzPuAZtv73wAylENrndTi+L15gQ2DUcKscO71aqk
57uV9NR222VwZsJvGdS8VjbGzEkIC/Ij4/OFz9S1196wqde4uWUGKxWLf3FErjEI
AJPw8dx2GlqXDRnUeN0QZr558hivUW+2ObVnS/2PhtucZYtqzzh8+d8sFXXg4dtu
kabXTcvCufVy6gQfl8xvw3dc18KAyfPATDOembgOK6EeNoYLzlckaxachBr6RTyU
o9fctG8cGjeIdUqFuxLDOhWiyUvjVB34btzmZdGyejkA04S4yu/i/yexKnbNBsbI
ArpslHeaGLm+IAue3XZp4vU+If7rjOI6iBT7lyn8D8Q/a/gmURSUF+Ni6iWD68Gu
fih5PTklX5tAv2txR4KWK0TXGg6aEv3nTxm7MOG1+dayNdeW+yF7C5SAs+j/EOX4
IpycKObAIL4GhGjOOk3NBsUgacO02FeGANm/F8Ideb7QVwUBk7niiQEeaoXQM3Aa
gazb74kXs7jQSx9Ijg+bUZDKqPHtbyALeCvqZ5owmYLfoF0slomjPj9uyy4TI5a5
iMZO52rRYficJd0AoJIgadlzS+bR+ywlTlO3EOzVA8T9Ra0TOC9x2jXzB8qo6Pzf
5ZzL04y51zY0CvjohiCJH5LL7ie4PKbaJJv6fICUaiP9nQ1LRKJFJl+0S5PAQ+hp
sKoZ9MhUzdYLRnzy8uFa8NCsKgOcvdD3TckUfZlzTlR7kPX7rzrTRMCpey1T1Vuv
p1FjL1e1cZgSeIxCwVqNHqtaBbKVh5fqyYXF361DEekWvFUSFN0soSqfWDxy0zvj
Zh54EusfwzV/h8KKtxI0lb3aaV09wrssBrO1YB7XZdltQyhEy6tnn5bznJ1SHK7P
s5OhkN/J1j2sDIvRsDAi0l20rirKB5PW1+zUuBL/+Hz00oHCrJqqn6ajXfYbBqZV
BfcVCUBhGzE9z/sUHySVgFq2s6DnlXx3H/3SwoTIGVekQsa5acXudJB1hHPmoleb
IK6MsJjZbXb/HnNSy6rHjSmZulv301o8NLTdnokceQwfyUyqQWFALULKhgcqVu6L
9L4YgLlKIE0RFcxpMjDq/OS3lHI+yO4UOQEYw9KtzXelC0EjAsRMb61yNBDMVRpd
O4tOxPnOOLY5E2oUL9LPb7ioc6wJYPBEECaRCKUNx/3M7NqQYTSYV2mWhGOytg0o
QpLLlHQgAeBsX0PUJP3uh3QDWH+1Esu9Wt1689TcNrpL59NQDd/8LGSSbo5Wlb8k
xi9mqpvuKxe/nGMTnjdUPOd2G640I52z+EKgGJ7bsKUGvSsF5KJ+Yvt47ibfHoYp
ob99mXcXcsfADMuujJARukQN5GUgTKvTewarGIg/gbxYC6ruvlQVAbpD+y0fNHgx
FHuvy3YfmSXShd4ZZZ1tP5Ajw9GDj2Oqh/Lx7mkweitkpjgTRbZDgVc7LtJEFm25
h4UepexPU1o19iX+khfxQd6apQIolHOt1bwFIgKwaDZflpSLrq7v0BICZA0zgaCV
YLkSjCMRdP1H7+xMtw9cE17YC/kl7wwVDZ670LRoDROTDus9Ws6bJxHgqWqxKaxG
QFLiWfNXK39YNut6EPijJmwf/RNMNscpDb48wMNPFpudvogrM0nfd/pOhMQ34wpK
nfSIiUpP5U+RYW0dKFHYhY/F/6bwifCswqmjO/5pgK/nQouq5BSuALXqqmzP2ZfN
HEYoaK0J6NtralvRWNAEe721dYFFl8wZAlGRfjnO5YHvKPPg8MM9tgNeSMVncusS
WUcQKLALa9oSIYdnI3oQJyI7tQvZw1xQjVZ5tjB22wvOyF+v2Zxg17Da4YyPk8/H
9ZOfN7HenoDw0yqzdm26xOG9Elu6p62BUy/fOivnhlEVEqL5nzq5ElpTl8SQ0mMf
wTwd2ZLLIZvyqICSGtEhnYLIybvBTE7E/DIqbveoMF2+IdeWevmGJff9B/y0ubBv
CJGHI/n5E8wMMOHMe4wos3rdDbT+XNWPx5cHreczr5YCKBUIzCVINS/GarmWnD64
h4DP9id9WjoXLFbHX7EcIyezMh/iWr1WUIxELFKZ2RnVRJBR2RVBjKrCShO/fCmE
Jdx+nZUaEHnqGxxD/La888TjjyP27g6pOGWCnni5wIPd2s15oegkxrXYiGjxpHW+
AmN2126Dr2zi2iVvaEYNGEFiTQk/s409i3HSk277fEGB1PBfTEDy0d6CIQxFAZGm
ZCQH71pUYuOfQwxgbjay+COuwsXdw0EpuxM9fhE+tXcZjJXJFRGJ4ZiIZNQpimbp
E/igb/G+6ss3oR1Xow68Rv5IA7XIKfgGpLvO37Lutid42aerN3B8iKpnAzNG/HYo
xnrQ3LV4hc2XfPofgjQt0XPpqvkpmyXGGHgFcu5jf1pf7dy/VW15NHqbPJ2wzzvH
D0oJA6s10rM5aZQBxLLG/xMF7obdF6cirb+qGgN/UOcBWFo6KE5HZknAQ85XV93u
ltrrOKKeF4IloDI1K7hVsMR9sfoMIab9X1sX0DJMR5zcp/oIvaTfRyVE/y3RrI3y
KVjghycAOo7f1JHn9qOgPQFP3tqdTqsXv5/ZLOXS1R+MGrpI2P8+I8F0S+qOWuLd
KxvifCZNXSw1A7Ge7MOUjE9BrIDNf2dqIGt2qaXgj8Dz7ZetY1z3h8LnzS4SpIl2
jtJEQM+q6Tk2tBMAkF9B7lA01BVXpdtTxdjGmIhpq2h7sHxa5qjgRvvk4MtNcRqP
dxHg/6+N72xYIoCbzyyH0et22+WB3ECpRwYcdBrWV31e0bDrBrDXgnr6KPRaHj1p
LeZfwO0MKGkfMYz2nUdPRV2Sb3Oa1b5f+xQehGouvRxag9WVhcwgQ/GQjvtsp08v
bbuRrpwyF6XwWoItyu67Fb0VSzEShuJEHPKkHBVJSimcUlJHgwCngAvPfWlu4JVA
aHT8zPIBFEgGmQlII1y2n9VhDQy7Tr9ROda3WnU6bkN/Azshl7bxT02CC/sMLvHv
gw/hGfVbTROhw+1n8qjr+m5zeIG7jLGt2T9/kh/F2KRfr08nVaHxlUQ4FqfcChJL
ay3P0I84SnU3sA1JfHqT08cvtrK47JaY1v+xvcjhzVGsl3g24xc5yBiSWdQhPtWC
pTnghNl87TwQaxjIT4KWCf+/kACLiku0Yrz8SheZ1DDk6japsmC3k23/Sl5kS8q1
hTnh7lhvOnjQeGutvT/tehTSkGO/WN+IdWpclnKj3jEAGMN2RzeMI4L8ej3mRlaP
TCCTPHYKGNVX+/gARYA2JcSiKVlgqNsx5+DVUsTU5j542vfQRYbdvPdXkkKq4+iv
eX3lLdwC+rbbsGko2q4EMRafm5SAf1U4MBBd2nL4Md+wHdPpYFLtc2r2TyZIn27Q
R9lAqauyyL4zKjOu8waH0HIrpgySoDldeDuKpnkcL1PVJSYr8mYm9sMSl68MeqNq
xeH5DAzCS/nH7gWhWdnSqaqUQTAHuO+2tA8470wLIzLk+LaMU5Psm2OlB17mkuj9
stnAfXMXT/fncnsZ6FxRjfJgw/iVWrWM0iAYQcsBjOzB+4FZEjhWCQ4RfoHmP1c7
S2q1g/EVBN8aMbFgfCjWhGGIku0UUKOvpujS01ShlDgz1qxs8Lh4jstNarrvcjv6
qPUvTcp7zWnItxATtcO6TEXpgYBz4hZCRGpcnsH/X/ws7DNBM8i3ng2rztSdgnY0
Lb4Lthy4MUHLlZyrmesXnWfFD5YdSuaQcPhIuUAsp/RpBLYOMC7+rMME8ECmcEVh
Ll227clvxBNu4KNoZ1rM/3qTNOseTOhk07dDE7gA4JOyqpNfxT2UGzyKLU2uU1ZV
7AE5EKDhBaub3SwsU0MS3c+zF1MouzEsZY30vei7SONvM1RbAViyiVwlacW8OPah
Q50Mo9VgMG3En8bR2xIm8y2manwEBfDeydu3eKn9rme7mflo+NYLYhlgEdQ/AXAn
VNr9UdyfkwTN6p9VuORLGuC9/MxJJjkWU/hUtDOzqNZtyMDjt0M+VHrTRrQUu+O3
SURgZpR8Elc/UkniFgWiiiH3uatZLnezIOqqyt2mZ67H1W9N/FGSVinWTtpFerBE
53g5ngFfXr7QETxf4zM3/Jm1LtpmpChMvDYlMTmsgOuFNUi2cDuNCoTLanHRLkGl
UVB5MUm1A0BEQ+gn25k0rFh4m71dCXvdyi9L3kUgEj4GHCKe9nWSiGsUpp30Xmdf
zr0I/51YDDq7JoWXCCEyVgapVQc5lINeCUxcPsk6vbJ9RQfsnLStAwlvtKiKlKoB
EFZFIfQHLUZoStNr6d48WNP+8Otn9UtLX/dNt33Th6hSzY48lfagX6uvCc2saapp
vv/ByZK37O36Qe+ZcsuYVH03BfpeXol0E7bSn2pv4NpUQcqHYlDr3UaAsufCRz5R
SeD+mC4qB8YQJlFM+HvtZTCf7hiKp1GNh/WM6DGJx39jYhh1QOaeVBtO0ACOWyo/
jM+V67qRb4ZVaUF27wsD+V1SJL/R0OejmEshhGErO0xMPO9RJbYAHc3ohrdtVQwx
p7dzxamyacRDc+WNVfJ6hDTl8LQRmV/jw1WK2b90Q726l21+iXbGf3uFI1ExFLZd
G/iDLOhk5BCp/cEz7hcdC3cW1jKrlRkrM1nak0DtjNpqZG1DKqQoqUdy3SZ3uqwJ
8v5lo5QthUr8n/wEn3U0yfAbK+X/a4H5MkBggcA1iPHnRpb2RryrbWsSMMvM+iUn
jL9QhFVMH5cOo7Xravk87hKqhMGibL3GVCI7ni3l9nv5NxqPY8DZTFhY0lvDOdo9
npYnx6cJSHMNJuu1KdxWLkwOOTgARvSWnggp4tNoEwxAU4ZebfnNgpvcKeeQg6bp
JheKmrBOKyLOATIVmgD6t+pYOKDt2EyHdAmKZCveY1/kqErQxR6gXU8fv53pSpet
ZEaOpfNXmEqutuAt1VGxd6HwGPBb7GIXb7maqQE7rhSlLT/Np5HjAg6UJfse+VOv
j5jTok/wyxRDwHHMFCFwPTEvH4qln8Y3czzfa4C09VLCgosgIDxz+3/KF7MSY7wd
fnYr1T7H3o0fq6E6Z9A2a88+QrzZOJmzwgfWXLpPLrvC7OaLwafk1lP7jZ17++22
lhxgua8YPmrw9j9vrxE159wfDF6k8wW4jSRcXju5iiniYOHGOQ84RRrh2LJrYNML
SZRW66kLj3/5rtIkFI/A4LPQ4VVDrqdwky+INDOVGICB/Nuy+mjoRF7mDYyE6o4d
OoxfJjRBQ9AG+WEmF93/Wy8dAV4P6AU+LhmQ6uwvdn4c7n2EVg9DN06XX2mFBX+U
ySBOUH9/t2WuMPxq2qC3DJWw7kU9Dd27MfTng5HgFxSKKnhW6vCRVnbKeQz5fVyB
tvSplO6fjocGeCjabM/Wg7M2b62UJXYuaJa/buBwFEE3eQmjQ7Nq4HOtgHOx7l/D
N8R0wkQ/YYg+meKcHkqJli0OfzpRLjcaZXc7BJwUEFW8lK1GxNIxtmIHaLjhhUrt
3DOr81xMK8+TnU9oXKXDEqsH2GyKhL2NCC4K+mDJgWVDIQNk2tnYLbYivJorvTUu
tWJzQwbj981TCBeZD+dc1tV/C1nPHhluB8DoYioZFWurDb1kDjlvjhIIO/a+Dtku
KFkXqrsYQ8hS1Nr91P9UttFLJkFQmS8yNTwqzRUgFu11yHpe2L9lejEFr/VKBfSL
18VGAvQ9z95rWeNoo2E4s3wNLQ0UhpTE1O0Flz4N048RYCdO/ucOaff7Es+gn3r0
KYSRj3URy3rSarA6KS7F8X6HW+TkEwv/ZGtaD1QFPJ//HVxv3zsKXS7Fs6f6Ht6W
8p8PLjt85xo7HhnFunJ8FqR106e9aelnbH2ZjALc5roWFmXRJmkA5hi1i1e3UOh2
cdGuW/y1azkcOHk0jTgZUk546eg01oTzG4dVrFZAWmFCOW0KiOpiQhP30eekt6Fj
7FnAOykiFog/ly4vHGffIzKr7H2+a/QYEQhkeCmj7OFLUBcFCZxYchdYvlmR97D8
ILmGePXx94TDsH82YgYxSgFke9iISq3mA4nJJtfyf4C9SX7N0e3f2HMVKx5Odn0z
9kOf0lAU4F0izLmIuyqXDGpIJyZW8Bqu+RltErwB03aHC9DPWLYQPY0qJrMMpIVF
JbAuiNc7HvcRYhmOsyfMLIJhelcHVH4rdUmP5AsdCMdroDUXND1MVk5ZKKlIVTYI
jD494u3U7dD8VfnBXH92O3tdWLq7jOdad66ZPyrG+E/3BPL6ncd35GxXd5wa6Esi
z3hw2+0+sd5ynPwse8bjRLcA5Ipl3MkmmD4TcwchGM/Cxl4WY03+kCcoIQGxUAcx
yCu5BtbzjBquLhMa5W0k2mMpYWfICUXC7IbB9hj59a2UjJUHulUBGzmHKucbYsbV
OA4LkBEloM88tXTGrI91jKjxZGKztadnbLh+k3EpaxF1MQ84plRnrC6qmjJh7qbR
qbqlVDa/geVQPY1uTLZNpSY9enFFmtimE1qji4bte5+IdNlKcOyxrhaJXONE0Nqm
WXPx9s+IpEbbz4PXCLUgiqVa6CdltzCtHYkhWFTMW5lnxsZwUEv376HEoUg9h7k/
321s88DoaynGO0wP0VI9tdfUc7FgZysFuR5dW5VVvY3PWBTZtjwnWBt/F/1JF729
LQsZlDBc/pxi3BCO9Zt4xPq7gZaliBAdfEMR18CSoNzSkZvfZ7YJUsmRTOHIvdcG
1Naocm5gfHDvemuSYe0ctY4vzyqX5ci6lV+NpVBGbYatJwH5nCczLSNeElgf6AS7
zyTUK9r8lWlXgNgUFzKFd6ovLi3+3Xqz9Cc5k/BwbF2zXYl8vCyE5UgZQTJfy0RO
GZ66mPE9ZB/4kP5rlCeAJ0zgTpL7ooPW4fy1J+lSBug3ReRT3PC4T6tkgoZUbLDL
sRKNlzMhd7lAqR+A2gNFTOPbSdHce6Lk4bcwMW5V3o9+7wJ9XNUcvxk655G6qidP
TWQC1QwrUitMPLmKj9OIkPAhqnTC7stKImt7PorGZu6ilB3ySvSCQ7ckNxQGtvOh
NwCgN6T0OszhcsApBo0368C3LX2KZF1HTRiBCcAbxfuNNNz36WCMZEt4VUnhtetw
JRuJa6yBwRwF7AaMjvt7hA9cV1l6cKSLu4Kat9skvPLqh7L2jlPUZKmA9ca7zmfT
diA7mitcsfS+yHM/Ovnu4LkmMHu67x312H9u+GFFhtKOjLDtI8o3Ni68K+ThZiIQ
Q3HcCE0LZw5f3MCj4krVWqoWq5y2vlkpYjA11AfDXzVRWbF2EempyOK5L2JBkW3l
pN/3M99ar1BPm1cKtKpPaipuoX+C0qdbrZoUwHE4io0T74+lWwKOz3As68JpYm3X
V+Oj8u3qoW5JamBG6xcNWs2MXyxHuKjj0uZwfyJ5fqx+L4co3I0jCpoMezrYC51n
LIKTXpLy5LKg83YoRkDdb+5TsIJfeup1yGNDIvsy5avCmYq/BrG++9fUGZ027br+
XaNHXOnEifjg2EbHP+/ONMiU7eM9vLBKzJCsR8l0CtOcWZzO75i3LEMqDQiNAmk2
mLBTH8xE/9An1Ss3gF4owKW2o7Jz/CqZoEJXX1f8l/tbRTXUl+GdjIbxb9vvRA8b
Ril4OL9PoOy/6sMC5wOQGLs2c7pCUl/neSoE8eCxke3uaEj7P6pk4oVZRv/nl0Xi
ZATLdXoBoMrwT69AtqKvh8TjhKWZUJufX792ExvHkE3lOBohgnSQMcOYiOAE46Fz
VnkWD7Mhe11fOPSBtTYVlgo7pa5owVUMIZ595FxekjV3ye6dfP/FK3pxL2xTZfGl
S0k+v0yoUpGJV8yNcwxUoyYA6DCOKzAKd34y45Iauo/qRX1aYrKm5QrTiYbPUcqI
IYszZmsWQmSDQD5DvLlbr+NMhp8i7vXs/NVoqhWRP81Hk1JTJ2O6qGB6UZ/1pvxS
tGNLVonJ+fakm5Vio3uOyrkH+rHGPqAMrReozO6NFWKnSTBuh6UIQSsLzI+ntc+v
mAPHhP3E4ab08+o2wQvdc/dZRqE6pGP/9GrXwXBQ1cSBhkmOpjmPSz3erUr3yibc
DYolAPgB8tjChpygieFF49yl2cPChM9B0UnEkSaWQVH42LAuzb1SiUn/iaKAogaQ
bUVlENPEPbfXI9/l3QXxJxDqAWAAIMT7gsTRBOH+4jy8CEF29S5tTc7+/8ZG+PK8
xWxMiIOeD3PUWlO6o3jjQjyhuQCRIELkZJCGyy969Is92Z+tW+2YbXBWGcjzMvRl
7CUR2emFR1Yfw50kvFbBYPiM5EprI+InphwdvmSKKt16e8w5Om4t8iKPxIV4SpEv
6kPns/ojYuzPx0POMbNal0KOV0FgvQIbPHUkza2xyaox1sm8aUTzWUyR0wxcfjIu
Ge64XO9H+eHjIVQh7DP5I86pJNpPYOzFKu3euGbZnYhZkf8MUkOm0Ot3IGGZQ+LC
yAvU+XUvbyywDGPonWeXi/0IMEZwzJyEba3Be4YIChdehmz+VMkIrtAn+aY5mt+n
AuNJ90bsVHb4GoSOF1yJ4WSoK1GHJVClp3ZDg1BmeexVhJMgJV6lEWsCQaeJTNVE
dvpaBRMkg6r6pJWXayXck1aLj5oyhHWD+xhkXy8oh6jSvnA9RduKRT2grIH5ONa1
XPCKAWI5YVeXyJhDo+2Lthv+XpoRHpANj82A/zyzN/KsLB/u3OW/TCmNPQLNJLvj
MqCWjoCxUknk8WSNJe5pXx/mduMZ70Mbe15zAkEYdFhlOYKt5aml0cHM7XZAYcf5
L0HQhQfoYCzwf1OisAYjPP9aXbvWDCP7yRLn/GYQ3birdDSL93RtOfl8QN+fTRBF
CMJ4OPFR2D7c/mUFStGmQ2sFYFzIK0xkSHSv8g9SEzL611aTC/nw0oPwRnkYhNDb
7LCI7PwZJ220mJrOUpusN7IlA9IWTo/AdrzOZS5oQ8RaSJYYHzTfp8on2gmGXq4W
IFsbE1tHnTvlNvcNDKG04O7V7pgaRSLlNBwUGrrGu9zvmmj4ujSpgMak2d0gFsBD
egbCrMM+KMbCYkYeDep29q/Ev3TeCS+E5LL9MqsbqdtxNOETIFBklUPbuYDe6nCE
KIeP8NSGF9mN+q43iIiSdcNJejGwqhOrtpONlHCtg/9uoajOrzXIhFJjDhfDh2yR
RsDsphUGMZYWD6uB9xIqsiW3EiL5uONtzdHX6m29e++otiDsf4uJJWCThyt/0s1u
DSvGt3W9ynXl01Iz1JRdx1nRSwhyFFNrUI7Zo5JMy4MJyVIBn3gtd9MNY8byGqBV
sIZBKl/GwevG78nbTiKQ2PzgOGeJkLXdXCZHZffMGrLIod4yWKtSAcN+FJnEZrC+
VaF2ylP63gjKsz1f5rz0FW8txKA8/ZY53i+tRWniYo1CPMUn00gnaN16qkm2iNNN
4w/QOJRTrLfvspQ7KGvjo9yoeLYL0c1D0LE8gq62NrYoVg1KJ2qMziOzb1TXT3n5
dHS8HXBuIBu4v7n+7fDwz4Oxp+tMjkLDHG6ZEHTQmINbOlsfds/zW2P3D55zC7J2
Z2MMCLJmWRKe4cupIQHYQ4u5K5m8p4H+lkxscVLkAaL3LAF3FxB1Zg18euh9muDz
SfXbhp4ZMaWVlwYVGH2Lf5S0y9sxCwP8JZs5r+5qYyhsu6bmv3Srea4TBipr9yYG
P7ewDEhDf596re7MmCMdFvVW7m89iibXuiIXVFaTlhGX9KQJ4RmT7ydQ9lk54hbC
YYqsKSoEB2rBPoeD/llf2gGZhYh3ikkhlcuPI8LQ+ypTXskRENt2kLi+puUEbjWi
z7C5KDQNIjnGeLPCBGw/Ekg4gP4Uq1YcUGNYLU13Vx9MdA5njaL4FIDu/MtWnRNL
ygLFZ5D5EYN5HEowCXHZuemL2CnkIqn6fUjCA16zgpSxutzWfUPUSzBezgkN5MVb
v02K+5JMu6piO3EsPVcD+cwOCRDRgD5txbtZXZeWaZ+BfbPpfEbDHgbcrudlN8ga
uuikNKy8R/B1xfu+0y6wKLYEdn+qyxNeGLdOGXISyPyeeSz9IVrSkDHdKxuVd8uc
PhyTD0yCEKsjHSuHfAhktbnp4dHK6zVaG8sNg+pisNl5NYLyk1tnHZU4SgDFd95o
iyW01gC3go8AdpukupoiENHC96FxCmHXVWYjSYZj14tmzGkBJnwDgWYLULbT4Q4x
UjuXdvx38hRF8YUcY/u9oYIEpaBSe3T+EPy03ePdLNSC+5ra+HXnJd2Bg8xUkFOo
Vr2Z2vFb3wLvsinDE5UXuVlqEHcpgrjRl4l/6jX+QyeJAZtsDXH+phd3Cw6v4ayM
BgS5VoZfjj7b1+vqcfKcpmfphxYiDZywLsSg7GiJZ4FOMUDLSOlBFFOIa6rgwRzy
cihPNIB1qB8Q1onUrv0KNBWOaeuPQD2A9l85kjUcgjK528pemitIl0ZnXtLlXcey
MI5Sptw+LmPf3VQb/53JdTc2TFuUX1vtJlLK6fa22nsSb8485GLVwyB/sO988caO
rh7zHESfj1lH3TkDfCUwmMbhZdzO171RkOMch6IvdCt8vGE3kYIabpRKU0U0EU0+
WEZtxpCv5KZ95auYKvx8N22N/HWY55sPVlkYgK+cvb2SrSjpCWwv3bsnc+1gSuUb
aDxBp0BlzKABStP82vF9kgbbH4CZ/GQ7AAkOGEf4w/El1mhqmZVbFtVvdXwtKeaJ
5kuk+8w7Baf9bLHnJlCcY6kzpFVB0vMYsWWy+OqOgjN69Bt8etgKL8DBOXc6Two/
CwFvRHd7ZuY2mQpDhTCvUiR1u7fYmB631PRGjJJjHpNNGaTq9PsK0C1mbExWum1y
kx+STj0esDyKnCiV83wJxCXEOnytc3+CILFI+03B1tcSMjanqG1Ep+ZQHqBmn8mF
TRzb27UghQIUjc5h1UW4a0wpsa7UYsIV/y0Ogf7p+TMhfPR0baLUUWLYOgKpNGtG
zZbqQpvb7uaeReDfinrQX7uspnVxGg1yWs1K4b1VUqI1C+gOqc/iO4gFXK4AlH0H
P+9oj3xHt7caDVCerPY7dQxg9MKZT6YmtsvqL6yYXTS9wN27ccn4ayJpRf4IfWup
4ZR8D/Pg5rvRq5JLyV5lkZAmbn2IhhqiTSoFON3sjgd0dfkv7rT9DbwqBED55hAL
50uiNfdsrwkeJO0YDqIAL0HWdvLNb15tNXqSLs5+aERoFWIgDJ4Yr2oluzMnpJE9
0mxdS3cfuML1O2AilXGtPOQVN5ZfFUgl/3yi/g8AXhpHBYH6Hc5kKkmSauE0bdJ2
84G9GVX5u8a1/HsVQKgDlIJtNojdKoEaoXVUKAjLIGvD4mrqhXuwFsVL09kEde3H
dHTkwhpnq0Kk3DzSQhOq3MYk059oCD/rTgI2RbsQRGP9C/VJPfQTk9iyeSJ4MHJ0
Z8IvdYBVoqtamhNETC9LGhWwvCibuEJBJMxkyU5NEWRYIwoh+N0NlZuSIbPv4tfF
lzq+ZQYr569c30eGOgWMJb9cDVVfPIZpD1hvi8M3n+U8/qMIBU0+eih4VejTHMzS
nhLlLfVWTdGBpQmlEsd9HtFnm9o3Yken0CVmXSLQMhHfeVpa78PyE8FWHs/+7MEq
WSi6Gi26yb++zR3qQ5HrxXiPvH03mHj34WVb5DSiWZ3zaHD8kvKbwhiOTwiD0Q77
zZO7qDt7yW4erc42BGnrBLch82iRzAdek1+G+tlWgZHUfK9mQmhKVAjbdHlCnLBB
KagU1d/gHVvQ9Z+KdSsGBMPNnighck5qPtiG3cGrBw5QY4Xek54WMBXwIBeXrHw+
cb7ncIBqU4ANad3pIEiFSdo9tuUDelpybuWRdeO42K+Wsy3q65qJJOYK76OE5ULV
0anzVD1gKqOe2B/l91phhLTIus8R8PZDZPMUUlsGhS9Us3lkclAsbKX+MTrtLPaF
bxZnfVH8NIS0pVKi8NCsYX8ZxOClyhZXv5MG8Rt73I46++m+K1TkBVOvWaj7/aOP
9aKZPLQwBcty9qzjJZHnG1Pf1QhoiIngnK5ceBXgogF3zGV56q45jZ+appapT+cb
OnJLvYj4TVCbNvJJEIxNmE4iiEr1DrgrwevRpUGdRobdQUoSU6q6AYzwUn5Pv4X4
9/kWLn8vxzEwYzeOXGNO+HIhR7nE81a4bXtyHQWbUmFanLOsxzHpeUIEZA+OmOyw
3XXtbfRg9ErUJDMcmFTApZ42O6lD1zR5HyjTfMYarWYAEFN1ae3VCxcuA6JXJCsK
aZptmL0aP2QnvIAGMwyJZmxOt1XygDTmiqOSq9Llwbj5Cpf6gsVCIklU0DYwzOqg
JvOjvz49z89tpEywkNDrORH70ddQhhQ3kW7BV4W3YySMyXNUuf7Mr5FFAPuNv4Oj
yTcyb49geemb/6xpzu4La83ybfKTwNHpcE8ErURNrC/orVKyPo7grRyZh+sFyp/E
J9NQ4/aHiO6q2B5X/1or9fe/yYq7btlLdT2OPZAmop5MfVFPXdqRcD55Ki9uGC5q
veshrubcGtXe1iqsvTinv9StkGiA0TuN8ZzfykMlUwZNiM8kk6RxOWdP2GLsVTaI
SLHQxpDWwrAN+smAjgI+bQ3fvMN6djtMj+S0IRuDYH25D0jQSFvFPS2rL4Ifo9sy
gzr7xFjvrB/qsLAx/zvs+4ybXmnXJ8T4lzCvyv5A2EuNcljkLU9S+DvRJKLZCM6A
B++odgGK3UwrTZ+ez5MlcXSi9+tJMlfAAFvPNXYz3g8MzmK0dbmeISZM00lhKS/e
ySOpL5nvlOxQJElORB6Pvm7ZRWiBmeBw1+6SZQWYV9LG6HljqHKACAF4x4x4Pfp/
+GX5q9ljMU2FS1Oq4T5JJ6qUlrgVOREsjH+ZrfrkK7cV17VcY9OuzoFRIIOXZ7t+
0O/l6TkUCcEIuYEX2djWi41PBy2mDy6Q+OdHUJZGkNflsnf8kv3gwUuz3/a6W/zb
Cm3b6jupDGP0EeJv5OMndwQY4jLTAFiiaUUbuxQFuNwZFPjHOlHJyE8sU7dDuZi8
2aYgMHxe1FEgJLNgXKgZAIuLjfd8gcGl2sA3Z8VQmcikZf53s76Hx4m30Ttjlk3D
KwPFJD3Z6ZlAjv1bLNc0JJHKL+IWCOfuFBdo8kPwWeglt2wV5vg8xdFsfPxLvBGt
1Z+/FTP6kRvErytWTjDfBK9DmluJRoc0St0h7HpEsY+7SH+w+rarKzthYvVQpFM7
6mYPETLsfuIDC/xjvtYMqBASJiP8jlhKgZN13VU5H5VO/HEu7WBgpCpkL+YiseDo
e6KUVdpDV8l0JEu7U68EWay5FP5sP1HkOd3K+EA+z7tZJT8MHk+G8RRs9zmzKfek
faMJzsXl/K1DGPXF9TFTS8DUVTgmNb91TXP24ElUzmmT8YVaZdMGtXRtLdNLm+o6
M0iJyOqeXj0R56hl+LfRDrGprzoiZYxJ4IrtYSAnwvm4uTdMe7QELsMdnbTqnnpm
Y785kVwx2TwBJGXcmjXaa81GHORn3YNY5U/lkZMEGdRKd5Ex7L14wlj+y3QWA8R2
06tf4Y1m+M1GVysUrJlQeGHCdw/bc4ds2QxJgYshHeNRabOFo/At/DfEDFNMBpSO
cIVq7Fm/MIG8VLprCSa8KIOaWU7ozbpCIpNfpfU7YAe8566mVI92qex7lCRZtaNs
RjYGUJiNmR1NbrHHQ2pJh7duZi1psXsb7K8ZnRthUqq/EBS0owA60LxnCsGaouel
nqmLU4Jynd74tIU03kr+Yzox8dfhjURBQex0NuGdc/eVWir9CEu1V5nHOHTqSiBy
4j8GffeKiIroz5Iv7rSGZacOSr2sLRLIlIXnE/NlptUyH86l9uMo4cTVvUJFwOTH
ccmnec+3ftsdhODPrrJOwAzOrU8lkbzH312D77+Oymi0lZ8WaBios7jmT6N1zc9S
UMO5RRtBG2ZEYiC0A1f0gMhNu2NIsI/qO3qm5B8j9yrwU7MkeRaoNOYlLFrX7Qmt
Bsxdx5mdRknwGysoLNkEHThx3knlwylYyWm4kDBkzr53SCS4QD4+rb7bhUrSlycF
AWBEg+n5TkGSsUbAaPL55O71clg2ioVepFcZcS7R2uV2yNgWDoDCsdiypaPwHCRq
bWqBBtP34s1DYSwWeG+bkJEkqmwbFZtfoSikYXB9+HXyQSw3eUgPsUo9001gb1jZ
9PG7TaW86oVTAFs6mUwDLm7IgiW3EC8Hg6HiiKFi6N1gDR3DddJ1IoQkBB2UTtNa
+0uABL1f/IWRUEnGSl9YLHslH5sy0vLuSWaG3RywKGWXXq7w9EvhEOgZUAwcqazk
w2s/MxV96blkPh8guTDvtlP+hLz2JdKJ8g/PVme+RrC4UB5nGqxdQPPI8VZt9YII
TFa2tz1EtY63Zxj+3YbbGWyV9iQ476DZtZAbArsJqfqfE8dhyw797YYesxPvTsGn
QlgwArX0ACTOlTu5xxGWqrGuEg71JGd1PiTk6y9fabJfNQko1NF802X7DhEk86kv
ZZXn5bdjdBh6djCa7l+rFn0FaOMhfhW4ZOtD8m5J5UVRlNAe2EpM4CS4IlEmBMdB
56/aDMirDncvFWbG3FVFgz4mlb2Dv0ReHTwQ/69caIQAM0HR2CHUNJJ6jbtqZxBw
EVKj8aNQQoxyXOhVr32VYubik+Z6/Vxr4y5rVZqESz2k3FkZvWfA/u3+QcpVAO0v
b7nm1spQRoBTvpfmQFNMOt5mhnLKynxeCPGPdSm6XUfMW9+hI8TAcelHUALIPV2j
JgEOnnpVsphIyQo29UqVGW7klGa3VOeVfBbQ3IjhrTdHT4qiKLbjWYRcKbO49Lll
7evUuYoRECImAzxIOldbIaJgkTbbRQdWNuZhIQ7xHnpIA4MArPfPT4YaAVGZnzBb
7AFtDQsNQL3GRoIfgbA+faomoaJIRlu0UUz6BqEyr9VRvvgIwIeM/eMLHhcuxoSR
ORStUkRzrvH2Vzwnp1JCdVNDSPJWbuOJXe/jkS0s7XLxotYrFsJKC4YaZriE8ajp
O7QbPwvYk3yq8GtOSc93M06ATNFDfv/JaYaWvvk4vH0wan/fmFnAoG0ONb7VJjYl
S7kB4GZXruMo3Z8zAk6NF0LfjHYfm2Dv2QNhQeyEuNlIItm9gu2ciRFnYONlDc1M
2caG45luI5NL5uyUHa+BXgw1FtcpGdqg5Aoe0SEub91a1EpNXKOMTNtZVnzPxOfP
Y07P7E5A9TOU2VpDDIMSLkLWaApCLX4RR7qWDhNUUhIn8g9EShiPpQ1iEzPPxTT8
cQkMzOVQlFBZdVsFL/xvNNsL6zVccbF68AUY67DcLyH7BCFXN+x44/lXsMgEYl84
MYOPt7S7Tr+pQ7ZME3PC6M/8u9q+XO4vRUB7wUJTBHRce5wekXSvGhgzfIA/UTtx
Q5fRV/uDcntUaxPicnpHcRl+YqqxmoS1KnGHZVfS3Zw2OiM7UHz0N9LwLch1g+qA
wwpO9ni1lS3gXYWgKBrhCthOfUE991enBSjWPpZlFSGN2kOFiRvdNlKA5O4wcvmM
BvKXHi/yXVlCRMTW2WuGQSa5tM7oqj0M4vmpxQvP7ZYEpRJE/Cz6+CQtaq0NOHo9
9TMH6DUQvtpAuOkqmIdOId+p03wnzRX8mdTMvji0K+/PjwZFo9X5R4g0jg8AL/Iy
NDg5+ETUFAqqg6oXb1Yh8ZowJIAGDewAIsH6GMVCGnoZ0f/NafFoZmApI41n/afg
eU58rbVW6sqw6HqpBiOG9RrQKvPH7LQ8TqgEBxifaFIMhIluJpNJBS55RXnKlVDb
tNsBYNzxff6FrI8XoaFguYvOfOVQy3Byb2k69gRaXNVELnzh+b/gvQfeS6g3jI7K
OmZjo1L5ARwiw+c/KfQmQqbwPnGWsnpvsPgLvCTEXy4iLdOrhjSGclbmvpq0CIlg
AsbGbjdG0+U5s5OM5JnvtpgBoSLdIPwhB90RbUHiZN+TqFDt62vkOdq4eGlYfgwH
J6V4kTPecaU1pQ9i5c7YizP+Azh7r9aQeaPr17trqzEuneOPktigNV0H+5sqJ2jK
nGbEbg3hOd7fbjpwAKt/FKErxPVgDtnaq4NExglgoyBSx+QoUIBrxBsrDq8rquLy
rZOA1YWUb90C2NLLoT+5esfeSffRmNhJTsZHdocTAeXrnkFHzXVTp3JhZzd4lPtR
QgFf582jL5k+DdtQDqp2tG5EDIqd/fCkow/9WfdGUnVBMIF0Ol2vV0Qbm+/7puOX
n4WME8REf49h4S1cphxJ3t4/jFglwXms3B0fYrsroty3+lRtW8G9SP51+kGWdGJl
hQIDkkWg+sShwKJwBUDsAeD+8ygYOg0hud7SKFXT+ZMrCOenIU1pMwZuQ3ks5Sj/
WK+rl3/9z0x8hEPmU+BbO93f/UYbpdOImVPr+I3axuiGkShab3CXicTI5IywMHOn
IgP10PwCTYo7g3orddT7Z88QbbgidtprrLEhqZzc7I7DXpHxlMl3w9VlILWOALt+
j46iSYKDTDbwFjyVm8G2YQ6OmFx6vWN36jmqkq5Zi2LGJr49hYEbKcnPxnFD+e+o
nqEGU9M1PCgNBKtrWI6Krbac4sXazBzyes56s5x9xio0KCFpSsPACKIsgFGVcN8p
ypJQDCbqQbCcMrEAiWwkRAZqdfcAIxhW3l9AT550pYkJjckj2u/yhFU33gE53gYb
0sUUtBEwobkRoQ4VQaqmsljCsD1twOnEZoCTcKE+7zerYIHSSH1JgU/zU/z4zNKj
A2U+yAo9y2ryH7NzT4kWEvyV8vck9J1Jeo6tNYjIvkguotCMWOVlLsP+cFhWh0xg
ZrObANQ0mKvkWQY+JC71THW6tFKk9woGeYBrqXzm4xW3B1OLLOfZUCD9nNscX2s2
Ig3fkCQm9JmEmuybAOOBujvarVZ63JXpv8IU5BG+qZndeqh7MWbtLoMyAJNYmXkd
asoFhlmqx2S1qfHBUpFGUbe51S+w27iNx6j4gqMp1tJnjfOTbVV388HJax+W7s7S
TIseUaNEXO18JjH+64UIc00h/31ynux/XXRuv7l9LToTBQDmxm2saQVr7O2AyKe6
nH1r9p53q0k2pPY8mzfOuXAs0mthmVCClQlIeSBPahiyOjsuW353tgTAaX/Ty0+d
00BiJn63KTpx6G7PJ0fWMZXGM4xP+kthtazri7/fvcEQR7fxofebZ1q0JHedVbYG
Y4FRVTGPL6OTTNxGS3Zs6lZejOGWrmjVXzEyTK8c7D1ygwqmxXvdGRSj/6CAEE26
AjmD6v7MetgAK7v+fuT6FuzDNpobolsr1SRROyXe2m+0LHDh9zRJexMnSJ+NcYPd
ZRGGsuHXYBG4+LYJGVrDGyS3eoHA5LZlxdoaeerVoMvTBpX0cuhSsBFH/u8dpGbX
6J7Q0RlJRLTRmKjJ6uRWp6zl/3hSjOpNtb69BvdpiXLLTwxh2uz4mZk7Gdl089lT
XFjHeRX3YNnJQAMN0NhUJnF+Ky3yi5zdKlTnxhM/RGJkkf3VOZLGnBNWjHjx91tv
uGB8oeXifdkQhfslAHHgp5SFxV/knkwezZMKY7KkeXUQMgkSnIGlR0+hBjwSdXPZ
Cf/8S/jDRp5+z38G6QyDtRXtIpNpcvd8IQrxxlFc2LPhk/1nGZKdzpET/sO2Le2t
6RXY07l/qNr0ISwxNzn5gVKGA7BPDM54Wguoz64xq8WllHi89CVN6ir3n/7D5sIo
BpP/CZwqP9Hq7Uf9qFJeAIRBtM1hMUq0Gi8lDSQnp7gdVAoAwosLp/uZ3tbTrl82
t4XBV3ZzLKpE9yVGpbKRdFKCGzqCIZt6T6T1T7URIJI/baxe709vTTm14hdUuOWS
eljcx/Sh1QVZdiIFGSZ+1vjfpv9ERce95/uhruUPloDP9viL95dbtx6/116wDtEE
uVIrwzcNHqK38OxdcI6OqVPQV9tVgSxGj8quFjfTgGS33uqiOlMWnLQv4g4iOyZY
+H0jRG2LHJkpn3U5kSPAboD1LUH4lr81IgKJjDKqv068P6FNvD8KmOxUUcjPtKhW
8kBzoaoJg6/a0kJS9OEBHunVkS8Cr/zcSPZV3dBCQfTjUChpBbV2vQY9KF/ppZUA
WjHJxQbEz+NwheQGDtEFfkS+5/EpUlYYb59HJp4ceFHcgzenNAkmwX1nCVd6B7GL
CQEf05SJr/Ek7ScBpZ86OnVkmC0eAL9/tsn23UqMUyG1FTsW3L3519AYQ5oGF24O
cBSUVq1IEU4SW/Oj+FjieF1w52vD5YjxfAL9JPR4gsauausAyX7vHeyotyzwYzr4
qPfhreBbrVH6B/C3iOW9Xi44UWZx+m36Si3eZw5icVPbGVy8SmXyqdS6/ZOGXbXz
0EaCFR+A6c3A9fOAn6YEZT4ija6Y5DYdrNahe+vy6853lMYBBeqEn0agMuTB4yw+
IjyrF/cnxel8hoQhGGybZZvHYeIgnFfFsRp+oqAw712gw18yVVXeNQX1Ucr31IQM
yKBg6hfV+Oewo3iHsgwAlinxpOmixrdwUhzSBgyHVEdBAUu9NcAN01tGW2C11aSY
G1Q1MnXLMJDnlMzV+x8WyCLOFtE6WTI3EQPugM5/Mh1qCtf1fpknE40oH671g5bR
qBLsBmchFu6nHKLmQX/FtJieF3YOLPE4DkLVSbJoqLhyqGPmN+UVTc5+CCoDSGYy
EpAECYFuroH7rgIi0N4AkVPHpkGdmt2TNK45GDnXj28SRizxmElyXHHvMC75Whog
+VC8xs6AbEb7fyHBZ5SPjkJINczJ2bk80iYQyJfgtHnIy+wIMMdlyuJUueMD6tO6
WTTcUgWDIWIkquS6Xe0cVpRErz6jGP+A7PA8YNEkFL72XfL7i5E8C2iNBz6ksDFd
c3n85ka8EYq6pw2izchclvwvywWJBOiE2lTLawT190DanrphPN8++TbPMD3kB+S9
upUb9rXIJTo6fsQPJzwUPy+aQIJpqpwKEbIy78eNeEj19uolAqEX1WjB7TPHixt7
//gDHeJDTL1ZszrPkX1Wi/VyRwpGpxmOdRVZwItLrZTjzrU4wHgoZ/MB03Xkwo4l
mLx0NQAt+MkOzkBBaEITrybYFY0vx1emHBhJFZUTxBapyZecU7g/Tn08FHY8HXYk
+s4c6KwPgA7wFRi4v6sIuUzjexDDWo38QCFK7GZRDk6rs/4lllbLvUtJfYF9ay9k
Tw7s0retcBI/b/7BvNzhM1kjewLiclccFSrtrRw3LnJDW2pIgr5lswu9ZlggPAkx
tcGO/qLH8IOj+QyB4hC9oNsTVCb6gMl2BqyMNz92+fG3nSTdp6J9Fg4AkJ61Mwf/
YiNbW8pkpOwvDGsRT3FotxGUjLIT6e7sttJGXxoLqqgueJy4I/UKvj5tqS7mQaRN
GP1pTk5wG/NCPFDHmm4uIGQQUTJQhDaj4mN7wlayTw0KFAIKjzN51DrUzN/DQJpo
KX68k6DHXH0JppUvtNiDgKVdQCDIOaeHCvd8EUknnCQUCDyWo9ehT96DjPKoEit6
vlsOcGx5Bxr5aTIfDKWmc68oqEYNn9clY04yRQF9oKGnqbNUa1Tep8ymwjhS6B9z
qX+PS5nbY8V+7xeh29Fdb2iKX0KqxQpEgM0o2khsTIxqMhZ6LKOLg1R2ND3VoizJ
0pzOGvZMLOI8hudNiMheAu6s58aZL1KrjhlT8v120Z9P2SicMTE62DswDTlBSZhr
Zws9yaa2RkuE3Tnx9q3dOiWLf+UNPxqFmqkjvwYxmsgCCPO+Szz7B0VxmXFo4ZDh
o5Llr89wXea6h/lKqiUxGY01VSkjbEDnNO+mXpw3b5E4WAe2AnUc/v6oEJPUGMJZ
J38a/y5pfayYlM7xgqBcHFg/XEhB3ts07s8421Ed9xe7i1DsQPHF8mkFwDDTl7Cv
q396ka9YjM8JrtVAd8fYu6932cisnnT/ltFim2XtLkZRcd7hD7c5jKd2dIceqBCu
NqgvuT0Gcly1HUMbB1OPuEUDGUVVxKoCMxRDGxLTz/FZgJlbsRE7ZtRB74m7Ldjr
4xUGbmY16OM5H6x+10sx/cP2DAyw5QyDccPRTyoG6QtCBst9FgBc7Zo4bSlRrd3g
tSE05SC29VDD6cLEj6nimrglYhl0CNR8XivbfPsV5xBj3NYS5F3gBUDwipms9SS2
aj5kcQFW2kyEZmS/5zWLhTEsFVKLnw/lWqZ6ao+laA5O45VKbCL0MoMvsif47rc8
4Fsvf32CyHQRG6t3awXadiw1qVwgtM9WL24+8LZ/vFWffnBrbnCWassSJPmmQK5H
9KhZCzTTzdV51QG7cyINafi9fmaRf9ZXXjnQl9pDO8vRVWlW7YwLeiV8nKq8DruA
qatqF00aY/O1csnHYoL1R4Bxe+wdrktQ4WjZ8OdTn3yZbEZabZTt74aKXC6k+MkU
/mlaLhBU82H/fMXZdPoxQyx7vG+M1tcxnwS6bsw6VML9ULc1K7ctzJHD+qaWXqGj
4ZTpSXjdXtAhdyjeH8issFhF60SmC8DIpHDSwg69klPOBghXuZoPNdSyXTkdhPgx
m8oFGaqiY1t8cML28nSfoQ9PM2R4uWJgxjTZsUH7/6SZkCB6t9zjmt1t9Vj+Fw0x
dYeFxtBLc69AgHnuHt/yLJpp0IyVmHPXJXn+0qEQxHlKAPRJjZM/MGD86zLVhqn3
X7fEWEVWJVCby2AMy4msbAep+A6Np1/N2JO9TdtPTV2wAFnV32CR6y35PthWbCBY
FnvrvrwNZjXCFNPGTQrwtT6mmeaYS7HL/QvBn6hBpg6N0Fv46TFvYiIdlbQgXz9H
pFAkRc0OKMjC7imNiVs9MDgXS5ntEP7AgQPKEk8XaUiStJiN5M1CMwuxK3cDUff2
3+f9kXS3OfxrlK7E6B1ad7SjZYax4EZBDbXWvuTuskLsiu4Wy86LjNj+Oa2DGezP
LdP+BbC1KJqmlWT00ATv2/ua0LcuKaNPMNAgiTcszEEBq4FHf46bVfbw0jIgOVGc
zuruuZXvTlvzb1c37ebgm9N9LSwJcCyowED21IfHJehMsoqco/X/fTKyHlzhDp2L
4nIqaQLeopVYaemjjEbxnqZCRrkv4fOp11vNBQwiUXvEkf8uX0ICLGXenGy7kdpB
/QHO/xi/6DpIbzGENE4sNgL1RebyToysCY/a4ZrDUvLFcpDPGsS3KX5DBgbcRt+F
wwB4hRuvmV4lKxrEUp1w6JUHFZv+02oH681ZtAYbzDiE6eqDuYLfAsp1TBF0ekHn
JH36axOQV6Uqr+WFq0apWpz4bJMYhLPmtxhDW9FOw0nI5yYjQhfeQr8aGbHGScJt
rXB6jghqrolh3JRUBRGOYKIFX1FRN9mxxA38zaBc2AVJ7f7UPkoT9HM6GIsD/uRg
uzrV8ifZe+w7G2boXpcD/J6Ee1wzNTomz2v1yRhFiviUuK/Vwy7BFDzSs/iiYC45
AUKCHYFVzotmOS9pHIsmhq1RkXEj+bE/FqpwC8YMABGEUdonstErM8REyk/5TtD2
bEQ34fdZIGWC3WQauPEU/9g1rPBsvnITSsT5nMHccfVCNlRGwh8viqalsHn+Ea27
XWkNbr1YMJCx06nY5TWGJaGD9hZsIQEaOQnksYVnWFP0yrRNwrnEMJbOBnpQV3dt
GP3uZzj9rfvgNE/cwGdbKeMaqG0l3msHI3n7UvFTvW/Pq1b4h5GFnr5yR7XzxpJh
4vzKxXMl7tIBACDNnbhvXNx/hikw48ZZOsQq8ZvgtpaZIQVBbHYpFTebxS1fa9kp
+LlFRE/6ZK85F9FLySwH32jP3W3lsKaXqW8f+MFbfLxif1kdzQ8afPiVOEmh0qe0
Z0fm/0tDYYcx6D2cxqGaWBSSMKLvRHu/0Q/5+FtZOyf47stT/wca47aR+S4EA7fZ
CwdVtrZoxPLUYkkZfvXn7N9PN7lu1lG2bzkQBahRIk4yUwAVclJMtJLD7kYVTrm5
HZSXt3ofQaOTABADtIhqLCx2J65Gs7i2YL0fgIyW185ibBBuct6spLm1Sypy7qEq
GVlm16IwVC7a0DY0oqRCvKlMiL8QTHz64oQ/F7m9Q23DAJcEExp1X0aKdf6jVF3q
ENKing3nErrTB59weHxR4lQ4M64WNfPgnZICUYYMhNt+MMeqIlo4D28wjJWCh6Bf
98Euy4GkOCbp6NKBSo02A0dBoYWMpi6NVk+C934oMFolmrpbvNleEIUsz6bk19gt
gVNWfbf0b7YIdV+19xv1NvT/FFf7E4tCOkwGGCOBv3aBRv6mOnnCL8kyRYrGPWtT
juMjGAaHrFeuJjzrmGXZDAsjUatXKbXyRuhyTta/FqpaxLXOpDgGkxZvhAXly5b6
xqwLdaKINZNp0RvIgYUM2zJHbnO1OqCRUirxKtmLrLNEHuuqHK590fMp3u7D2mxe
+7gq7WRUO0/RKLs1GhVxnBm4X0gdrMQmOT09UAs9aSv+aKu9PyzRyYB5180evjDs
4Yq8eWjktT1gWPnXkNriukIVbEGJx/8Tzy6lQsgym5brcwp5k9WSSOckDkjZtNqg
MuYFTQ4/QqSb/HJcDzQjgTKSEYVa6KsYqsU9ql4WJ61Psi4KdkktRhviJoAQOqji
RzDwfq1mgnnQi6y1cmMG1YGLMjb9AqQ2XKXhwxpVsPOg/CFa0zJT35n+GF4w3kdH
7XWjPVq1ni9nNJQyxBKkPylDCCz3JTfyg8i+04Xkx7Mo3DnfBu3GgCq0Li5bTyeQ
zw+NshW7Qj6iTwF3TgcHNFBLXfqlJjiSKdlZZs6BXh4U6NiUxbP9wXft3xFA5avl
3wx5uxXU5R2UzcaLeYeD/FT/fWmer8q6dG0VD+HAPLoxjrKTt23LBKBmI644bcnK
tO2JeFN4G4OZWqBvppP4WyLv2uZTmcMTDVBYWtAIHOVV15JdExcUbLdLtl/DIZgW
csUoL12+RX1lLZGD+Kj8tn1XyNma37AdadiLQ1qCwstiEOZ7GaNmzE/PRkw811GI
5oTu9l2U5S2zcVb+Y3Ep38gYAVSfsBGTmN2XVj9+1mA4tf0dc/QmcqIYwXKflCoG
GFK1x1VwuFb0FJtBRyHe+ar6xGp41Hy3GzNIwmZRI58q/MMSUc6ZgEDdpg4Gss3/
a3QxkaJe1hxe7n5ndLiPR9bhLgSLrLpzle4zilTVpavI7O8+QQx4kV9EM3gQ7nWo
gV54lfRIFuK86xLwTOqUTnU/EVD3IfTMkEJ7EHDoPAoNf7WMsm0BWwd+Y5dYWlN4
NVsFUh0shMocIu4O2/KwLBLoRptjTcF6PAL18UbgT0kjLn13QWL6We7/zpLSMVhu
OGtstukj/IIGU1bgMeBCL+4aN09bX/aSJaZjpTPYdV7d6wIJ4UXY2uRhIzD1wrod
KhLtItpe6Mg5+03lHMJNlKmiZaoQgNe30tBbVlAKDfqr+jOrWQzqF8wYa+GeeVz6
/RMtu5iIXSxxyRHNV1aejEdalStxa6SbxZoFC0ts+C4cojbJxrjHjCu2NV8Sa7Jy
Bi2ejRMAA1VQGOPclSBw6A+XocCh6thMi5DD1UtxvyH096jiHvO6pTmrx4rCdzVJ
/ua3Yz87Xxr8U7faROVxKlgTq8koCxknSAoKPdzcZHUzt/q7m3U6zraQB1htttkQ
fAPmxfoCDdQIaE0dRUzMdZI6dKf09ojq4HYA/UNso9A0ILEqJc3X0y1XSyCMYsmD
Q3SuohTddE+v0BDMxlie7LefJnsWoGq6mPI5RSnu/6Ef87XjvDVeBcDsoQuUXvsT
jFq1sW4XdW9BSKd6eGPoZC5tXp/ibbGHjuaHOWcy7cabJuiWHCYM05aXlSqs8B6P
uP61myZ+sBvF7nqr6wxL4ejscJbBDzYCVfSl324jB7XuSQvuRmQnStPGxdFJsIXH
3uSwqDprjtb9eqyb8loWcsqvpzfHdmcXedbPS4k5Cgpn/t1m2bCIvKCTGRJKkZ45
ReX8d3oAtEUUQlRbcoKnLx4h5H4W/UiRQ3AKF2d8vV/0VkATtnlnbFWIQ0yCTBxr
0Sh5b//gF8EFrWI2kFlaTdO8UlJCiJZuoWD00/lQaxge+UAdBYKwSGOT33EdsyWs
QjJApIstShLe7fjE9h6joGNkTAMMF24NRMiyW/RpqT91/NVy0qnIgoML1+aEp3bv
/R05O74toV2UJnkkHZPwj3OU4rYLFp2HvrGi8c04OwyiqiMZ4/a3yBv4JAyeMKTC
oXWrsnP2zK2s/S8X81qn5k9fyxBfR1K/MVZ3pCDlJM5r0jpwTOoxKtEwi1riwdvc
P8DguoUOKtjHKkBw8UQdpf+We7KbDh7OvHRBlDv6xhKZPJRIwPh5kZxov+n4Eygh
oJZfJO1awPX1RzUqOIScapBaVI8EkWPS/UGi4cZFDycTZ5sVCspcBRqsJz0Wznee
l7EhOkLXsqYsEk6HCOx9++jHwZN8QvqtRaz/U3OTkJuUGdtbxcFkzyx5IEQxiBER
yXwWTJNzRLHXiY7sUbL/C2kkP1QNW/d5/ip97UJ8AMn6bSM5yWxxF5pr8dUZBaSg
BiaD2V0CrMMgmdK4rOtY4HZ4svJXOBa/bti47xhuvEfZNUbU3nMogQBJMb0cwCtP
Cu8Uqi4P7KcgIwkdGqDTIJfmivJ9pP6OHlAu6HoQBv7dB1hpFIkf39QioMA44V7a
UCsxV+bj/1eYe0PH6dIW+wiNFhGrZkjUmsLuBywqJhpEXDEmva5foXNenxsPM9JD
TuZlMXRg1YcdRcxCfsJgiE2rka3TdiI+3YTODLjPzF8Yz20vsNr7z7QukZBqQu3V
FS6LavfpGwFQQJkY0tymzy3H4/IVkJyFapXccsmeIuXiHvfcoCQRaOVkFzDy5hKq
zYWiLrdZAXXfogI/3dBybe9fUIRcU2BbRi0kwhuo6pn+eQZsTxhiMsf7eN6ctmCX
nFXD8UzuZBI3bPkFgjkayUctW0iMQgYObuHUe8Zg6KiKKsBcQRmiiFqEKlj1UDIP
Lf8gjWYQfGeeL1Z3tAsL3qFDYCzwGQn83c02YhMYHp1sYUsF/q+YozYzo9NN9oOV
E2FyLe9z9ybeqLqffTyWYLIBlJ3ERaTQw35S5nTEKghzPWDXdKZ0Eb9xXeHc4ieN
kzKxPXMcPu/AWIq3qvCcncj1rjPUSFU1kMdxp6gw5lfQTg49i2PrCaS6uAWkoPE1
R1Ccolm4jyPWkGhMPkRfwMmjGuQT+Fyo8VJ7wrK+e/+3PdluIx62hENx6GmM9Z6a
AbB504eYjlObWZItR+xvK+eVm1rYUv+/GDRurfymtOJ79o3Z8KegIbgrY24EoFYi
HqHc6RYaqOUlonQ5pcm/QrQmVUbQH12XBqvr0gO0XgAowW6ss2r7Y7RVWqI/QDOC
2GY8Els6D8aP6dQmCsojbZEiN3+FhlqEpzJS7bq1E6nmF4yRoVaiB2f4iuEgZF7w
X1YqH926lvItXpoKHcGI9WM7MiXSAH9c0H2inzEmkbv2yz2BxrLeZjoWzvdGJ/Bb
sZmD+oLTchO9HLbeV4yW0Jl7/9YqAbetJwwMNyC0psTGUsh7gbdcz1bzLe/HWgSN
mQgGswVHILUHCKTtNOxb2gJBWrR2rcJPUb1CHL4J3+2uMcxeGAEodnamWt+08kU1
E62xdKkLbs1Agr2LkWhG9nfukR/3hhr0tqlE49UPC+Pxs380fMikfkbCyDkM2kid
WIJzkMShkLFXqgPNftuoF9vVR9mBJen9YcBRpL5dJsF7F/0Ek7RmztG6EUzttDR0
jYLbU8Zb1tHpQOvjZKzN7vdi5J4/Y7tuptqVoXTdU9keblRgMc4aMvDeDE36BD2y
q6NIw3ylvQM0vooNCoq5vfVJfzJQ9Kj7lhBvWkHkFbegVd8o4OjilFVje+BOWIj3
BWjzI1u6Cn0tAGZVH3W2nF2djWvL7SJU2qOkR7rW5KQukbqSQVJoOkCEOTH+yf96
9B4CKPyoD0XHOjdp1c1GompYL+yN//ujZhD71ke9U8fdzwyw3F40M6XCIIJCP0PO
11Rm0FV8qtQ+XkojxGg8ls8eR75Vy4kqYCGxZwiJ3JqSnrdiLfjf/XV0tpwh9rVI
RR4VJpgvXEzIV3+UCvbcuciyp/pXURa7Hoti2s5+V/ewLmzNofU/OLKy/Wvb511m
uthQFTcu8Yzd4PGuam/UaYCBnEnGd9QhjHNNprGo4V39ZUsw1sfIbGeSfeKEe7gf
dhBCx5KseNKcHHaGC4MwPZIbF5PFM4JZLVLJdJkF80qiDWS3vvB6fJcL30X8e2Dd
zS0bJsIswYgd9WaxoYN5P+GSHXkCIVio8gwd4eU/chT0v7hvo0G40eltorJtUeji
Qz7UV1oUFQNbrQu11J+lnkIuk3YK5vU++HGnXgXjZ4OWXag/CyIWjG6j6SinTlWO
OlPOOvwk2rQPEzYstuW223Jp7VnhP25WnnLgms5Knj+sNRIm+hv+mOdSt8Sb1T78
Qn5PlL8VKLJP8+N9vWUx6pymXnUGltmLLt9lbFKqNWi8S38TnsHwgFKioR2hCzWm
y+2Qzhduy1VZ+0DK0dlCzCSqmvcgzYwtYKdbP/U5cwXq0/kN4WGinNgKoYd6EBOA
K/36shxIIirNzECLW3ZtqjuHMn1BUfwEbPE2Zs7euuQu0CZdwvGUvizx8uinFt2G
ZAIzc9yf86+dC+A+pBE2O8uhPF+n1/2EiNFwyh2EB9FwrfEvkfgyWlmd6Ll+a/WB
RrSwhlZXifkz7d0ZYullRV2MR5gO6ujufVq2IPbHyMcQqkdPlTKdO1Q0eCDbajlZ
S4bZWsZ0Hjm5lVvxS4kiCKlM6X3YISU0nat4aUu/L66BEuYyZAv2vpffdqgVx8Ok
eG0uxwEiyFIrSh0xBJ7qgqE0e76CxmJqDzBUIwa08KiJO1hAoKhlcw3KDPWbyurr
clfydU/LpVFAnLjmlkR/YNQZrG1cwVBJw/woRe7SL6dnsZ9JxvsCDcE0l5OmI+ie
lD2NCNmw4a8dHI8fxuC2bdpWPp8aPzk6dn+lv0ckV4bueBwwX20kzotReD2l4aA6
2gX9OWT1+96V0TGYV/xqkelfum99jFqAI0aT4WnFgtdDsgZurbO+epvTm2DM4MgK
0IBAFHV5YKVKHj83DLAr4Gmc6WbQFBsH+BBNLi5ozJv0kw99KiyXKzrdBBV5UIpd
haqE4LDQQY6qANTJ6MIJ1JH+3KzzLSsMz9S2HMo5vqP2DfEcbiE4sRTIJJBvkPmR
So3VG0ZTH24fzP8+bLkMj6Irgh4TvCtrdbx75bx23rc6Hu5kb/otHqo5D0G97bZg
9okqN4fQxJCppcVwRs5pEpG7Xx3SbBiuqXVPK63pGpuJIyuQ5eyojZanA3CuUaiZ
fv5yE2/NQm8jYdHR2+CSr8PX8sOBzdeiJoy/oVXBmZwv+wAiyQOk7hOtBF68oCqo
d6+ex5G7ofPEhfw5TdeOwiLCJw55skPDGAC1vU3kANkqQliHAr0zakaWjEp8DMGd
1nLiyghagt9cQhcMPDHzTE7Kb7FWA/zGN1h24RZHGiZV1gKN+XRMYMRRjfCHIn1R
tmqosPQrbAKNH4KnSdLEe1fmGYRSAPujpUB59CQ2ybovpDVBSTAQAEpxNfsGHwAY
CIvthOqlrKrA691yrMDaiVF23ZiJFdt4GROTWKIbDCS2tI7lcZSs9xBdbXxGKbRW
nJv19NEatkAIW/7EuvACNdNpkH7/L+NjQUD2hY5LZ05EuB8wk1pKTQ2WZAGSwVh8
/irPYn+pbVcBmiIhGaiWnIqI7Zket81up/HbjZ8NrhmtfcjccJczKiPICJcUjsrF
BnUlivBNif2sRzMTARK+fwXPiPU62/yglK7RMaU4cs0ehJ9Yh9p3rtmu0Y5lK34u
DFk9l9IUnhEv8glZcjvQ7aUuk7or12Yom8sTk4MgY4AMn0SaBsS7eo7ScRR2Wrv4
36jpmqbYkSuMWifKp1nanmRIbemw6P6rPsbMLkjuZQeX7BK5fKQfjBugmEw8YD72
VAu+2CddkhzoTx/HfmyZeN0KJ/KTXB6mUnwkPLZFUbZzfoIisUpO/dKMAKVW5rEQ
k6yGN+L66EKd4Hyrz/V0eI1t9f+jtLd/eTgf/paRewMqpTcLLpTon/NMSUm1NdeI
jcBuuoQdMU381IPelviWTzIrj/WQPfPMlpbZaBbYl3HfHcr2fUFPJkPsk1NroKpn
NM8Inwew6yD0cJMEInnwZzs1W8YIEePAzh2CRsgnESJYmaB8TlJ979q1zbIsTvjx
O0xp2GJ8O48J2aAD/3IZJukxPnNsgz4y4iI+bp8LilhBYz900v2pBnMjNiGOL4UZ
Jej9bBgSNR47+0jWyzl33sT3M3ys/+0gVX9BPWikFGlIUo/gHFiG5C0ewyp4XEu8
+0q0+bcigzTLxRb59ipYS4z4jSE+KkJIED3Grd0yRf1MXm2uraviXNTrPiejZlr8
yvfUVot92K+YGUyAmnf6/+CeL7pO3urwTWZJV8zlCMJNTH7kAldEkanuCIiAodhr
ocYKTLhcccrPD+6ijDmwaUvsj8r1GtdhtHtDh+lIZpKi2DAijF1LxBiddm2QL5nK
uMzj+Br8qVZU+KuVAcpqHJe7N4MugvNjM15QF1VFUQDLZIBzuMnWtEVwkRJa0wyM
w35I7fhIRu48kAarrTXfvKb9+jCHYuDBg05/2JaHejpYEYpkHy1Hj70KbTWBCpPL
pwfK60HfUsUP1RibfMAqs8GbwdzaB6q2Gac+lKS4+zxoxeOSkSIN+WY8UBZ065Qq
dE9vkcki781DmcWzvkAb1Z2qT1QSZwJHqegbjnIgfu+EHtUcuFsggF2ZbGhWYe1x
6XH9hvHj3+sgUjJrZ0mmt0vowaBB21AX3DTbu64QnZhEHZdhkakrPfqlepz6HbJ5
1PZ6AIcdrT3B28+x35zlaPpH43RNdHTeu/SrWdGzkCCXcbsXz9ZfdX7LBw2imTLj
qSyDosiRO4EWQcJlxPbi0Ye8kMmXcfW/AjZPotFPit+Q02+ZxgJl4rwlAH9fNaaa
PExr+u3l1xnD2/acy7vmsL9GY0j5tuYgXdqTbnBxkIT3d61AUEqldG8JKkQYyr/H
B19aI7gb7/pnj92m1R/+hD9E04YgLwqUUJpdyD5cgp2qpql3TjwQ9ZuWDKZ1ejEZ
2Z76iLcnN1DxGGFEApwRB6yDQzfqAtjyzrzO1EOoqIyeHxR7V2O+m+yx5z4vUsp3
UNIA9OhtI+voCQTS3VVCgGZ/p0IaP2Q1cOMxRGKatnO4NqjDCX0ekN/4zr8MIMHI
URZy+VdDehguG5uqv4K2wWzU94KlElgqFvZpZLIW4rdquC4wKUhzmKfJXoVIlTav
bJ4J6csmdk5KxCpCqKu6UY1mkxParAWgEKhpw1K4F1IZfpZxFp97m36ud0yaqstV
TwqeeipzWkevZlyvkqfe6INiH9ikK30OYqP+xmdOKLgni/suYNg/psXNxpKbs8/E
ZEaWitMTm1KeY0NkjmPNSuIyDEOnIla/ddqOUvLhEZiP+gkbKH1yFm3YxMpt9I1c
XyZpzJTW0g/9NYh3L5cbo94lCJ07BKoq9thCsebu45KOZv6NV/6y4nWQ6zFGGQ/Q
iC8pjurpsDhkK3vf6xjMlFYi9U/eE7MQDTK8Jv4sGm3+VYEAC4Bd4WlAaUDEcwJa
aBuQKJ+aXRAYQH/secbWDmqyLSmtZ/X3aZaXPRiO1dY7m8nVrPL9z2MC1jbWr+hU
TJ2Q0WEVLRSdW4kFGFG3y3BrQLonxeQOBIXm5aY9I9Nresd4nvix0lLo06UaMYV6
bHKSGYYaehSnnnJzTPinUAVxSQ3rZydtSoD10R7cN0AiQq7F8LZb9zIt57Sh9maW
rkp4fGitgTcaQNsCAfcZUA4T54eipfKH5biWXND0I+8m4DRbgu/F1IZSBLlm8lhU
AHAd7fN00LvYw/CezEYWqvJxRv6OkCqyyVAtfkqAKwKTrRuM0tCGBdgoNr621G/T
Bs0mVup2khCFtcwkoqNjhVFmOJydMy23Mz96l7+mG2OSi7AFRoQwqODsztXVC3c3
mmuqqnREsldyFWhxIe/D8m/rKZQBqy/53BvHUrSe0LHlLAKUu49ZdcrjhGgk4zpV
9d9azzincV4NFJcY9Hed7MtqCAj6TKvu2UZ3nIbVh+yqcV4oaWZySUYcG9hai+NQ
O1ZclCWYc6wP8hkO7EEMipi6ly+hR1jAqbMN9I88Bekb+69EOG4sn+j1ORCYZF1Y
X9ELX+7MxY7J5ogarPz9365dRYcGrBTlh4KiuqUqvHBnIjMZ/fl1HjZ71hyuMWJ4
jSeXwn9izCHAN88aJw8ZZR2rmWRAkEfme68+t8ljfuZz0B5xYUwyRKajuf4WDG70
pB1ENus0bKyyBbBnPg+0fAVwZPTluS/PXzzq90QiHgsD/PaQat2s9gOaviRN9V+a
W0ggiwFHTJGzp54YwynTW6fC3hr1Wdgtr8TxTvGt6uSELRkPuFXQcLqzaMrAlhaS
bUawhTCGqOGeQbQ8p0zyQxPazWuE26YMH/gCIVMMFR9W/0hGvkW/SHWyRpc6YZhY
qyIH88jGMzZ6C8RTRztHHVwDQ23MvdN8nQQ/fPVdfWZgbMQejm3fzk3hkljZBie0
mZFOO3ggrIPaWC8YBoCEoIRRHkhDS1RhhuQY5buyZE3v7oaavWOXTPI1S1hTxrop
Y+InJTI4vvy6uX25cPauJKqF/hdiGX+5AvfHRjEW/V7u1ptaqXT2bOqoC1bB+kXK
3FddrINJyT+sGmZxyxLe9KLFVU1DmLjKW7PpUZsrDhhFpqZmTS/izP1auL/LxZhy
yeeL2vKs2a0aZ97nyODxta8D1DCs8Le3VNCp64ObDxhdIefhlW5w9G/izJ2435AG
OCqg/RZZxAGWQhIPhGq1Mbi4Ys7woHWVmGLCM/rZMNO9hMhgT3BDILcOUI9MLmsn
sLDuawhjXVKP38r14fmc1k9+kKYnku7Dk1kswcHaGkQYrnnFilrypdiBLf4c6Kyu
LnT4SkbMGqvEFj1+qSRfRSFYNBZ72q5QD5gnAnAR58h4tywgC8VwFBUlAbCtc7kv
wX3vedquZzc1hK3wAA0y6E53SSi/NJtKspEtNvGaXyGbupEWClRj7AQ7c7lhPzgi
zb2jmf3SmtPyT87bZY525SddKNxQ+7EygSdeijH/KzecyDp4KMyxk4R49Bju4DX/
kPE7FG41Kmm4QCReREQd8PyJW9YZidWx1Qq1emZfBCA5g68txEbwcMJtMHcguVeM
yM/TBL/d/lFyNB0lcpyqhL5wSCF2evLgVSLTZ0vQqcbLLnJZ1cc+M0U8yelGGbyC
NXlbFPWRDUrDHUMy3Sgw/ZsdNjZ9Kn6oq0Vt4bXMntWksSyriNLK+ESoACXAwVWu
rZ6Ayn9WWBubei93JKW2xqjCtKZz7RXP9/JbD4k6NOfD36wxKQIhkpzT37Sje9se
TDwHCWDtOSb/q5HI+8aRXdjb7g8HltgueWjqcassnOxLlQcm09j40H00LD7ASpiA
KWTBC4tI0tUVvVqOIlfzDoux3pJBvyU4GXi9iSt+fZhb/6bAVXf1dVD2Z36GWl5a
qb5TaN7tWy9Lgrq3OeT5weDHCvpm/NXqX5KJt1pU5EkZwFvQIOP+tw3B4XARBzY8
CnuvR8yG2NV8awn1FX0UWlEbGWDAEeUxPCOANSQLlSssMgXzsNmjpZrXkdlNRB3H
XV2GkhxV10WWUGuTSgbrvrzu4zwHBkkUPeGahVvVYzvRil3mNlGCRIrKL7dgB4iA
DiK2IKSYJ5ntd55Kd76CWk4p1cFHdxMCJki6zHZxYvxl19Ao8ha8lV5R42aqDXZ4
BChW9o6ZhzcGcRZaIH4wz+Xq+jofm/v40MPKeA8qwKjI6P39hqxsbmrOgGSAGJOB
4cJOjjWKwNtlu2qSh6MCHjcX2TJJqYlC22TC0tOPMni6lFTIxEK7kClxpZ4wE9q+
8+d08+NgMeWrz7RbeHNvBGv3jvPCrsMZXoYaz3S6zWAGZq/aaE1yYOcJZoq2acng
AzOGpabCF0+nEZfqrfUYwCV90bU3Yx0HiUSMlHqTPfw3QnsaNQku523anvJpfnQD
ykcZSIyDqzPhZ6aCXcH5GSkjeWkSJWwNo8DUP7xWPvDldW2ZdDvUL/1p5vLco6SS
nbFUBo7V4hfSl+BqbHJo1lUAUdUfCjWW7i5XgmjWbrYm95+KMU3OtLCJzpNDREIR
r52xlnWTf0PKOxaspWWuX8d9kcDvnzAjPbjyE3ASQgcD5mF3aUGOAOabg0EFnhw0
P5TDkIXPSvUWqXeG9+eGIc0VBNqc5TLeVasId9IZwzxsC23Zki6KEH+uyFEkmv6U
5X1eIRUFvs1hIoWOWzI4/An6a+ew8vDniXa9lkKId1MSt4JIMZQ2smRj5fki1ns4
8HKCPy2G9hEzdkGEL72RkTE8Vlo94+uWmdSM5eehVFDLDHXrbUEnxdsCfV5j7/A3
t91UxW/q8nafj1oFakLS4YWCvhRM4kaEOU1ElbMyyOPbLw+wHQAk/zuqWAOSlxL4
B3zdFQdt2AmagKvp9LvRmfdROeGxpG7CGHORmlswqcUUnLnnR/lYywmc7fQeHimz
J6HMhmO1+H7nT49Xca561EtLvoSdlAEDtRg0mm0hzQRvlBvRq41jxODhSUC8PHVE
q4xe+vS6Rh05rkKONQB/vRoR22HBoPxt7HiRZfE35XN/+410QK3TxfQsBYd/FYt4
uAGeaW/wLnAmSRiG5Sk3TNjVXnYnlyCOwLSNwXuib1AyYGL9E0AhjF1RnHqEPvcH
ErLVx3yCHk/uLjFANONNWy7fkWG03Okgg0ZGLjOmlf2uu0diU3Z63NKTyWSfDqkx
hydwhaHIUX61ku2j5Mz3i/RCP4yKSzVBDVLI0MzGeqhsl8ly0Db/GPMbr6vZVClt
oj1oFZ+qR8oux0KCC6ZB+NjO+iH5XZ/pF3CaIr9S1lfqD+UNzTpRjHv8ZbsrGdFd
9al8hek4HsDl9Wbnf0yxrpwfYqDK9/mXt3btU0OIBuI1y3fnWftPTopcTv0HjOJH
TEnHu3UUTaLUuF5reKBsI15tBbrfgSGAB3WrpGU3BQBmF/wJV6K+JEvpW88dXS98
XINuk7nXYswi3e/CDfqj+hqvnuwVhc7DBymfrua0n0GW3YM4+9pTA88arnU5QjTK
NCegxkgE4AbzINoUcTzFN5zVaJDpM9/iFx2JkBusrXt4DzT/i7kXagJZs45oXUFW
RmLfzNrUosghdyXOj8weBhP2R8ZD8dvLZDiLSz7C5yLAXt25qxnM3ls3ICBC/Aqf
bL77NqvRhF7+2VNJ/RxzswSgt7+wU80chTpL11mqwyFJO0/CcHiiNkUoVZqASET7
5fITuX8hlF0ZaJCUy9b5Iz3kMeJIAoh5X/j95sZDomhoKuv0Mf8Iwm/seKfqqEIO
ldj7DNCwg14VaDQs3PM0zDrL/Nd768S+sD8lrvlyie/rH8Wwis9QuDX/KFYW7lUH
G52C4L1uc9c1Gu99+brL/fxcn0I0zvhYNoYxJ4KNYIcRVkhfzuuEHRLyhMpAn9K4
HUWBTWOoLBkIBraFWnoQyOyimS/dMh0O54I7y/Ra4KVz9iGxwgPSJj41oTvl12gg
57B9oONF12aP1RS3QiLTPGhTsZTi3C/X9HOSEX2FiURmyyZIsJppCkvH4dnjquJA
aoSxnqdimz9DqwhSLceUmVPa00AeFCDY8C967HOAHS0N/z56jchhzX7W8RTn6qFC
+ypSvAUSWVJUrc1dz0zMnEIjGtrJUq8i2PElXENu49ODBmrl/sxTlSYcr1i6m7UY
sQtLB1f9ua12hNSKqCDx0eP46+JDn2regIo+HSaf4RBeECjYK6y/PB0b48M37r0D
SWqR0V8bhjV1dygC/N6PGthlu+hDKYVpxzNq3UHdd86Mt0pT9SYdTuYz5MqUd7HL
7o+GfugP0A14reTo319MRqIoIm0nVF66b2d/6UbER14PqKwjPUdo5C39BneCeRvU
5jcwICvTA1G0WqlDIBt/BtXZzl+SUywyf+AhNImIuSV9m0UJeqD9uRFdwVL7/Q17
26CSSbu1r4Eax1eN8tzzaK2Q1IQsPtH4GSZncN23S49t/31tp8IwhBj/jQ4hbyUK
wO1LSLzc3MVv4k/B7mp+ESHiwUNKy9xXEj4NVOVToC0RUFhdiCJvjI0rYExGndaZ
AxTglwc1dPPgfrCayC2xRdvP8PEIbzncbop6KFGbaDgKIlptk7PsC6HPeSeOojSx
rhNma+vAFQuHXEjfVTGpcfRbJkkq5OJkQxmarLXZFqTt796J7IHGR5am3f14KPDw
jon7yp6RPZ0cwcW6ZfJ66hSVdJ8WxscFb8tAxTKCoMDmGIuHXsg8Xw+A9hC0T0iv
i1n04sQLHmzdzwueKuCm8HcDgN+F7lmQk9enqg34ihY4BmNhhqCDg0l8T7rxsRyC
R7RB6SKFj9cMVnDuBBhHLiZ7QRRu/vI0TLpJ7dMTvGA2EvlbsG6nhSf5M927rg9H
KMyAAFvuWZKzJcspTr05FBrlEu9slIIrTc9DGfZURHMdkhZXSh3ZLJXVn+HBnkMq
espKgALB2Vnni/mCxCkn9zrMc0+Fe5OVWe6pyuZyIff+wPbn5E5PB2DXzIOxx8R3
I12SNEaPnH+LaVkl4c2Kj5CoJkhVt2cA97ta5oIwGVuODJcgLql+Va/8jmDL0CV1
Wu5pEKwMcHMCyJ6p2S4p405snlfnx+nHHKircAR1cznEXghU3Yhd27vIWVzyCYik
nHQ7nQGE7cSAi29IVPD21LWP39aId4fpmyrD7b0Ehx+ORbasiO3POSWPRyTbvZVX
tvHw7nITqlIx9zuJ2abZ0Wu6OXBbWLKLV24j5G+mZka8Rkygep4whJ6fx/iSNqK8
fG4Yk2jh3ZoFHm5VWRlK03cMnOyos/z6BYJBDG/cPlQHNJ3ePKNWyOs1Tc5hDIin
DwMLWBFP7w9v97ReDs/PE0sLftRP9hsftdAL8wOYDxAX+60rK2J+koPH2+Xu3+Uv
F1gHsBiLwkHVNjZIjzDf1GFtvAlNT7Jifs4So2yXUaEEbJwy+0RBdg6W8F9IfGwY
yQZ9g9oH2RXdyroe5THPon5Sw1gP/qVC2Rhmm/VLzzsLclJv/Hse8Tbks7zHaHHl
o3z1a4nZPytll9T2z7wwrg9agZWCIPBkCincbHpOuFFYVBGrBoK3B1Wzo1/mfyyF
Vyn7i0MSSV5xmfLQiXjYSnaTyTSPT9nLWGpM97zok0PTtuBWEbjOSbgPbvfyxPqf
7MNjI4BHgF9u1H91no5EyHdm3h5yvnU859TZaLYTpDKzBwp/S3sYSIHqioqg9g18
Refk/EMS/7NwBS/dud7aG/IZinkTn1lLKatQ6KjUFC9n86266bgJjuiLnhhmO9Q+
STDmbODouDxJGKtTbRgSlY7rkJeqkPEpmHFBpuBgX3U4aWvHN4Jti4DmcIVFySUQ
EVKrphuj8/m3nrDkdfBfmgekWrR8Ih4aRR6yaBeL8xBygTHsp8GmIUb+NsEYSueT
t2+bDBHQDMeqXoOGSN+bQeXJb3OhVHI/Cnxo2RmXkEzCOW7FVLORssl+Jt5umL7k
p2TJhIFPe9DFGH3UAirvDbTieqYPZfDXXhZb6OQNRmdmr0GfKyfWr9IrObZcOxdX
qhMIKXqHrY18cm0sOXc/bt2F9CcasHMOVR4pwUyiGNq6wEOwgcoyJ9L/WO+GzTbQ
vBzZKpytIv22xyNLariGySwZFTeoGQ5yrYwvclSuHJrijnNDdgGl3bMVqr1LDQVK
hlC1DWZTpvqH2rKpofAMNT2qi8t39G3BR5vlr3zanPod9fLcNYV2Ay7lgK/6dWmm
ZKWipzTQzjM9SIBbRijz4y8gHZ+r1fXLzWtKZwxYgepZQdrapk7p0q4og08kcNKu
cK0+aYPmUxMBf12QbuDHUyf+iuSuhDnCqal9rhnKYJokILowqAbZPs5s6X10ph2H
+2hCheYnnaLcHz/w9JG0skBVKDvLzn058qIGJDpW5fH5ibiyw62Isy/CMNfI8hYb
csp9L3bBPOmNcTlG5IWuXNi5mPYimEnU7iK1rT5JCQ3TS9FME6s434MVsnZKsh6v
yTXjJwjIw72oFTG7R8By+JTV+rzRNPUl/De9AEWsLzxxhYV4w7tkhxOLLWrzia0e
byAqc64aZNfEXpqep6vpfW8tNcgPxayotcpuv6bEfByu+2KNmnlnolxkqErI26vD
Rg/HnpE2mkN5FfCrWE3d+Hj2ix1GNzUB6cjfWtHKPn5fIhdjQhxh1KpQ2VNx1vuq
N4p0RcH77ohJMAnjJNczB+vqeRgHNVDhNzhzPYRk/WNlPEma9VXarAIon0wPzHfe
Xf1vY4UMD3EgKwME+mnFsmy0w+71rnUuqQxgR93ZDVhKQzK5CkU4pUC/rqUh/vPF
A+hbPjRsjOH0gLa2I2O/CGU/WkU50QNBU57StHu/oJRjfd49s2+EnU3dexMrSwmv
hxZPKFpDR7TAP+gNSE4oBRqFkJPqZBR4i6/8m0nUnJ46AzBDPxz/6dOtdy2rEt14
ywkrz1aNV5Cm+xTN8XpmOe8htXutOwHhJKBFT7haK6GBnpql4MWzWrPpamSfT5kl
Z8kgQ9xlk/YLGCyoyu8a6TGXy7qvSpWkt//A5ojAfaXvLIfcIEggew8sCMw8AUf5
qgKE/7cV4qSttS46nEOzoQI+pOzP+tgoP6DErr5IkanjR2VCJYbaYWu1Wjovham2
o+P4Yim2xDITcgEAW5YaDAx5LBEBRSmtyBzBRrrfuiAraGBBDTLoiGyudpS3KLVW
XWRDN6ckdPAto6GvXUNURxUJpfQpgePFD1dUS5YQDAbttuw/XXvae3ksCSMEQYam
ty98UFZcEDlzGSxMDR5R4wtYa/tKdxSKYz11eI5gsscAIWaw2VzNlVu7ikEjvAL5
oFgVJ94vHZwQs4k2KLQsPDdcD5KiEYLuqG1gDFc+6wj4zwO6+kesrjfDl6hrmbSL
s3532I2W4pOdr0+sDHGAbiLLxoldlIhVEvXsOYq34VeIw2p5b/C11e3hKtz5nQQ0
y1kduyUwOdSiUKugdBqM6OdJvj/49GwsMWr/Qz7dBoAnEgJ2RcYj4hgtqI83ACRS
asAAGWduuzzy08M4W5eZYI/X/HBjL9gvuX/QR75y9UA373k85ZUY/2aqQ+dzd5a4
6VmYKOUUHMqOcPvGyrs9JbIUmBVm/BNAPY+hewZehAryCzKogQq9+wr7h/Q3OE0Z
HzbOsKf20PoM6CCu9vj9VDDVA0QV6BEWnjnBnYE2P5dxO3L1AXGPwfsuxMY9Sdwd
gUDoaDwrvLu0iVonexR8pQ1bGMR9ZpIKBPbiKHzdnVQHCZe4emp5c5rL6qXdt2MV
qn4lt4a1w5chQfUG3TlSoeOyX09G6aFR1ee8uhAgarqDdzzscoHdJF09qh/aI8Sf
gTfO3lUKwOeln8v2kBNIV4+y/65FlOFZ2chVqbfhY4Pe7Nh9uLi9YFK+OSBCX6Dh
OmL7pq8pM3e5wdpEVxPe/IjJ4fDv2me7O92NsAWGLubwGpcZBSaDJp8z8ecnyyVi
5ukAxGzWQwtoiQQYhZe+bAg11nfZOaIpm/CwsRgrp8VIHmn4tnsRJUrmtSuBCkoP
WMCzoLKHdBgRrg0U4a315WvWloo0f2CCqKyxZ6iYpGb8TDO4CcY+izNHsLMEWtV5
ijM8ZPt4R3ozaTs+XBzMnlPE19vxZD0rYHZer3WtZ196RcGWli88GSbwbV810Ds1
/E9ZFEI+HbD8hXRkHZcaOkAqO/2zl6ffLT/z7voV67xY8DNKZ5PhymjoquKNTXDz
8ItNmaa3mokEJHT6HWU8mpASKDNXUFmwfxzXNKQOiok7QqxJQ7prR+m2SYm56aT0
AKsSX2WO7fwF7PX4pV/Wdmnkrkx6+zRYovko+C9VU/s9f3vyvf8grttTuWiOD20t
HmfttkP5WGXk7Hup3zEDw9aS/jWvpnw6Cp8I6B6V/U9mlqzbHfERcblG0c4za0jt
O2yU7NGdI2cWfyb53oxc7rQMc2g1CVnhwFhWii9pROxnP5UXKaXeHPKFwUg5u/3Q
hnAbN6OZ6zpWP0ub80byxEjk0QtMk7RofnlGobWLv2ltVMvITQzxw22Va1RRbkkr
P2UMTnKy6SX9ZsFEOeXc2GDoC/BKFnn5/30saGV1wk8wJEse1j8i85SL/n0QonoH
nSgVUFg3YnKkykduANlfUBZjOYitp6gbr3LuEmIbZjttd8qk5OcclcSgJ27+bwV8
IMZsoM8CxganipS++VAcG78YcT0CIJ6TXPvLjf17zEFiU7ZxyTDveG1BzycduY8p
LQ6/Y5GskKwsTR/n85YsrvCnVCzI2Oi1kHe3tqecB/B0JB1hQWjiCaz8dXlaOVbj
rOBms0a+Hu+QglxAYbA2D3zKKpP7bCx0ss4Ic+H3bQfNdrO49sZp0c1RTDRrICyl
qljUU7AIi1fwo94+re4Vas/XP10B21PS3tN9w5KjO1wkQ3k0xN4OEqxGQgcYVyfY
RHiaK9tvw4tI3HxHyo8KHTUqFQvAublnvrJUFIwfN2YO+GXAl1Y9OqeIJs+sfBU6
CmDdedJGVwX+qU4VAxKyjfAX2du6TDcEz5LvPJqW3NpjRRjZcDyf1cliMIB53e+T
rgkQfcId1W2B6V/63mi99pjLTyaslA8uTvEF9ZVH/99OgPMBAVzE/TmJ4y/9hxYH
lOMwjrJHVH8G7hdR3zmb1e9/3CizMeArRdK46RTHaHUABleCfRoNpm6hzHO9PCSQ
xFuCM+ECY16QrfCdwYwm6MwQbYglOSRg91oeZEg4CZwAK0MGjCmqKKRPgjt4XFmg
RxN9w98noAhojZNCISNoZqgSONP88bl4vu22WQ/3YF7ziyWrKRVaGfzsk8i78bYF
JQGu5dBmVrzBt591/eapeSnPn/ikP+6lCCBmpvpY/FJM79TyLzz9S9GxEaRQ5pam
4/kJLJZvCb7sdKkN5y5dOpAuqXu/DC6MAxlUrQ4Ba73rShoUNm7cI9Hh4n91X5nz
4QJhw9gTcb6P0l4f3YAeAiolcKJS/Wy+gaCtLgAwdfX0M08ddJT7lFFD8ZxuE1vj
y6qHFruAk13sLe6vN/9szr7jn0+gXyIGBnFrHeACqXtSblzq6KqY0N002+PG8XXu
N09f2WmlA0bBO33JN8dglP90mNgOdHTE4DcBBE0gADwgajs3UWc3+FmP82EXPBWs
PSxIMQ29tOHlw14bTDSTTAKhiBD+UM6nnY5eTFJiYNb7iLzTloDj+yOl+HeJ9+kZ
yKdYyDKiegeiyyjS0v8a8MyZqC7kRENmkTZIBUIU3NUbQVgunkh/fXJxMqrDK6XB
HtIhhGbHFdTzUiYNkWWBJefs6IxEtbxTkqhuC9zFNMqiJPuc58VEDAF8qHSXC40C
mooESJR/dRiJrqnanQz5aexRlfAqYu72NrhY1Vw3GR+r2hOm6kPMRDSYidnmX2tx
9+Mtwmldt34K4racTPisDXB8/JdWXe14BV/QgxFreOpb4quL9nLTVpDdKIMKwRo7
KVT8Kn32MajaDf93lBnKNAfY5b76V1Dc/EYLFq/LZkUST+f8uAmLCLPJEJwj3JK4
U0z+0WwHU8nNg+Gk9L8XABMMB/mIUfsOFxZG+rh/IsAhauKojjsLGsK2P5Knl9mu
C0MsrxxqxpL25hSa9ketgOnlcwdx4nAdh3FK4pnugX+caNeufmDJ/ESONQ1ETN8m
VhqObiJONY5cB/HTjbiigMSXCLj8N8YTNr99hrzNoSA8ip2JNV79qDlBBaq1kKcD
h/mKTKyxKMUu1+6Bu7bSCmAP17oUGQC61Ig/W+Tj6R0G0YBYfoiWxm5uBLB+VZ3A
YZz/rEY4FUT6j15eFKuTnzoCCmOZsJZEKYqIwgNlI/ljUfDDq5nRwnf53C9YqgKv
0TPJRsTLGP2X2eS6JWJs5OmkMeGYTAPh9Ky35ifxZS7KA3LgBAC2FtUsMrVUtsvP
g+riGSzLclGpK/b3/84OvEr6DmiLlgDjS2frNyphJkGSZIuVfafnns7W5V159w7B
moc9QCsY4Y0GFwuF/WqXoHPDjbkOyUaRkPsY2igfpqGBZkwVIZCtZsuMfNNpTv8z
g+aMt7SiqagAmSGPFRjO7bdIJIsmZxCuN4SW4LSxtpH6jRw/fzmD/lp7Az0EzE+1
lYRTdJPYc0FHIjr5hek9mUun9qfqtTetJXOneqQ95xk1OS7SXJOaxeXvlQSKZimX
l85xc3dy2pnBajA2J0o8OWjR6Fbv0Dz21dZVeuzhTAcEd07Wxc2526qyxv30FLhl
n2SwaWxSzUOTf0+gAKmOs36kFRJF/xvopjrlrvY2cKxov30Va3MQ44KsmqUFJhBC
trxBmcs2b8sRrBMamBWchws7E+FBo2ZSBxPvVwaqIQRViYBQro0FCCTe4Z7wXH2f
003iQyz7qi6JMDB+kKj+Q8z6fRcX4yd0aLnHqrHmeaqZJvdrQ+SZeNhp3/3G6HPr
FInskFXbngFpxijfhg4fVYYrD9iTARgSvTRRDl9S6fbBMb4i305wzVgiNdZHP5z8
KDQaTRvoamOrt/uDPo9k0Lvryv5MFDF8ouinyOnmV7EZOmJNaGKAvwif78YInY4G
QEfB/jb8oYLsDYstrzuiuHdtoHUTrwYc4BH8fn/fhxrtyqwYIoM8Q00+rMMigPbG
Bq5wsu1Qm9cXZ15UeRDeHT62Rd2WHFw3yL3IPnx5PmRvntsljcT27h+gDixOAhAL
Dv33Wc9gPJFDbhBUNjdjAJZR0SFfYhuYuXihED54LCNS+66u8TcoFZ8sECCt/PLz
dIYmPM5yDcvH7grBvGhCnerg14shAZBE/Erwjy+7LBcqvFPKwBAfOSJQVG0xUbrH
cCwX66ubxY8pqIQCLstWwk1Dml2NeEucAhvVGdfmYhpC+CR/VRLpNoz1fE6qi9Us
0J7cIlgub6sPbuc+6KaeOowKu67ETbqVYPztxXVH+qSgURcTGIKA9ebj50HdTPsf
EkkqbeGvQWjZzw/3Xm0kSNKteQ4WYtaGAW0Fm227AnElg6TX2xUdOtzEG8B+q4X2
cO7qTNlDO0eLGqRUYte+uyyWTlUFwiygiILEgdol7y3L0TXoJg53Xy0EeGE/0g39
1OoG7kpQzr9tU639p3xrZEAZZacWdiuQxfPBJaqQh99DozZU+Og93UPtnEy9yMYW
XwFi1nKqdRMzWMbhLiX4+/0vNbBXBIY5TRP2EbaEzbZ5Vh970qmz86UwuYQr9NV6
ak4LLEt0ZzWb7sAaSfiSwzU2oohVD0mpVip3nGUIrDVLqrTAZ0p4WSXnaJ3CW2ZR
j3Vg5FXugzPcxGgHkrouJx40nT405jCczbQh2h4zwi3pxkYeRSHNivyUfeCoWCBi
53hIskR/sGDoGq/3jbK86Kl7aPUs96gvJrRZ8DjqRzchFqtWwEEofE0VUlGOBgIw
DEW0rjcDLeklafJG86qLNN9Yh6xWpFX8fXBCq4Rsr12voDj3xMEM+cF0Cdm/LBFM
EexkyEHesxIK4BJyi+4QyCVma9D2R+yVj2M37FpqYIm69WN0PbgqNCrtybfozUZk
pGtiL4RG66hXLSi5Cn9+iA1ZGwj0u7U6Q7WaKwU4XdijI74biLFRwVDb1A3HlnRQ
MOulHVRS4jxaQnhedyMn3ufpHDVOWGL73QFB6bjGszcJL+2rJEfbWeXCIBKxCFdt
wbUBvptNtTyLOjH7FTFz8KfYcf4tAcHE4NQqmhjMgou4S77whzKDBnVOWjsM717F
74/GqjfZmmLrk0Vp8LvnDipxJNQG/aqGkG9PLU5a3iUOrg9PkFNDsMzA0aa3oJ0y
lbWuhno5T0+E0p89lSV8VVl9wwgk4cQAD5TeP61VR/qL2mDS4O4s5HPaCCUO2f0k
DY4KHmUaJlo95cjbkWaAgXusWoR6SB3aAfy84yS7JUbmqq/EWC3TFRYTJSgVEqXH
qokXyrxyaG1ePNHxOmrH3hQ5ak9CLI7J1f78+dKHmHJc/uWY+OYi4qQQGzqRWawr
Jn5tPMse7vjfwRephX1nodOygjyxEHGJkhKUmLI+tgXQgYneKDXHMR4KL8+Ev2vc
uYdAc0kJeiai6ixyczN3hfZU6H9U5mNv9pyPWrqbECywvK7u0YjUBELc7s4Y1hJx
Z/QS2xxIUBRIZNjYDuJdAYuEnuRWy8vBO0b2ONtKF8znaE6g/ck+VbBmB6TWeUVl
qD9PQ4yQHj4Ppi20zDUVbJL6Qy2Ix6BS8DGoH+l5KuBp9L2t/XuPuNucORO5va+2
zHj+TXdDbyY7rHc4Mh+h9Kcy/JU9p9dDuFk0rqQA87IADfgPS08xBPoj6+q9kPaZ
SIuZNX8rPw+pUwF4AXBGG478H9Pg3e+ZYMuZFWEefGU3B7rPX7oUNWGNBVbLRrwy
G4oQX9QA4uQtIG9KVwwkLilngDfiYffk3smx5pwACrdzWsIwCk2LRcmUYO0M9ucO
eH7vrz614zDqdnq/CLVoV1h1c1imjNZfsUk142JsmVAiofIpzSdidhRsTm8Qp3Ua
SAH++cyPs3Qemu0hWcc2ujbAFbycH6N3kJIsuu45SEvOfrGuenEugEAxMsreW5Ci
gepzEvzmqbhYo5MhvF1367gYqmGHveRTLTX4DNk8DA8WVdXbEaVLwy6H/iDnnnpw
dlsk+Fjpdg27kvU9o6c/WKi9Zn2U6gVqXtlOvVbqjbxD6uRqV3eWNdFHcUE5rJpc
7P12yw25c2b1bNt84vtdPzHCR9O8zKXaPyhX+Rfg/SdOvvUsTYgMGX+0YH9vcKgX
xNbr2xb7K8oPcHrwkGgcK67hiVlvis0qYofCFEGUyGB1+4AVR7j875vVLoKAqraG
4z2ATVEvrYGCVuoM/ODawawfFiW1uPyTLVjmpJ6bJC/7ux2O1CVfZYznHWF3HqBk
BgbL2X3jXM/w2IadnQMr4L1ULdFZdFHRp1ykmE6/UeuP6oAdEGqc9TreOFVaOO3I
sYq7eCCLW7Jg9/O5ipwmdZXNSw/kSD36kqi9hxPSrJnCC4yaIr2dKbppBW2tSXY4
azwHfecUEYiyVV6m0lwvWMPkwZkVOou//WKl9mYc/nurVTu++f2vHw0tNWJz7jba
IHcoeUlVAYKrOEgj6da8Cik8wRIv+T9+oWV7zZVVJL/tpicW+Qf8MLmd2eVah6yZ
KTiIaTZQhzoqv67xvjDkyY2YLNrjYAUww4icTfAaN0/UxmbUJ9rxYvKPZ7EQbKi6
ANpyAMU4wOWPd1H7lUHT4gX9riV93MR/rwKLZHKgCf9saWEaPRQahClinOqXsrSZ
1lz/KllS7Mop0FaN8JvfnNP8uNW2WQh3B7bgOKCRrnns/0ipajJqkda6wzf084yC
yebLfLL6P88DJI164AsFjCU0XypHmxzM1XBTtdv+7cyfiPIjeq/8uG4VTBg0wIuK
jUhj6gPMN4Jp75t4s1vL4XXgCuJlhvcvKEOFLa8xsTMvyAkx8+i8onZHTWC7ugBz
sLOsbHnlKlK31UVF4UNulW8oj083GspExfa3kJkMkwCV/S80ewI7zYYG9sRWBZTN
jmJhz/jYXaHmfqVwgNkfwqYBBdkT8r4oEybI5EEZiNmEOHorsrIzIafVJXg4VqfJ
LdALc8E0uhRSzbTnFk5WTraez+Z8G2uwu/69X3OhTQvs/bWWro0/oifTZdwfBRxS
RDmacPEN1Q/YVSjmP541JApBrZ4l4kVAImXJDXTcrxBoc8//9LRKzKn3mIxD/8xp
o+eBHnBMwkeCR58FQwUojXXTPZxRzSJCBBSD+F9mPe6JJmveKYVRf4EkJQSlN5O2
kqw75d2Z2xDDtGFLpseESTQIrVXQoBhQSm1ktCGiWPp4eCnsdnUxhNRV644ww4Ji
n0a8JVqcBweoQ2gwUxaVnx1ZK29fyzlj5Su13GoejG00GUJ61jg/WDApiG0Trrih
0khu1Cu49KxlNEXKg8tG/+Ze+jszVkCCh132cBgdY+EGWdznXRihP6K9jso9PtBe
9eRRAvyrYc8pEWQCq7GBg2W/3UOJnZGugg585u6BjxzdcAxp4uGr0Ljuk/t4NCfs
jl8EJiblIVHjHJbsDVjfy+H8QwYbhSRGWmtNLCHxtrJhz+0ra9FScJWoSDvsNWVj
UiAJJGeu3rEUSD3n9gdVO3Cb7E2LlKLXv49piIFzY5Esv2nVK1ys1wmCypl2IJ+Q
+ulXW7paXX51PFBzzS8oeJkepNy2nDM+Gg0C72cNQ2J/yQNoAdJW5kVTtjbF0eJY
AWpDEQyzFEticipxEQokk/vyxVLbxeKRzpfKjmdzuiTQALbHEJF+rp5V2ojahqpn
h4NMcLfiK3E0otF7J0L8bqe9yZgPrOY2EgcAcOTmcCaMTB/CUHSo5vgbgQ/sJdpz
eHous9Hhxi5VV4qE8Y9qYRKwQ/eQ9OZ9/OO3lUUrAxgjSkNLU9bz8Ihajz0pvUOb
ePdZIa0tTn0KqP7ZYZMJUPcLbrfRL2xmR9MpciB/eBYzV6amg8068pS1pDdM8ZeT
AnTShMcVwYgP7pi6udYPYws+SxJwMA6j5x2HHo/SVtpQmB5Ndxa+pctiOtDa84oH
x5hxLAE+2cUTqb0pOofMzr1W/2jkxIG/cIGs2TwJmSdHz30VtMaNLI10lVUDqoW7
7i2n8r2ujpUOP/4jWkgXo5O+IaHBpIogpR848S5At5dOTiuMcc08+EQm3Vjc6tZH
O/Yu/JcDq6WjMJlpXp4jB/26CQo1uf9xrrWg9vpFfOLXMvrn2oMHtBLxP2DXsqvm
DIa9Mx/Gd+UYKoN5hiSFtQHTljs4OemJKtjU3ZB0A19kfm01dPpbinP61KGcK9rG
MC1E6K5P/mzHgckTsElqHBBaeSqbbATor/mvdewdQ1Lm2VlOqhL3SBnQ4ZRmb1Jc
XCZUjVt3/RlUmOuImEqGt82hpDzEsOmrB1fkS0gSns6kVaEnpXWRi98eW0MqvAxK
39pKfXRjpf9S5SaDz9bOQrUnYWlc2BM+GquUu3bVzAczj2VE8CmM1NTAN1anFVK/
H2lAmIjQ8vymg88WFk/+gEEat3tMjf6aF9dVBoDozWz0cPDExZduy30Zn2Qi96WF
cBkIMSHpdsXO+FPTLuk7norxYK4n3uTiB63zM5UWLGu6hSha5HQN4bHvD2cMdf32
3zX48DV2xuOZlerHXPTrJ57o1n7iHcBlJXjGO0ycoBtbkL/X0bTaX/NyHpLEYh4R
FLFP0F7AJyZhHCcLogOfj8YvUxdSCTnmF2IT2Xwfoe+XtU6DSTYo1M4aeKlJkQ5e
a+5xN7T0R71Y8mWDb5IpdxKDQz+F9amyvQLL2abQZC2Pa/RGtxWQpchvygLBJi6G
xtJTb4uO3cHm06IICMOJvacPxH2pcGhAlbe/vOkaPGeTe74DRFWT02Y8ZlbHBE8v
zPjr2hKpnfRXNdpjEstHV7q5unD1spXXmy71Hdzv7K2xsaxSGpZikgqWjdW6+0RE
q9aKId8R9qvpbFF6uGDo90BXsdBBnSPDPN/0ILmeM3l2NlJqweNetWvXnFHzTA/c
4nCZl0zh1ybrz34Xh+1QP1OlVoTnkkgsoLTdgTf2LGTzNxmTNh2ui73MtSEF1zr7
RWfpXJpF8J3EVGjZKm1tWwGq9uuqUKfwEslVZ1cACWWml2cnY6cUL8wmSAzCVrdo
o/DLtmCqR6T6yqH/fpFjUBKOmJiDhjjZKuvldYHm3t3FAbeRpiYYa+8y+4/4/DRl
IvqgVnMNzSjMqZhq1Wog8yxTBdeDPRW8JtYVLZr0lVOq1wbrBrNMhKjitFQCpVl1
LYmWGU6MpotOKm6t0YL0s84/HDUcG8bztIS8nK79+52AITtDPozQBZsmCbgNtlr8
voPlUfJKXLezqXlxv8nq6RyIlmvTO48LPywA9GQ4u/B96GYH7vBeQ3CKalwtZJhJ
BJ8bRjk/6Qr1vGZyxoNlXWcXYkC1LYvzTPjGUUa9lse0kq2yDAcN/3rhtdTcYm2j
XMTO19NDHvxOKp2Qfn//6bbbgMeIKjjc7b8j3hFO1KWl1+q/pY9OKf9kEBbd0kZT
hKn8lA8FBWiB4cQkJOuBSBs/AOHqNUWyFZUjUom2dDpMYsks5IEz9wZDk6WrWf4k
awcZtuR4h8dXcMSBFt0HNR6sLUP/Ji4ySMs7bUZVSXQQfzDGo5VCJeLIuCJ/JYka
UW0Fr69mYGmMCtm7/x4rm0uLJG75rYUCXhm2ygzcgQaWahCB/BKVSChJBkVlHtXV
IBqxnMYqsj/D5jrZ+26wEN9Vq6tdJfIBFXQS6GTbQ/9erVA6MwW+zxL1Y4tKiTkk
jQGgkYdPmIRI1QTAhd111n3JWjGRnYiMdWjgFQhsooFfVNl2C21JQiJwcpiPdu62
Su/pv9YiFFqSGNuVMIN4uzf7P1vtskFXv5nbs63pvzEu9BuJ5UmAeZe2DlxWzFnG
Sa1C3dwajNxKF6hFibRGnbPuk1r3azZoky6f1TBYDmFkMQawZwIqb+i1491ftZ1c
ety79cz1qifSkxSGEL3lBY8IcdVxyiFj8GjzHktlBS+eFxCsIpPgIJg9HYOlIWyN
+wsZCFcbtY6dlPxzg/SPUQ2lMpGET63ItmzAtG6euNQzBt7wL1ZjsuzoPa4zHAbi
3hoTkWTDANz5RSaCnTUEtCr6kmowraPsuARDIJeuP3H3nhEhZ7pwLKWShsusmTyz
Fv4mxlyFAF2P0AdjXXPsTG4694syz7TW8RDxxSPRSXrtYnpZNWSzLr8tSWwbxgrx
FuhpkEpXezASvsMOjLc9dKNIRRwbRG7c7tTxxp0TX140jh4l7PHqMyetGADiVcpa
1BZullv4ywzeOXXJb8NTIWDvzSvFqgPxymuk+JX7TYKF/pTkWXLa5GNIWymWQ/uC
F3aRKZRoVq3eUMcpRb55V15MQpel8WwxjBjcv/ZuPIKJl/aRk+2MN+0VBV7BDxgw
Hwt9ZAhfr5Z/a0XVPCPlR4Se4ud49VhjjlDO7gBg/w9/wpcJN9xKD0zsc1URSOf9
u+nFJmDFQTP4bIob0jxDyUULNy+xpOR/Z0OZ4eioomCZtE0o5WdntwNWi8Wbhk29
ir7fMPUqLqrn8yD542rj4vobUIchHTW9R2ClZ+FzmCuD3I5aLMCl/g3x18G7aIpC
iLA7DIqPuR/moRMKKTtAZxDCAkGFW+ll8Yc/769z50ing0rDU6YYTjI6h1TWYVUQ
q6UOVztCVIblrBdsnvVKFH/eIJbS0Fjt7vbztQ6so55tGuD7BMfEIOZ7gdLLj7xP
4hLpXN5GgDguamZNkfyOnRA4LhUrvJ8U9QOY6v2A6pO5AQHmQlSyJ8LfPA9pbOhw
bW5Z16BXvpvmrvrwmplD1M/S7YNPd195bAxnIYzwX98pcPdL/qLv0NQchZJ8t/Rj
Iz2LfKsBDxc8xRyGyOFo8tZ2Gf6CYbtvCN8JGwRQDDqgDdtz++1DoMM1Pm0o6xA6
KZqkt29m9XQSfARVsJwmI5UBljX9mFEvoTaVcNj/AF5ly1P08OwpF0pn3bqWj7gz
Xk0RNv9xoocJkNsv0RG0M9GFGkstMOOZi6MqcWwRqibKZMelGAFNRqd6ZcNvgEci
iZBvq53VTqEoOTJNL8+GNss+k1faHMW1Q62ySO4gz4W3HtGuaXM4aRosSruBUa3D
so3ylK1MTPvW6+6CtGrS581PlH6/TNcQX1t1/MiahiJZ2aDYzDtXGYLke2nStOGO
rH3pdTf2uMPVz4YbZ8zgZwJkbBZioDHqDOYj7YtHofZoQ1oFr6xlFvOw2dld8ZdC
RP+FbUUOJcc2peLyoN9Uq8YtLr5BssuQdJ9YdhA+cmli3JCk+EAW46IUOv4PMQYs
S7s4jZo2mA0iUkiihEPjoAyliK2xO13D03GhUHagv2gFIE7xFt0vrGBVCRIEBFpu
nKvwcuzh4v9W2jta9tOYFydx3w8RnUN2nF7Dq2PRdJuRW8XSSQbxrGil/0mE+3Rk
Yg78PEMVO8cmGoEJRC7ImSYu8HM3MtiFb7gynqcOukRFF1l5IeLTCTRJeHwkV3mH
kZE2810PgcUlfI2SGPv7jIZ3pz2Zy0xhilmYStg2B0EDTZQoYGK8uDR+S9etm6yX
uIHFRzbnW0LGXzWztcaihYbJX6HxYBwsb4NcLo9MNQNAG64QXqIF27W+DmxowQCv
YWVbMtCul9D87vJ603D1LGIa+11EgQtB6sZ4+VUGCy0esSgWZRRSFyE5xLXVImY7
llZ7WI7ZSPMQhPlmZm8kfd8UzbYnKRobe0WkWWmyz55CUTaGyFEd/+MXmcVUu7/J
ucdGep8XELzgDgCch+j7T8gJP6g8RuBb1b9WtQPNvJ5VxsVrUOlYqD2pjG0+VFLh
UJCiRU6pD46B3MVMA5t8J318h1dVPxO+n718+lD2LMdcJM5wpvNXkGCkA5YbBkIR
kcHq0bvf0TrC+4Jd0GWqQ54A91PpIO+hV4fR9XKRZemka7urvPKC61ZhOJicWacF
wizIN7rw7Xync0upXrimWijJGUyHi7nsagVDi53QCMppMz1STFJgPIIW+Mgbmhfo
eTUNENKT9cDCPqEosAEkJxV+9NbRNfAjgyQDSojkyYqD/Gike5zurc7xIPkW/7q+
mS9yQBO787lNuBlm+iDxiHVC60txCFowy9SHsdxxToA/NO9fcK/cqBa2KFr5+Hfb
83a4u1t/XxpzNnxl+ZtP+kh7Pgly9N53237aBBISIMHOs2zrQRNWHhpkk2sfd9HA
hMM38svp7wDj8JRA2A7FuuxS/I/VOtCBEXWzJThgzaw4XiFXltlWUzWhdXbN+SKg
TQWyOIrKIpTCjklguSxP5yisig7xgOOaeJ+44sXYuX0EoqeL5SoE49nDWQxqZ9A1
AfBD99Nd+fHvV7v51U4B/0PYlDclxuFgwA1bNLzsVQGlLFxqfpMIxeshuEBPGVYN
+3zlkeReaNHF1i8HiOj9zXFu2a0n9ZonZcJ5GQr6gaCKYvk65EzTcXwdupB3Gz4E
Z+Vt0mu/344GSMgYTaGIti3NZLiyYYiOGGUuUVsCNcJqrhoo1b8rM9fQ0YLJxhVG
WVYTZE2gNplM4Pj28FRC7j70sPdnmSbhe4VktGsgnpiMcfdYaJL3jXN1VDGTkSSW
zjdYWTW5RS849xa1MBCUOBxyzkkPCpgY7oY9wbaiN91Fl+iWxQt5Bs1pLZ3+mqJl
FCPi6FW1lrefa5nqxqGMIZSFP/gv7E/BsOzIb6/6TMcmtm7BqxVKRcN0kSLPiGKC
Eh/aP/MbuFLdGrkzDfc22LK4CCjpkFEc8Py4i/PjMAz3jKmKc+8fNmcJ7QmhrPgi
HBCMRiHjmMcoMnZMjKB9hGZuabKJ9J4ZWSqBnapZDmn11weMhexXsDdGgrDTgFld
DfVyOPA++B6cYUhdYR4LLLeO4QEXjjXrJURSPfodzv6eYE+hdGRpzrCVbhlc1H7F
Uhs10/jC1oFX0adseZm4DG0MqoyN7qfKh6DSCgRqMrxZnj+DRIqZALmbpi1O38e9
u62zXjj+BhsEJu90SEL5HfS/iMyIwXHQTn8NQQ47GG5qYXC5z6SmwdbNZI6V08HH
aGnsyyK2qnhI3aloFCRLbyxKlDuhHOlBM33jXGVAGR48fSmgg+by36opKN+/Q+HI
L+HntRkc3Gx4g8+jg3yrl5QOXLyFkIF4HS5ffB0kMwfy0sq1tLZQKSnd/oXdxOm/
weim9+LOJ8c+L9CYz5Ow2PnSnyCg/WhKeWapnhkxfKPFOg8iG84OFM2GPU0DRVD/
nVsghaKxtVpnigpRw6PJzgPWtFUTkXx1KjtmllvXYyqg3heD+kNHpRDh+x/4zAOv
2wxM93bjlOBsig6JsjFLwGGG2ax4HSsprzZyJ8jiam8eFVY5lsxjCVzZviEPSlAL
S44ZmDALaaGI2K2fYI+4SnOm7nZ/YAS3jXniexPaTi4aPDHDjndajRlDHae+dFQ7
ErzPbgOoAHT+Rj8o7PbmjkQ8mZ8F0P8GxM2jRvOkebsEeCnvXXZkU8av3YnQuP2x
/KVDQsn8r5vsQs0tWpxjx3dgEM/CyZyr+KMgWzngmXWus2TEUqLH5kbpZGUhD2lq
tuofMxYdZilMszolSr3AdETNJYx4LJtybIkvjQSJQkzhReJJGSTJ/TlS4Ow5Czv+
2hkyUK3vk7IFxLAlgLp0bNN3d1gUpo53iexWYiGZtnKHU4Qt6qCHxOtzDUkQ2M27
geZ/jb5JYNRZAZP/N1+c+YuSr2kGTtKmuF5yxc8Ggepy7+jasz/RB8Q1HKNT9olo
cLAWOstko+5P5vPOo5tzBxZMsrdSwoP0068zCEiL4Oz6B81DhBcd9+FstesNg+Jo
VxVWOMTGhNqJXVZ5bIJ2BhzsfF7EqXF9Mf/dAkqAito6hX05IHgDOx1r5XxwfSor
OY7h8FP6plR9lgP0NvVKFFYkmvyhWmQpdLTD1nwJ7azTjkEgaacVFtNoP0jB8x5G
ywA8nL3nIp3qX18d6J6OWPlNjbjswvXp6hb73hnP+3iqXnBAgVPrNPjeP0suMSRN
3nG1bkc703rkMH8tvZ03gR5RNu3wr1EiOiXvsEZ2UmbVAFOZ8f5iQcErXWCnhK6h
VnxKaI/Q0qoWHtffcoLgBfOu0IPyKTrz5Je4MMUZ5L8mHMs/2oCjLQzaDu3iubBv
oFpYI1guCru9rI7lKgtRyhz9iriQ2dRY/sIIXZibrTZuOaae0f1SyOdz2+P9cjt+
YGmDtuY1jUWLxGaxCswcAb962c4Q5KLI0RBlGwIIxWFfE98jecCiRR61HujvhRjn
V9T7ff1beoKbEIUTvtLXQEa49ckESoELyYISV/8GPDgHm69x6H04hW4D879qgOax
gDB5sPkRHMDug4ZnGS7FrRgZsh/tnu/kzYzNvwK34/bGlssI0H2B1T8QD+MAO2BU
GpI/sOjG8jNfEsBAy/F2oRXAaHFh1KIbfJEpb5M39c3jenDGvA+gKqCRES+w5sW5
bK1+g/pvXfP9jlwpJZn/YhMQVLM+F0Seeq4JZQ8M9laI/9aBreCaJagGQ/5LnnJQ
dI0YhrB/XojLs3vjCgKfdvU5vrWrppaDwSRzud9MDSMb6Be1jmAv6JuWnJagmxI1
wHR+Qr+OtNON22LhhLbXr9CIZt9HPQfygvrBF0d6KZ4tM/dImxC1GK34mAhqRTuN
YoAj7GAA9nLfaRuEJG/xno+c0ueJgUkIiopc+pN5ne1KNtSgQdNdsWs84w89KEIz
275VUYUJdmq1gtfmDmBj0FgBjqy3AZVXRvEwNQn9Mn9PT3icZpaceHajBIEAVc6e
EcRq1/a/KAInia0VVjXIy3n9AYRcsVIfslG4Uu1fYj9jy4rDNc9vlwmd0+XBW/JP
5/F1Oz7Z4gv7g06Yb6mm7NK/kNEBvuQRB5+4ccHpPjXLCLdwZaZjYYB/bgcgXRac
JBioyO/S7V4P4xfKu9FsK2Ca5kEF1jggq1w4XMxl6sa2L3gdnWdC5YIA7qS92yJa
YH1fjlOFpdqJSSAlkVHjOAegRPmkcApnVW3AD5DhaVROqP+7vyhmLiErLo4zjh3N
N8fBXrGeUUAUsILpIa7OwKjraEUShwII1rVSWJgQzlUiwqq69c8l8FmLEEvAArgZ
2jXuTOrNrmnxAwPMaXTEbz2elFCpMXRkNTpS85RISMRIPps7/2WhcQi/YoW+E+GP
oLHXSxp/ttLIMeDDqrUb47gGcxGR5S0/cWUDe/AfeQ8jm6DHmXUIO1VtU6CB4F5u
surClD3kHCVdl2RxSeXxWLtNbhBTk2Gtzw1lljp/TXa7gGgjRhGbAV+0lEm8RwaY
iGob/xihhylPIx905tQsJ6AzrPDUHHuYLMHWG9/zd0dQowYgjesiZDTnOqvc0HFg
dAEKPLQNEiBa5K/m4rSI38Bu6OykFx2XaXRIwEHSh1cSTZe6SblUMxg4ySFPTY6F
AR7dZIPish/hAhvEUlCadTX0XXC/Xk7ptTSGLIOoaZrKj1y6RBSikXjfXCxjT9Di
3auctxdvIvyQnJ0A1CvncpVzhBXinsiCt7YByf6sNmJbRPhZW6BQ58AJX4mWOUI7
uVorE+byKue/9DAyxUIFbgigxWu5Ozk6wtu1UnU6gn3QRo/dZzCcIm23jnm/sg6v
YPBF6Q3aAYb6XaEnWn0MqLmzndayMzo91VGy/U7ywdv2mA5ZRs1xK5k6E5zrpmTB
naT68RolkXb0X5fX1s3DE07YrKuNG0sYayTLQF7As6PWHRa1L0On+TqJnAuj9iDd
toU95x/HkM7Nq7IwLlQoqVeS/ZET5zUkAk+fk23imPhvmQt4Jm3NoDeSjJmlqNUH
NZnDD4NkS/rBRRNGJD0VN4+6jZ0D6Jv2NxGYN8S1vGrygf3UEI8c1MttCRcuIJIC
HSegNbL/MN+IwBM4cINgp1Z5LH+IDIRlUxizVZ3vG01lh+V5wfi3stz5pNBshiVW
DvyhqYdKa7Z98RQRRPotwCsR2g84KWNShIz+gM5Cl3x1iPB4fYRNlM5lc5UYkqzY
WvAaOQ4pcNYrrzn9o+P31N0Uo/+KxrNhjuOY159rhOR3Yb3ziJh8EQNo/I4r81db
Uuvdg/Inz28RxmSw8ojlHayMAxrdOD1nPBcQVeu9CgAIxDzhL/DwzM8FgErEqunZ
NYnc32THiOFXillnTTo1O6TOJKLmZso4LJJM++qWr8PH6oXxFK3kkDpNULsIUaR/
KgtFy/WtLO7stZBqOB/utqK32Pkk3BNKfXgzPK1vlZ6nwELPDBLLVkHrzK63biek
mX7o7pHcAvwp8cFEHzvM6wvlheDn5lRACcGOUbVaOhKo48rw5Ae97aLGc8BQwxZF
sbCuUbD/3h/dA3XEkYWrdxuFNW0o5YrRZPRC1GgO3uo+8mdKjkyt0EkVtmFfxgzB
MhI4TfdLMJNN64+sq3HcvCTOAHA4ZeFXupps8WQkK1KpoFO28hICpxDZAy3AxSfA
WTm9Ywprn+fSVLp0BO7FHMSMgamqVMzSTMihvGDsi6ibcTB8nNpOYdKZXSqmluKK
VfeSexHdZIa0YI3HGLxRAGkxjZMFxWDQeqNltIrT/XCjyC/BYmR5b8pLe0aoXAll
TfwyL5wF1zx+Jyro6r/4pLf2Jofdu1DRTLsqKzauFtjIGXbvBSE3XfpOw8H+2zXA
FZCPNWufY7EUayzqswe4PzwTlAUAbJxV7goq6ysPYKy0isnGb+yIPL1Zk//YqQxT
gAmSg6CU2E6ybWf4R8oL0SWRUH5pnp6YqXwMB/Y6/123diMBCdyjHRArFp6QPDSv
eMbOQXAkkuCH7gbgbHM9uvGMdnzIH8PhS97pYnPgO3dyHicuGTKG4u/LGzdZ33JT
ggZdBQd0tY7vQJNyBclyOihXeaMiDWbAxSIMDG1dgoZ6GYKbi0Sqdp99yHzS/evb
BcFagQGGHR2R4RYyUdG0bDqfkSHbdsggVkbPsFkg998n3/so0i8IEwlwhEyPOBQS
gODZiNwa0e+IqOJz63YLvcSnjHmvej7ImocZ3LCQAYjXHiOWWJJdllAqT1P4T9uD
8sMTvUfsEuH4K3vFZhfl6BPx1bjRoqUbjgpsovlweFnAgLkezFgmnhRQpb3vtCJM
rt7fFXNB9obFnAtLcU5MYv5RiU1pXQKWqjMll9L1C2AdRRRBWp4yzxhO8l1dmgch
qAOv4Q8JjJskDjagddU3QMgl3UYA7nkzjIIGkPAZV9HkN0LK56ZMB4pmAeqLmH67
vArNpdsEZ7EbxqdilFjJCNze564YnQuYTb+4qd0mGN2z0xNq4WDaH6jSuBwpWo9K
H5T+WS7IDhEo7Q+RlLwNS6vW9SudU5TlUhR5khCtbCeGuNcsu5gUcHk/e0JkKakn
vG7Q4bzIuElGCP6HfjVYlUViqx1h75OC9c8uuensW3qevgCyuRcdbwVIhcX2Fv3G
WsLYpCXjHNyLxLr5P0IlN7rysHTfWFEwtSraVUJ3TOfvNPEKJR+8pIsuIwMTxRoo
iC+dPu6mg+tIsDxtetF5dIUXBtStSdFi13cBaptJW4qXzZ0Lr0LI2grXeiHasx4H
GOjPDgaR161mC++pmO9v1QN7KLqZkVVxQetGEZdElBZmYEBUCsNpETTvDdfOgY6Z
nUtZAdOUjWJMrN4aoqxRyOWKWY9wIqR3SaT1tvYmlLlv/ZzSb+aUrgzJQNW0kcmO
7rBNgOfjtkScsNPyxLwBF4mGYYSeVAMRMZgNJZDC5Ut24Io7nxyJ+Pm9T0viO3Se
HwhTWO8n7JCkJaYS4+n4MLQB6s44HtTIVMGFbJCLe198ntfGbC8vPO2jPeSedXIV
hAZmtyb9Mvy4cJ49RxaiM6D65NXARWmOPPQaurR6kb5G4t1ix12T6b8PkngTdf+T
JTBv8eP6p7iADLV1Gj98ZyzBuGBcKj+nDCw0X1RK7Gz+SKah8oibFFAN7IAk8K99
hEVYtCoYuIeAgke2JpjDV34UpaVGg+ONjRMB+h9xjmyuwsgk9EV23jkO1Vsdflq8
0xSGRPCyvznkHEbKH8GzuDsUb0CsxqLuaODxeB+Mg7syOZPaZdDBE+11Y1YLsWVy
a3peEkXA5Pw/Y0Nq5Z1wO+8/zT6tI9ynIrjs9sHWhw9qTyoMpgGHsQ0WX0Sf/B/F
L9+VoxhPef36gqSIZNbYVPeLvNdJbJ9MUyYh1M3rgZljSgybIKMHaMor41at61+g
QCORKSuY+dvxGacUWvBTdshwTgaSXmcLYfC3CxPGSGvg4Pxda9r6Vq9kG5YBiT79
DN6b6KLc3VER/A5YKnMy1W9OXQ2891KPMcGLfuS1b8MVJQv3ZlEdjyUw5iMI4imS
CIHIiuAex+aSPCOpeMcGZujkB2DoccfEwmS8cXrxQYKp4MbYm4vd1gdsD+7elrVV
+q7s+FdEZwn9ctPDx7rBfRyLkZ5zynaXbMxSvzKDXOTBzyBTOXNiT+gDkaqgtcky
wlzSxtJfWb8at3tXjldTSuzgepoedhmaHajlK2IBHH+sgCFfXoNxcyoEQ4eQShPs
rvEJw1wzCxKm6LSjfOB8RxIK/hEmT0kzU2PfHglkuthREwG0guemn/lPFsPddchX
2x9nxs5EftD2g7OK9GL53TLBnIIlkccC8l3jfxMUHcruF0mNF713kMJ5LaR2FDwk
nf+Q3k+istp44pw0ZjPY7enARuuo4dIvJfJGHBq4PPpS7hfXekVX1fb1svbOhUAa
yijOlk0+2LGwQ2KTtpo/22SBMAFVzOY6AFiO2T0pjgtfir5NgvnJAUmfN1Q5fsHy
4HzIiDkHzBpY0y4xNZxcafT3KhoJyNH2wt/sYohQ+VRDqCJlGq9fHh8IGuEhIrYZ
RKTyZySf86X07XrqKZJXVsvUa4MQ5GxLOlSWCX46qxlT4Sl4zusWklETdyKV8rKc
V5EbJ1BFxRiD9p2mvmJQvKmNbab3SeqvrxVZ1MUwLqmgOB9mb4kP6VP2liovThFH
vaB1jB/g3lej5x7Fxm4iH37nHbGAaP6YTBh97jUw27JyAXqZ89/x5KlQnyFhQjpQ
SwXJA9eRDGnSYpOgJB4OMcXGAylUNq5i56MBlVc/mRgFbElYvfnuairZCtb8kA3Z
GFC/JElC45XR1CtdXNNgs7+1SJmyC0aLjtuhQg1GtSgvQd64nvjpyDcT1rETIEMI
MyJID9NnGEUClx+0TQAWxryVVnV4N3yFjuJRRjbiIfw9BycPiPsWngcZ7SqEO07c
3lbf794/L9DzxCcz1sOGRhhbViL8aYVtX7prPdJPqK9apuB9AWsKNcRY3MbbC7hy
R0P7jgl8CFHGwXjvY0682ZIk4Ig/L4R31cegbHNgcxITqmwVFzyLj4wu0QXJXdB/
haA9l33LDcA90Cj7xJoyZ/tE+vXKaftWbZnvNA2HECbBRepJgD9hWekBR2zjCQVv
1nRtkVVmIDKv2lDNBWNL8NXIBPwZev7Av6frg3L0XBQ90/0fj7MKQtqw6rGAPyEE
kY20kqNMqQ6w3W+4OUnalWdLAJxd4DibNNuiqgpxdKLzonn56cX4Y9OsrOOJ95mY
GUMIgr1IjzqFtyzlr0JZLLGCSUatxWX7o9s2n408S/3Mcq55AcP+PEyC7/ITGR07
ot6be0wXjK6yMgNS9F3OmiiU/grwaCQCv/QAwrQMAg5+YfP32Ts88q7tB9P16P2w
W7Oct4VkPAj73ytFsWVm7b9BdvD2uTNa0X+gqnv+huYgw+hlCc/SSjAqqVGAzsRX
v3iGF3sNBq/AIkL/I9HEBSNUunL8ZeS19R8WrsU1IyrwuTTr6cPPr5At8LSuyZL+
EYTn0EnAT5F9tKd0WWPniHqPZMzzYjZXEidWMiB/3ATg/HGI5hmjadzCCSDNk6Y1
tCvE7XV0sPRMJrYHUALa7AWGkgG9UO/IzpFfazHhsTtCQKLTyS0Gw47Z0tMSyhWO
s9vaksSQ0FgT5hCiF4fh6c+7QvTeEa+Af/zby71tFH0B80RuOJlx2Z53ycHPtiKK
NvX0ri0Lu8+0WmCG90MYLfqxQZvxUrNqCWjz+2/IlcldqwOLnenIrqPD2iCJBm0k
GUSs1bhV5nuzTtkShwd4ylyYL+lDmIvhlgLmLAa14nv5Ai55KqLzpKCWvVdMfXZr
fNucNvupu9qdlrxEb9DNBpKlkTHeW0nL6oPBj+7HSqlBrrpvnV0Qk/+/XQVKyUB5
616WqXnRxdSN4AfQ3yPsn/9i2sGv8EoZT5dxzsyW2X1z1R4nQAe7w14hcAYsQXd9
omw/gr7swu5CFi6AGesTob5CJmH2kVH2ohNMOcJFnRf3f+1gNGH/hTaKtY5+N0Dt
Zha54sc55HOUeVMdqdHmhIaJik8DhSzi61CKN+F+zM5cIR7IKOIS3IWRVCZrlKpF
F1JL9N49sR1Sns65w3+bxnxGKKAIQ8Etuq0zWjpBv+t8KEonQnh7uBhIB1A3Aq+1
W/L7EFvZ7dW1gELRks3o+vhh+KFUJVg6oZr0IUcvAmH3dL3GkL+y8vy+7vkpDdqe
c8JZnqSxwCaRABeuBZDSnwZwFsCvthAj6ACLgAHCYykytAdl382mhLZNtEpYsJRx
IzMHaZCNjYIxRljkm63gUgZN8ANasQUApwHsSfLYn4UeWI1T1eyOOVtSL1uGYjln
gLs0q4ChGpCMJ/Fckthc7MwNcZQ4YZ1Mk+RVzu4L3B4rEDqAWPihBRqkUcTgQDs7
ntX57vcOrXS0t25ypopaIV+1ckF9orGqDv6ViIaNrvjGUk3CwCPAlbKxRpSS62q0
2fLdRv4cNXXElP54JAc+/6VO9B5gKBlo0jXzjnBzUDQKkSzUrNMwxmk3ns3gBWRh
3BB1Qyq23ckp2rJNvdJLgY7BIbSkNn6JGJd4gVZ2nP/NqpG6UyqjssgKhKdhubd7
EGV8jXegT6KsBMBxTBQxPolMWRMMlhp6nBkbw2b5woKma+U0BISmlD4V+rNiEF1R
yaFyowLXhSnrOkpUOIptDPuJpUgILTlmgJT0ciBoXKgUzswiGRSSpQEMFAZ+wuzs
mmz7yTDhSa3ceK2k7G3ADTjtvPwRRR1tovLintSDM1sGMgWIVP8ELv2GsXTq2Tg7
BU45k6meqCSV3DdjANfqYwYLJhIUP9l7xK+39RhSKjqb7xRQMdwXo/xD64bVGX/F
WE5fpkDbRdWaXlDtfUzls5i/eLXb60bNRHvOQgtVD2eArXmc0RL0AMf3AtY0v+Di
LCm1z6b5p4xBydJwojB60q+/HBZPiN38BeA9ryAtkju86RB2KkTP3AimSmZffAvL
kxDxaRg1eaZ28vZkAH0P7jBP4f9BEKNlDAu3qp+LlMronGapzcI78PLMZNzn+t2V
N/WTe9saCLQA2m0uUq4k57MGeBH7+1SGpobit4BoNXwHd94ArbbrTJIVaTjVJwEr
VXoGt3KeyI6eZoIkCu9FOBq8YexwWYPesebnwb9THe8yy3srwEd7FhL/AiRTZJ1b
+amDNHHsWrVjuBFEVJ+bYHR04+HKz6Qod+v5FgPvVOxq6B+cid4D1UUwVckGGlNn
NivXyRY6YLJH6L0gRfqdDa2Uj5GY7gpmJDDVSS2SfUawHLJfjqakUuWWX0GfmiWJ
8Sr9EgQLNUgKazP6zZk/nOaxsvFh1KfhUD8oR8TDr5/3k9jVao3jTsJ/hbAWpudS
7u0Y5ri1bR8gRkm41udlJoqfLvO4MhB6sSmpzdJkzIjczWmdVe+k4qjvGhwAnjLB
GDqbRKX8imtbDFx58npX7nVhrRn8InPd5fbrKo1xnVbUJtZLIh5TfZiq72+5otAT
NJtMCeDeyvE8iXZn1hw75tSh8JNzPnr//Eu0ZwfCpjqlietk1pqPmOfOriQuJ1UV
pC/iNFqhd++5ZyE8Ie+PxeVyRxf9JMZmehIOk69BVe2Fj56yIKaXAHMAHam2HHdd
sz15/CdC+S+6QLwj9/01nKgMgUMWk8no+Pc9kZlW8Dw1hg0LYtWQ20KzWvrzdvw+
WJiXBvyWQHoIsBVuDXJeBzVLfw+n55UqsqyXZ8Akli8L4Xiw/Hk9wvyqHsJ/Wg0h
WeGA3Xnx5Rtc0YWlfODx6kL8u1dUR/Be+19MemB3QmRdayljTUQskBKbamDGztr+
WzBeT/17FFFFocKNjiUZyc3FEC6abn/hMxMeiol+/1y/AdMS96XaSqYEvhyIPIr1
0lsmQi8yE5YIVEc5Wz88i1jbIzOPfaJlhQPxAQfQcEssKcdKdyDtQGovKH7PMzow
I27jPnV+erajRI9KeD0h93LkLpiOZy7xqC+ya1sDZuy6B8x9fcasr7KepP2i8nmL
Ac6IBM8OIfzPbskZSLX08sEe8X8F+IQ+ofvHEeQYCF4aXniRhWgdpXPORBio6DiL
OEE1PfITAHgMtyxLaVF1Nmtjnfxx9HM0ZUukMAeOYOP3AtlsEOXMYQxw1c8dubvg
QTo+x7HA5XB4OE4pJrB0X59rQdMMVTHl7kOsakTHmoz9Oo7JiyjkvW3Kf2/FD4DS
Kvtt8SDbkP+GxpKlyL6bgfjWPFgGE8E4h2U/Cv2E0ewI3nxqF6yMfFIG8WSk6+4L
0wP+P4oGzzb8tlXJBxD2BJxeuV9JuY/XApxNd26k6fcm0J9wHNXwkIkEKvvAsgYG
f0VIr4eyZ8IGroTQfFpt7r5W7FUY8akMzg2HYBcQ6+XhV/aYD0nHFz+vl9Si0Lw9
th5BTzZQV7qy6X7yyuQHdIi/P0aqPzN5ZrL5VOfSkQQg+JU6ffQGnlLAWnerCN39
Ja3TBG4qmP85N3h4SlXiU4Hf9Tz02iPFmBWqPPCnlNJHQ4YxSPB/7YjGZZVk2pOS
yCDmX8gd0Gk1ZZ1goA8bH/CdvVjhqvXgrzUK0FVajYC9eskT9DQPa+urjcpfIlO0
TV4Mp16QNCCZSCmm+h3kNk3OlvGdYAmdEwLsfmpVXjxrT/puygyI2HuFm0Hou91e
Z+x8HMz8tfuyDzNj4/8N6UchDHzTN26j+xTptMGuFlEbHLZOAnDCazUisrvuDwhT
dovZr4J7mPULo8702+S7D8TXaXJ8QVpYvvuG54+E0Mm67HnYLEZP/30A2iSiWksw
kkvgE1QtW6nTHPAmeBnstpYpWcpmWjypmbxzCF9hGj07S9j5+/yv9Fa8q8SSJbLO
XW+XQUQpCLPoDmd3TsFL3PFeysDFSoamPDVd0S0AJrpdk38eOCGUhDiPIa67YMxG
L/kXgfd1z2y9yqWCXIp1NwwgU+RrWkPslsB8XBdTtQV3P2VFdUqN2ZYuYQstIan9
27ae9D4tti+I3RghDyqMMy6YhjhvkvTPBNBgnmMKb1Iu4reWzpXBYn8O3A5mLBLa
dUCwqJQgCWd97Hg23GmfNISAyu/BfaZWuPzUMq9X5k1eBwzyuTC3gusVH3tnXAXg
RPQGQNvFgY72kQT4O28LAFQka9WfJbDIGv8XQwXi1BuujFwkrzoCVUzoIm/oT9cs
Ua615z0WMNF8ygJpRj+tXYj3/BGfOQoQC+ZdGeV+zh83d0IV0Lq2WhVBtUjEdYwo
baBShq7NXp3SQiRXliR1OgjSZS0M2/S2LxLeR41sBCgvaWXUeN+7IDpxNc+fu7U+
VRj+DO7FUEZKM7wTlBDlOhNte/p9FG4/1RkkqECu8txkkY0NyeF9nfLu/SfTZong
Fpx3mKS1RVA0R/ElONCovamwJyw01ZKAR3VHO0j2Qn7qqwRp5+uV3OqmTGD/Qpnx
mXNrg0l+ZyjnQxIeGCkmGjgjuL3NOVyTa7ntxljlFyxBjMjWRPq/042nS6GpwQ86
+XcgDJ7eH5GekDXG3Q8qvkHiNqKjLrZ0DobOkAdPsI74J9QZCTh7FtqwgmUzE7cX
sGfr1/rn+Rmmp6xhZdo4nZSi+nd7XnU+cieQQE595Ujfo5MPYRfpkC5EwziECMA8
7yPfU1MjPl9dn6JgQpIn3SamjAt2jnSIlTkWfMalhbGnDdrS1DuF7v0GsPfTkZhB
3ZpOqscHDEfP3w1CgLdLJZs76C4EQkNaM9ahbOzKe0+liRN0SmoBtREthixkWCtE
bz0bZCwBO8QZqsGGqS2voOt3pi8kdacSYAkgjkCAHDgGf5I5U31SZeWGgBLLYNT9
8iQFUoSAzwuJTKu0JiNveUo+/YOhENZWawNumngqXliev2FH7QQbnRMi6ENHvaAy
Y2BIiugEbzn2xpo8mVZhyS4kEqNASDuMlp7gyBtcuEjfIZVniyb8ykhcVsTWRp+K
Gt78OUIFp5z6U/Xgi4JJAHq3qmrhvH/FT2Z+ST4w3UnINdadOLo8HAleyDZRAkSO
Ll1XESIu/45KD3eTRufBcquu2g/zWePnUAqVbR6yUIgkx7J+DxB5EX2dgLA0RxKc
1+cxT0vzDaU8D2so5h5VfDF4JvCexYXFndAQFizKxecoE/BKOo+VpbpKV79ELeUN
Yl9FOhoNOQL+mD5Th23nfJbB8qch+Tp+29x2gc15zVjnWkLudt5ywf+rkdfRnl1T
8rKzDrko+IobjOuffa3GHCkJbsWs4KHev0vpA+cMH7tQSLn8v9qe5JlIcQ4Bi8zt
W1P8RZrPAzZEZbTw5CljuKePPK402imSIMw80cgyTYdqtg7SnQDVuB2cfbgeyXER
3VxBkltQBmK/IeVvwZwZ81Z/e8sNUesNXuBtM9lFVve+2Odypr5SFhu439k5sqIc
9GrjGJ3ILCNsusX4ihkeVmh3zpWcyD4XkZWnBWe35czRqR95tn42zutVJVVrvBk4
kuiHXiFP/Llt3m6qNNM95GW1qIkg35OmwrCDv8D9W6hHrsBXaEnlnGs0QQFOnkHF
kowyBwuEDcSTeC8ycsWy50yaXdQ0e7ZxkMfN6LDZgzEYcfOcSV2plTfsWv6MJdpB
Lp3UOybDAOX1dzPUFQlmEgOKZa4QjuCaUOsEygYJFTiuDmq3VjPPDzHZnLuE09KH
TejEgtjDTIWa7inNx8BB4tizG+uDFyWmXSCHRXgeYEjyoUtTk+R7934LW8wN1AWA
I5pnfHQkek0Cx7/0Edb+MJ5FWmeyTxU+x2M05EK7mSS13BmGyF9FdIPkggBL5t3f
WAOXKL1thHL+OIwLFIm9RTUqQGn+rYe1tPkK85Xi64SRhfST517EVAOQQigWHl10
H8ZskPY2n8qYOgCiZ2BESAgQ+KZl70/9UYfl/pQTIoRIjK7bT6ZRI1k/DIoa591l
re7vbJhdNb72Yb/1RQZuKT8qHrgVGgfSbFQscZPaxr8hm9N84No2OrM6bIPl/pVE
iz5mTNFxrJKLjkeVpWerc4zR8RljtOLkZwAuhAb6wCv5smMKl8gIGIQpOvE+rKRH
Mtdfp1QQEJYdnBsklvSs3VYJz5q1ufL5cm6sNXbsVnBOE1fVJbuY/q5rLdzOIdL0
ZojxvKktZ2LEiLTsnPkMSCXCMVqqoQNpUqgGsTO1iDZJ6NAgSJ0+G/BJ9HzEG2yk
fjnbLkG9tRgmygSYmFVh94VuCcrUi0VTf5Ar3aFqRYorUk3OTgMWFdwYv8wcGcab
oJHTNbwJxXXttWr2kxknI3Bu/R+FbA7+yas5v1syGlmCXPDwcG3f7/8rRMPLA8rP
c3iQql4xGkZF3x2dtb/yMIg5yKF+JfA9IMM/bWEUUeFvE3zl1BzJOH/1GYyg3gOE
O9BhoFRJ5yh2sRXsmeW1cCsDAa+r/X2oCvS+iZhmi8M0RAsbp8c0jsiarJ/qSqSj
vmhv34qnbR9GyXMlmlfZhk4NGPM6BUiSHzynVVrXuUlsbd8Ss6TguqFP7PjzP6KV
6KkhDiANQ5Vzqao/vh/7MuBIjquMrpDz1uWwT7B2Vb/I2//Y9K9bqLZAlfzweoBG
TR3MRh3/xPSYOnzxm3aonAVPLw3KFIhJHSgGIrGArsCweK8CvB/cLneAMtp1dzeZ
Ghd8GBUjKEIBwjCZDB+VUoVD+AYXKlVqxWGVMxWK78Mb7vBy7V5QM4wqdb7s+4a1
pyxpBQJRxWcwgyi7jzkIcSA12/bHIDNFBMUOi2dqRY/r2HhubdVfSFUe3yb1utt7
Aw1cils3xXn1F+sOWPypdHQ/UAUO0d1LcdeC2H/YFTKK3QrYNO8mqzqQ2c77JudY
5rXOB05w4B3P5Uh/QfT4+tY0sJFamZ5CG09SmCWGnoJTHP2OMtOeRmG0CRzduVmR
aFI/e1GkMTuHF69Gpfy88V+xeQZffjNTSR1yxK2+WvpZGCKFpvbdIkgj/NbWthnX
mgK+W8qWQCIcKpGi0I+FKaDLbTCIFSmeffFpYWzZ/TFUuqBmjOUojlKPv5+eFPd1
2kANyXepNIgC7PSPy4HlZdJnxtDloaSv8BZheu2/XV6KD9v6gx95RNoDwiIK0DMo
lKzBaom5gozpwJKszdHrLmJWF5bcqxeOzyU6TBF5rZu6fcPpqjHyr/JYg4a7QB+A
TJVoS9fE6Gifi+H7M7DYjNtXZWtcr+LQl028ub1vRtHqx6MZp6+koozzBmU0gerP
OKUlaWqsvsNhkxA+fIqBJV/FPtL9FffY0q2zzhtr6IJ04ONMMkAeqZZ9TA5/V7Ds
cWo/J+6VxkxvwCHHHvKRgpO/9oYFovUXFNDO1fIO9EP7L4/WNC7g3BXlPG8DFTU4
oihT1b/0FUBWuZesPe/hXdOumutOWYnyJuUsO66E6QwLkf8BxGjpKc3zVO03fjgn
FKjxdYy6ZGoa5IxZ9TdGg68oc+dQHq42b77svlb1WW8u6vFwDUR3xJGrc1xKIfG1
rlVLT7q6bRrf0Kso1m+D12jA7mb8e98QEJo4L0kNZCy35uxIfQrFGPLIY6PASpvP
yYsr5lbyGb2ry0nFYQXzf5IOeN8Ifx9sGC+d5ACGxJ9cwCV3FoX+4S/Sum7bQvbw
iZGCswSk2vR260YxPY05DtnMvc4+6yOFWPsaMGOQmpF7drJZc2DDPLu+w8O0XaHN
uLUFJLdvn2hF8CDJ6eYJtxgP0cwI1ZfEUDJifS3qmogJWRoyIWVu0kUPBvHobWeO
+RQWaTcIUnLOuQ9VypMiIzehWT3Tdbb7cKtWQJsbSmYrozbYq003ThWbKFkFgDcj
739GnJn1mrUdVy/gXNhguAoTWFd6KDaiA3nBeEr4kgYmWY8miDiyGy/sqRCed2Gb
zO/vaYPKyUkkyK0ss8oK44wV4/D9oiSIdB97vtyHRWMowcUfHPtAR3npHG42xoUz
Z8iJkC+0tDkjmHXxaOykTANTgRbY0QWdOp2eoUtmK0Hjb0sNqbxh8Lq2Ha6bssjU
nTyoRUm/pEc76wo9MZhgpvMlTrYnNoYluHlbw4RdEzCSzNfzL3FdTotBxls4KaHk
b4DtuS9nezWUKc7Vp9phvSPpu9kLReCBQYujq/aIdqUfj6AD4kxkyXc8IZNqk3g+
6LzjKHHqSQZVIaBQJpsaQed7K7BqpaZXfAsr3OsI//mxfym8b8Qv8s2SkNblpJ8j
IqgFN56K1OstCUxyPeQN98JjzyP9seif+/yDRvqL936VGAZiLqvN7fKsIHHSCoul
X6rC0ArZTXeod0vuYhgXau4PwXWCwXwIgqSsqoSEZ89NZ8aYVUznaTbZgGryx9RB
md2VtLthzowzg9CxfNUAdzZUDCg7RqkDodSDWdFVxENOnqgsS5DDL7SslDLnx6mW
xyO0/Yg3FfyPQC1mKRot97W6DichOT5BpxHLhgBmwJRpAt2IUGQdjR0wcG99yuGe
SRjzaHmuohWTKBzcKVRDwcLPotXtt9zhuKKm+CGez3h3gfOROT78u4Z9NQi/VJGZ
GgDWxpPDqAEQFY6unj/44kgKm8ZTH14UpyEgXKtfk7dCPYeTaUeY8GKBDZNrfi6A
rJdxVteub5NIf3Z+lqiZ4yICqPt5YpAlA0MPDYDj5MqWf5TCD+DhQiMPvQCIjhZ1
pqsBp94nzoOKuYxI7ncGg1zLjbt+zkb7dMUxKda/vmv/oOdPoNh/I3GU6Z2ZCEc8
f8mQwqqJ3vhn/PgaQxJ5oD6bbahHlZ3yGRNOSkCmsu9jHliwMQMhOVDlrAEPjfk2
PCsVc6OJd/+lRVN7cn2yhLv+78h9MT2Dz5IZsh86aFskVCUpuwS3izAbzuPYz3D0
LO29oisW343VZf5MGnAfPWOT3ZtlxaAHP+ygtCBx32dCxQgKx2x6/ehbQwtY9MIn
xLZoMPEcdOZwS0gvrja/Qio8pOJdY9dVkqpjJ1wnrg8dTKs7W+JOmucxloIB78Rc
pKHJHO0tWgIITg5L2rTLzmGWIRYvt3xs2EIX7n/Nq4Prvy81XriWZGqRgWqUf3hb
dVlNPmpfFgw8Dq5gEFqprGAZwjBatjz4f5WIZh418CZNfS+FJ8LEhjV4hyrozXVP
mr01INP/4LJVKh7tW5hnktRSYPCzuJSucCaR2UAC9F/J1t7FemlfU3JkzW227gfW
Ttnh2Wq7zslLK8e+YgFyUQj1JvU9+NmBW5xKMb6RPB6beJTtTeWQPUflStQSH0oY
6WXmJcgOnRLWDordeGS1Cv5zKBj1ZaRl2ciyTgZJtcteZPYfVZRg/0sxhcTvu21o
lAehKaHGVgNGDf+iYFaz8ZrIV0BbbWJwt+BcdFdo7HAYfTC6XKG9+qm+XHxYAgCa
CEyUa3+Udd63SGCrqWma6/coln/TrvJNywK32W4Gxrq3ZIIYWZ8ZHStOCf3PsaAE
FxN4qTwUKmtKLHTvJXhRi6SylbnSSIw8hocDgQqbSP3hUyH/LUKRlB/15ZGw+3N3
v+ClwfSNPYthx/qIMDBhCVitjXGFGebivLGRRz0V58rbOjnlJ1+Ioz2AcE6ljTvk
IEpVWoQiO2j6LeyDN5zZwRXDiCdDRzycA8uUlzT/5GtirTOy6F41T0Oe+V6ANyNa
V8anbF2xttuarbT6tQrp8mKfmN6UqF6yq1qtqqp4O2Kr1wV4ZqNP8zH4/m6BCKOk
wIUR/6rvk/kaRMWQkV5rGxAi2gyEd5E8qSm9UaxpVUfiyUGSMpcH15I28a7qwD6T
chkBXhWAZENiEkSKlNizL6LzkbMm7bl4rikjgBwrE0ZM+M39mCuxtBwj9JTCSI5p
QezF4hvMBOpzb9Ja3AngKYUh0dOwxat5UJzivkFM1WK8gQm9H2Qt80yghd3XC8Hr
mMQI+QcSFcoE+WdOw6Pk31j08z/KYyNVhQC4cS85FcI66mUlyXREOZ782wpcjo6h
uWuBNj9u65knitUzyq6VJXVz0muc/kpW5DpMdqC5W+cNKqXKa9EZ/MEIUeTzY10/
UFZEKXwkCy8+j2A1NfbIOSuFbVzecWzBremJvLe//UpX0CJ7JnoZl5cpIVuOwvyo
mnR3VFyfncgmY5wltCrstJbnDLcXpz2Bq/PjPwDb+xnj9+uFeqUpWmIARl3MUd7u
5rCb4GF6/0XY677BE0Jl4pzh5Fdt7n/koBhWoZ4YMoQoAsVYuBVW/LHCpyq5SHhv
kpIRp6Jkt2bQnILwEchYKgjblf0GJSDvA7ne/BJztbf2V5MeLQvSjrXZuDwbuN6k
FzJwaWihbW3ZfGfhPiA9qFFsyysAAecMufnk5VGNxC5O6s7csQQBm35f4dk9gBHH
h8GcOjjA24t2aP0x7Mo39RuM81GzTHcWmCYwUFdakyVH2xRUg5eg2koVn47Z+qu2
WhZ58gSAwHqOZn6T3ndXReTywYQhW2A4NDjhbwi8IjhpdEo6dcmgHf4AbJt1ec+E
2Y8vzSShkiB6hQkkze5iMElIg9thUgsOgqr8K2CLnU4wondvUKSiGCyFQEbKmhck
Tmiz4Ie7oi4nNigJAe0qmxKjjPaABVsJEgz4lQaB44daZvCS0qeOUfq2drr26iEl
oYfBGvq3YTEa4kbekRzSxrpnGTQWNG9ZXQuQ/Xu5PAQ89ei7ZzLzBp5ZY5DTBFWc
01Ccsk+N/xMe6MK+DgGe8X4M2jRI7Nj88OWRPT149ApAY8jp/r11qyUGFWJD3uxf
IqJbo3IYRKtgKYcpblJAzdbT59Msb3MWB/oELGp6wKZ/yOiEL+3CG8SYlJY77G4O
rbAkNHs7YfTniJrkrQRTTwd8vf7bIflONodjfUebEGrqXHy2XaqcI5rPgKgcxsHU
af82DQAQkBN30rW/jc1BQHsiJD9GFpLQfuElVRwtHi+es5oLJ1gCF5Sr0PLbLEHP
s2cOlej+OU0HAfSM98S9fD9wgB3UeECmuzNgUTG96gI1T0h8CI0+MkFZZ0t1XU2U
dXQFkdgQK+qDYdq82NR1yD33YF0o2S3IYLYM5Y+Jgw+E1AbX4bbn4O/zaz+3vYx1
KdtFryY1aKHGLzCnjvBjKXHTFHj/Vo767Ir45nvkFZSQMAnfLoEBL9q6zQr2YTzF
cEyjaNgkNX3ezY4AggSelBZ949iTrmrzxYX42X3nfVnMeuBmIe5V1wvyawZv3ilG
GnASRS+K3mtzkN+rIZNHwBlwleP3PV4ICB3XIr0kVxUquDHVjqoJJwFs4PgxJ1y0
/Q502ebgeRmo88cemdlEO+cWDqcmZI8L/zT2d8mMj8Uojxkvgt6N3sGDKms9XAWF
Getu4ptsPuLjAEZPMCEsKY37UktOKpu406c0l59xrliOoNAJmowR4EriUgvlKwZU
RHRsk2PGLwDClEjiujgH2KdCkGZ315DtNs6fUXj8iZNJGDaxbLsIfqoqjY/c+Esm
U3v7QD28SFjTwNMTEZH96wSFgP/U4HSuF0lFquU1NWXDpAhB25sdPe/bth/QuSeU
9EcVJ1uTt9HGO5DK2rwN+VqpxL0CpBb2hWJcZhAEd3RjwlGU72Wkl7u9qwg2a2yW
eD8o1RMJ+AnYwjqsKBBzC9cfKI/7ZRpKfSDujbR3Nx8FILW9IZYK+UzfP/rFs4Df
YPlJW0R7E6+F98tmRVUj2dBqNSs62QGo1muYyy2JttVtSDsUnNoXf2tq8mNmq7HH
zkWUxHXV9JWc9YmHy/ra90YmwsFqT7HjbHQNJXSGPa4n9ojnBbv3nDh3HvXe0o24
aLg9oEzIpnI/uK6Ikwuq3UBWR2N9s0qfc/r1LomHkB1dNxiCIHtD/aUUrMiH7Lo1
K1l+TmKrLe9MUXqHrIn7Q0K7lCdolKm2GfvF0IfVjSKv0WSCc+dT1UqDCg5pyNqa
dHErYxoHxKyshMcTqwKKyrrfF/wd1iZOyp02WnzyrDGsSIr7vTAekfm92hZDX8av
ywQtAX0Hdz2o8OXwnIXjBcGuDBVSRXfo4N6Uix2xunbGIyW+G6J6F7Gc9Z5AJL96
hlhbNNkJwKK1v8uXpdXRB+OwMazxX1nCAA4cDdMo5gntuXOd2qzZEzMavYclQVOt
dXhSt0ph9Po9XOtnB03uaCx3XklT1wKIRL05A/otavweMJPwF42k5WWG+EJR40T+
pw2weML/2CUfbdGEKPHWF/51c6BEQ76DlcQ7QcgSlt9egtR2RkECWXE+Ufch+QvJ
ABEgU8A/EtHP4EuSOMFBCR0mDk8gmFV/szcDfPz5rtsMtChiI8abbnCkQ7obbBoE
ye4t3qxY9l9iUYaTjt5ERY6sueCA71WZj6dEmeuvLUunZJllHtIy/AnTtVUnZ0De
XF7PWKLIwR8i7gZT6qWaLENHE6iqfRMYa2kVraGSxBou7Ebw4ITOwBJYz4J1THze
dMMA+mCgYvwzPY0lwzhBKlc5eSAZ7dfM6HkVtvfAg139ehkByENJ77+rNMBQH4u3
y6clH4BM3K29mKPknbZ7Q9bOpSZT5xZ6aMAKuQgofcKvwSBemERmZgeJXTXCEsJA
5IJQdZJ+wPlnNP1g2LA4AXhKW3ieJxscjtPtRnJ4FsjpxoZV0EpWnSMPjsV2RMHR
8Q5faFToborWIjhVT4q+SLZBfKabmn0TMlkj4LldJJ+KbLyIKM/8w2DkhsqxYCgU
lea78Uns3yRoVKdXcvwVSdOjxj3GqNlfCui0mzPjk7bPIRMFkpPs4NB2rnWUvId+
SrcZCsSHtqR/UFuVSn62gBvjByCaz/85znAUXyC4vLsGX4ZutyviorAF2mJRBSjb
qwtxZfJsu4s27CWywiQguXH2N1N+4rJheRO4xQBJ//iWDQYUYKITomINFPXNXD++
6rNys4buPVdKBI+f6r3Ui4nXkQMaBLgzSAzPjqS6VdsTT4kZywHI0P5jGdAYdPpx
NQuvfnjPtEtudwNadnZS+c6Xu3NSyaCeGUKwpTabUQcEGQzPvbIXzDRCZKEmMKRL
WJtXNALcMHh/7MvyGdPnvxUQtvkZq3nvOu/Uytsv+QRQUPdLDuaHnd86E/KI5h0B
0ESL03kW2/rzrt2H1wmw76XxhQBLMc8fYI3hXFY4XfUnRuS7vSEWxQioz2RUT2XQ
J07P+NWQ7R+9fkSw7oP6oV+4gk53tGI4qrxtNqTRdaEmP8iiJUXCwHT/2F9NGiyB
B03cNQGvB7eCKsj7SicK7psaqqT4e47dpQCXkE4LvIQ1DUKaDYrLyBLdE9MiTiGW
ogRhE5G8jSf+ZJ0FhKr0VS2gEUkv5x8ll3O6B1rynoM/ApDSo/9RQ+iqVSiChVCn
BS4XB5xuAy7wyxu9WFFklcx39Iqu1yrzr5rx9w/eT18jmPYmVlM4b7vPZ36qQZGb
Xp14Le/y5fPBvs9mueTb+VGxpMf61UgF3mX0ATDErN7+TjqwlwE7Qqm3AU1vzEIc
esEvUoM4XuCl3asXb0ptc439qgfaPzERZKG2iGgOYUYvjaEh5pV66jk6h8SDnoSd
ltqRmVlM9CZecaXy9p/Y6/pNxI5qEAG0i8Gpe8nLC1aPr34290RxKAVJsB/ON7xZ
8bq5UYVUogQ6vpPrQQhgSgFnYmRaUkqJoR4FvhG4ejpJjx4ElHe1czgGOoYVow+u
F4x4i5Z6gnUY/F6XvOCsbfnZckARFDHYvJdBNvtMs9c/SE0qkflWKIZwYZi9xzjq
1tJLaAp5pej0a/DbnDyHjyBcKEKfnhtG/tQt7w6YJtLjyDr2rhbNt1UV2eRjg8aI
oeSOMYtvkciZGschmRkD+ZB7YAylZs5rWntRR9d7EcKL8ydRQmd4RgjnYAQ8xXs1
qpMtEiisNjsZ/zRXxdQ+ZAplQyI5Rm2OIJwnbdA/9Y6p7fnHsOWk3jhHKTVCYZ/Y
yuLbT9t/vf3kgsf6tq54oIvKAHkK/bfmTonQvMNh5g2axQMAxHhkzKpPr2g5BoXY
ME7XUBrz2sbFbdQpGCeMvaPUmwRxollOlzRtz11UlZk2h/PhqCmk2zoYlFN6uXcy
5KQC2ctNAMS8/kis6ZkhfxezHJQUysYpLV1yeU72OL3O6InA/KrGy+16eQFtaB1g
VoWt1aEyr2/YYn3CAlFFXQOsaKK1OMY7e7ePQY1Zyd3PaDNm8ruiALpLtW9ZgQeY
QPlqhorZcmq4mjvrfHOPy1YY5/aanxSeGJ/0dyLXj/HIKgy6pEUNv9faqLx9SALy
C3MJc0s3QWuHf8S/c6rvouoSySfkdlmZqm5toS/HngXQmrYCegY9+ynmwpjNNQhT
EAPbOvMWQjSHiECyFMoT4Yy66MUF6xKZyRbYz5NGEdQB2TSxWUDOSlDMmYGJDhEu
Pm8qmI0UkDjQAs91pZPsVtsARC/8YZ/qdByuZjhdBDhGSIpEK3bH9UujBACl2Tok
2Ex/7xNo8f8hrmQt65ToREURACFFqk9zfHvJJH8qytjoFQQPsLrN/kmuACTyy3pt
8I3wEncSOnjHFm8hWXoZiOrDeESgjCh++ga6ldOgbSApLXWRJOL33IGhRN3X2XYg
XElw8R3kijrDo0u9xguCFaNWEelAVCyQ+Nqb5zn8KQKZ5eQZONeYF9rnfPMTfLTj
S0VAu+aFAoIRhj+yw2IVk/0Pj7NUmgBJllRCZtsykpsqLlEjIa9EKWKpZkjvqN63
27VzY7vGgseIo8fcbJULOvS94l1BAMi6EmyTxboC5m0MHZsKadUhVHBvhYfGDSB5
bvU6Rw0DllrxPL/Il6ESMt6Y9zIOD0T1OKtj2QwFWbdKsgBgnkso+fb+wSoThozS
AV6+pNIdTX6mjERHVRihmTJskYv7akh5+o9XIFS6SrCqVgWIJ2ItqMWBLTPU60FP
rQxStUAt6LV1mTAzL7N3+4VyYdj8am7OgsjpOPwQbArnQsRt6VJd3T8giHcKD/5H
Ex46mjWBoeV07Yv3DYZeLdx3wjP+UcCFzl9eIFbOE7k7o0Rw8KtgWNfzR0uiFLc+
foZ8AwsZB3DVElcQOatYA0HxSYe7IPtj7399JI/v2xv8m/KXta2WjXMdrzd75Wef
z0CSGAYxwV8gScRe3FSR7bT7Q8S4044iwVfF5xLR5T9YjmSj1cOQTtSL9XJBqRyp
CLuF5yORehtD/qw8dv83eLnVkYSM9UAUvQYOC1ukmVDenLe17IgXrGRr4VPlQPpl
I71G8OHrTm3BKU3cpNDFhY4R+4oRHj+zrNxRXF8mDS1LGk5MSLell/GDqh1tN/tJ
xCut4lGdDKh3EEXXteUdwa7ND89tQJytp7m/aP12e3qkyD6aPi9ANCILwEX52lQh
60nta267Ob1WnVSA2t49EN/VuNLOPZ8dGJFIhj5xn8PzNnbM+2uKaohHbOow17mt
nU2kqNuPOj1WbF666gxM6pFAJnn32qbnpQZt5lgCfsPaQY3SSfezbEAcI+8fXKWu
xG99aiMQuy8SrwO+sqV5MSCrrBIZcT5jFeAndr8TqHADvSG+ulGqexdO6HvqeyCi
9gV3LIuoLXzKQcOnayEV6Tglsr8+Io3pamyd6r85f2Mpiw5Pn17wBCiWOI7uyYP8
aoV6R/QdHICmQfnwAZtVnCQiKTOqb5mTMrdcW/4OzOpkxweYZDdyZzw2LQbdjXdL
4m9Dv8srcd5Vil95s6zAMvPGDOlYbWW3WILZlaEvXfOf/u62hC725NM8NA8nU7jm
nH36/pt8Yho9BsY97tqgEPYRPu8D8AlbvbIQnQPyzCA83qU9+y/0PmfJDYULt8kZ
tq+c0sA4n7PX24lQHcirCmY3iJNI5ze4HuJ7DCr4WrBsq0OHlNgX6IwMoHCPaauK
FRMBCEbeE956IFXyya5NRrIad2BdfDuRJhSVqsSRj6REd0E2dMWFidsFyo3UH5Bd
cQVpm+LoEXUhCo2gypyHp33OPXU6rE5vkOdDb1O3G+/30+fo9v1Rnu7ev8LEixg+
HgiZTRy1NyB3xMEjiiXcOmZ13la+ly5FTv9fhWvwOraSiaAu90HCXTi7EnlLIUZc
CZcdcCo6Cv8yQwtFf6OAvGm9xp6CCBPMt3K3XnGNOJ3SShKFifQSatSi3ygivrwt
3PYa1J/AyA14gB2sdi8ETni6dq52wj6JpyjAdHIEi4BnzQ2TX9Fjca+7iJ/1nun4
pap+WmqwqWx1NZWELI/b2iuls1EbTvPN6K587VHxu5ZF39D/Pbeg1gsINv+R7W8H
ZnTYw5+PrJAPDlhZccLT+IvwRo4pk5n7/FLxFmBmO1fH2IP9zpx8Aq4bxicCvdwZ
E4CiPtWdKe3Eev9LMsiQSFthMc2WlQZ3/Qzpu0t7zo7MbemWAYL89xzsBfAyraoV
/VO//loY87hiDDOYhkxDDpmsqYrjRsIpDT2zGmQ0AtgCPi4A8y7JFdREueMBRJbx
7s9sQ/lVk98i0xg8WSIZQqxZr3JsLQg+ZwCoI/ITI99oG9HCsqYKrXVMri/n5TGW
v8iI4DMryQW6BTXNyBrHUiay+SE2bAJwdSJP1iW3nJW3FYVXZf8zZcRYDbzW+QUh
9sqoD8Z6vWv96DlgXq0O8YN01p2SvNLoMKxfxGqSUXZ9htfe3mzgUIH4moqdQoaB
PT/Cq1PKOLhmMWHiBH2KgldDDrHR7ctYkiPVn2RIIlTsyv/kIGyQh/v8tWbPn3AT
DjcyERh7EHLLTIfs26Eo6kn8RqvDDyL1LPDAMA4gKuyTy94bjPSiyYL4aGAkyex+
lte36NrW+OeBC2Pj6x3DH3LON1/gxR5JcL/2nImpXchnJ593Jkx5EWSgqdUjl2BK
3gCPP3YLrhI4QMUnD8bAgK7M4PJdYVLvg+CUpoASqeGuKrcqr1t5msrLtNoGqsKr
eYMVnsgASkAstJBjYuLZJwsZ73OhOllyWpR4g4x93lXEWmv1fk/oZd8nu4Nt+1Pa
4VSSD24tTTEs5+I7+BII0gSH6u8iqTWSfxwDY4xDlrrAtdVh9TplA3uAsXBPNaFN
7y901KLvNjKZe45rfgKVpb+ZccX/ssA7B6kt0/EfpIhrOg055fbT1stJUlEXG5XI
0rVcqt6k+X0QCwXWu402jfHg4BKR6ah48YuEtDSFhgysM185e68xka9roooNzEd/
O/ypPo/rWSrvv9FGLY0bpo9ughfVvtqcg+VjgoBoKYaj/whPj8LSc7l6VT8CabYO
2ttaWVRunB0DgsqUqqNu5xfT2ZbqqFV+v6EDgE+4SJPYFbJ8VaBGQXi83gxSKmiX
3jqUWgjUsAhlVorGXIVoUctspVgAizkzlgRH7dRgXYAXNh3uLKV0ulmg4NeeZf8X
8bObDnbnspSTH3Dx38IjhvBeEQzz3lUQPGr0X57jOyAvvIeepb/+0EapV1DAb4Ga
hZ9+6jDq06hxfm+X32Uv9JuS6P14SFxpHC6UC5qI0CyWBO4y8yYw0tW00yYKv4O4
ZckjOCgCfcfvs2AnHSj+7Fl3cxgWpdcEpAg2KAG39L7uQ4WWfLMhpizKISFKos7N
G329GJpVldLdmHVbvK27OfgypHu3X85vn71s6xMZApOldwGXYZYVanv1fvcYTtoI
gX6g2XljScTYqFQcvEFyItVs8M120EXZcjulD87Ku2gk7IeAkJxXMAw5Gy059xi6
FBkl3FNBhjO+LD5GErM561WC60Myc0b6lZyTb/eB91rR2tBXZofY8ZIQVXpbIz0F
Y89gdPAbVeLBlNQFABBBpMXHeG3KOl602rD9mXwS5JA3CqV9zyd3vnhvfuKFlWwC
z+0ZTsqchnulrQhoAb5OIXS0pP1uA4ZEeVuYZKXPVaCdOqDHmMnBkoW6DNjwLL6m
fi5TUZQAzC1Jmk53rqKef+1lJF+Ru43RNlwLmUMlRsasUb+d/uXG+I9d04R7gxIw
4bkfoNXr9sA5yeS51rzq+jOx2jnxIEIJ2XbEvAPTBrsl2XypY9+F/0eIZxTDokMF
PB8iyf7nKhRuOrO2u1wi0CmZWwzeSSD/Ykp2oh5ckKrVTXdqH+CRrxos4oXsUQED
WPXsyaa1y+reQwi8xNQNQ+ft1o4J+asLEd8ZQNaojIVAlkUk2Z68bhhJo7IeKUuw
kGZ2ddP4SHwJw3ODnWASSu8K4WSweACxpTyveyU8/afVQakiJ59JKKtj1+VxdcRc
qDplwAQl45m2YJ2MTO5w6DBkjK7nHgdNAbT9SxzYln1pVDvXeZ/EiB5k5ESABrA3
y2Roi4DPE3eWE4hDwY4icbLLJrNMmhWGW54QVGcodujfi0qN8R1c9az/xvb+oRhd
IgZROQtv+yRUN7LcZKAhJ9A3GFFTz2xbh5pu0Lqupv+y7eC/bQ6svc47Lw5UBNEf
N7jAe373m24dw3USPKUuSBXAaNWBl7BZTbBzjN+XbgKofbrB61YY2QPuE/Ua4Jnz
SIhPZgQALexrHgcOdibbAcGoTse+3vnoLMqVN0jl3hMULwB1NN2DibuJjVq1YyFH
UfB1hs1lzNoAOhJVmmt1BDR5EqjRzOFRVb8WzNo43sHF85+1MOKSz5dMckVodSM5
sm/0fvW3C5/ryQjk8ghGMA==
`pragma protect end_protected
