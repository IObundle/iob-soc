// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RIrmQrZT4gQqibTfapbxU48qLvkr8hDrRcUYxbBy8SrOqYOMW2JQpkmFPU3r6F4N
1YipMYXBQ/vIo+3fs352bFTcnlIsn5iKpQyHbOn5/gb2O02oOnmM1h+uVNV5PwLX
wKZAv0ry0+udzzyxGPNewvp36GDudUfNH5YYZOjKsdA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6352)
TGNYQyiKY4LPbZSADFqDcX6eR+8/+9PhiiOvf2+zOjPXUWdteJNvHlbFD3yM3oUU
dwDBz8gZ1ydBwnC4Vo6rvpHdn7XOT51Sr8Wg2jvxlow6wV8BddCeR2N1RRy9ModW
HXPtz8XmOhierGBvgVBfCDkK2xQYaaahxUmuI2CdMFirHJ/KvtoQsnGBfpOstoo7
ABbC1j8lYrVF/96NhsGY2/iPfpUmeKPTS3ReUgRZ4UwdXe7b5Z/VrcP/AY114slo
8pYit68dskUv/KMOYH3LWhE4CiDUiJJXNxAV5/wXg6VNMHN3BYqSItq02RXDWFd9
65w3rUod3Cz8LYrd0uYMwUdOJ9mq8dtOg+7KyBIvwiefHIc1YpVuQ7ecE7XuuSR3
1L1wxAzHjvYHyDVOQ80TclvCviEFLU+xTeOFuf7x5HndI97RxsD3BeaqmD5DtBol
fEdoHdPGoR1ILDQrcoSiVRgRwXddt1LFmkFWZohqJfmJXzf3c7ZctnZ4KZv9/PaJ
W6M+37gZR7/TfEZKrpghU2AfJyp9n2muykGuNy7pNsHZt+mBIIR7p5CNcX36aABL
F3LgWlus5LPNmqWUkh7t50XATi6tzZeErePlnAQB8gHgAH64pn0TpHzjtaMj3OzK
D4W/kSW3y7J3mLj88ZshFbldF1EBxLtNZ0DoakkQUhQKQu4q5/URtP61gD1nTHWy
zJPt4b/o8h6A7gM8THH8ZtFKKkA7BaYEq4vrIADl7Bqxg5aWxxebDdafAPOk7m39
fR45bI5h3MPyn8xob3Lnlcltq/runu5QH5c64cbGhsRl4aB+5SnCaRrnQgwxJ5og
q5/wHsMVbJ/YvIOQ2XSuBzt7J3eSGzk7ZJKCRJHL5l6i/2tY4E2e/RdSLkFwBlYY
wPoWIEKxa2xmnkj2q0wy87zIT5z8eSHXM8GnojLULjl/eTOHv38NpbvX3WWSpkSr
219tC+8mmo85s+Ui2oVidgtjpdzqCZATnbBipHk3kDK2w7nw3ZkI94hduqkxMRQU
aXkT7E9H/2BRy1bKxjt1u3E3HIf965DBn/3rMkvQdZ+dzcFO/EpbWeDQZN2GLsjI
9eYFwubEWq6sVcru+yhBz/nB7HlKuX4WiMUAJpU6sHru0BFbPChDfaC9fLAQnDLs
PUmYp1HOQKxKaJD9DIEaYzg76HI5HfJibgFu8uy3s2zQHEsznldrqH2p7RLbq8TW
u9aDuxm4my8BZxHZMw/HGLm1xgQvG8t/2wNHv8LTHzlbcJcRH65AIsEEyefrOU7d
0TlrooLyncqD4ZDwmhtTQHPrHecP1yEWuCYjibumxj8tiXt2OITtsAQuPTHceCXd
gsPXzpbC9z+LkL4HptBHMbh4eO6cN4JI2OJD60UI3RyROfUULeVD+kgw0S9SmRqL
3RISGRgeCh4YYv8n8sJjiMN+Zr3q+yqVJ6/HArNR4SbLHSmeOztMnmQa5B0xXFGs
NkBqHNVLxoFkAqoLWSFqVm2As6bzU8Woqc1HZB+u1dx+fNyaZPIpMXQuqZi5yp9+
unz8ojzJ5WT1Bc8d++K/nfD0jsw0N8vwluR8ATG8nlTBeWoEXPQh9gfiPzw6llkO
adDSTWlkEo52wHywedMuclDruQTD9CE57EhzWFgD0FPutm6JgyOGHWCcSUI/UeN4
DUA1mHhtqi792eLwKkDMZFRZbaVuSM8KcTX+1AuAVLYe1M1PugCIDEYlzYQhlgv+
nm8bmon9TLAXUVX0HuFSo03g/b9uy01ILSjd9HWBoY3gMuu1Q7rYhZrG4BWQGLGC
Hx6b9n0Axwli3VTIhL/dmBsv93XXF3Mmtb1lLG2K+YkhdIft4Ur4pliuDRLNAGnQ
lcFJ5Y1W9yr9M5Y7OO5KwM5TKH6SuEA6AkkbUV46wuyV0qg9FYEuqYHJVfM0iDvO
unekCmF/iEpec/3j9DA8JzwBdxfOJWRdsHV74Edj2DLCE6ftVVBoHLdLxIh5Vb5t
VTzAfI6Xhr3eKpSuG8VSgnLID8cki4tk7/UVUAa46V8JM0YAC9F9AK07+h/RZz/U
gM0NADyqsdf/gN7DUl+88Xkg4g0M3Pimfva2tQY49EX1ftAeWIoBKKyKQYpadU4b
+OXNLdYJzPNHPSKYxBSHK7W6JiLgueRrEuUnXCASaliLeY1z3uQLlQ3TsVBhlmUS
S4jISqzvtxLV71coIW3aMxqahLFM8H/bG3o+tf2ff5EaczgJiLP5um1HiHGYI50m
+f2PV0prWai1MZ9HAHHLRs4LaMasObycZcaTJBWzPu59BxYDWpwvV6zhWwfGNCF3
Sgx6ACus/rYVg69IyRqORtAY3yMVcu66sh9S9BB82MfT9+QjDyfnFdJGn84av1mL
0U5i3N1TfmJy0L21CLEjnOA598xUO+KmdoVPHS16gyWNwcv7bD5ZIhM3eLAmax3+
Q+v7xdHS0W8+o88pUtiiYANuf0jpVZ1ACSrw0s5tTz4A3uAaLbXxCaGFzqcZD2R+
nldGpMjGgT0n9lqP23vsAHxpEz6F9QB5ZP+mttghG0nN37MU38D/hvzjO8C3TXXZ
eUebsXUddXQNTMHV9pgDhHXPqZqteqYbk/lp2rfDJkX6SAqT22GzROg6yhxIet5Y
iBzH1tBVbuotCTtFRB+0xze+mZ+fSFRu5PP/gMfPnBTsCEMexEiVmjfuYe1UkQZr
nXlM+aa8z89gTRsUEQ8m3WIN9nmr2dNzQiBSKfDjYzugmmyIW/U9Td3k0X9d0dTL
WDdNF6LUMNyNHPQ+OSt2G2GyYk5W6pX1YwaVP1s8qSuxSamsdtK5nKh4dr0xJdeh
qiMYC96659bpR+zXp4kpGhVWCmxzv0hdySEwQ7MJkvLbaSFFitQ8uaY0K8UX4B4o
PUIL7TyZOVee4kW6BfC/ITUuJx5cFzlth1IBfcnagKDOnN4OUbxb8cWCRTOkRThu
ZSHrXpGTQK8WHFCIBQcQgiasFSPcu5P8WjBm4xCAkC5WUtKa0zJZb+6dWOcvmTsB
KZ/ykBYlQSx/2SaID8gXvAiFh2ivnbfU4vBEDri9n24dQ6THyyLC1w1raCQofpNT
OidMUyhoxSAcfuQuOryhEQBV1WDCV50Cm0XwEV1PL3x5Yxhr+YLUZ0PeB461EkEs
ZfWIbhxQ1y5XDPUs0IxioJn764bqVlOdQCS3yDtTDY0wsMAgv53wFU6Wu5C/YpKd
O8jT4YxTmXnldDbcoOeUqhRgQrOHmK5HOWD817Q19I4GJsrnBkZivVzdLS/mw7Dd
f3CNgBqK/aUDc+rIhNNZ7rT03Hyepxc50czpXcGeZNdQRwHGn98HZyM4Ro9mLVi1
Ac/eHC10fdqHo91msSN26sfQQhdHSKwUSq94brthY6Ct1DoxWxqbTR5JzWXicBsE
WeajJQ6R06XBP8w52zYx9/tr+NA1rrtoI02ypkONV+av3qt92XBx0T1LfAgPnrDO
4U+ZGWQ9rOyPRp1XGLmVFkmjSiaNMve9JK35e2F2/C0hKWRcWjkopmdRCPbvkpoo
CPiwTubTDUXpSXxjVoYRzdxNAxf9NwAiwWFyv+U79x28oWA+E7x+a1MFISf/surl
KFawv7rWEDeLEYZ4koUP51LKirPSe/wIihWOAxjKFhePp21Xj0rWcRdKjZuuz4q1
N+xYlNIbjpeJ6VqNX/uGKl16725olT+q+de3tiBlPusa5/Nei6Zg9HuF/QZ0WW4w
35eS7d/pljb9qKmCwBnLsSlJHCpwYtMN2V6vhE1W55sgecDisC+KN1DRM711VOTL
351MMT8Sf2cux+l2y8DEr31Cq/SfS+6W4PjKkMgB8o6O/q8U4xNlqsjcSCuYAZFE
3HQ8c2bonagNIgWC8Lrq3L5yc3BtM6XOqVJ48v4ip91RvE/XgJ6/MQYhzojsAZ8Z
wUAjaP3kB3tCBeJuP3zgaACFr7rkwtQNQf/xjqoiUa9iH+nYVCivPlWaVEaMaimz
+OkrCercD+hemb621ZdPiX4QwiL//+sr8UmTSWy+TpuuQCEJacJqYo9K2AHP3/5C
r1ew1GR9XWLvUbNxutAGhh/Px5E4G4yuyw+WM2ynNDzG4kif/VvqXNJAOWRxNubS
eg6gFadsRcNJZ8DvYKtSLMjXCqX2yO1oo4yxISFmIG7SblXU+YqcjAYwwAVbyLr0
MQLpGC3Z8jGcYqUvjn6O/suWxXcX+ZhMsNHk8vR/qMvTR8RCQcI7S4MNRyYeGLG7
RsTHnFyBNozr00FPTHEdVff/Ab3hvwCExd4gzeiHo7kQURq8GGPciUuQ7tkUwVRC
DMK+ykLrE5xYA9GqoYd7BP/rdEv/sSUQK9tb2jMNwcWL5ud0BtBsA0YoKneRVJB5
lbvVKG+jHaF+4MW2RqN8WgDg41XqkbHXRDzEBNgfU4Qz3d79Ek0o9cxaKrdhXo+U
Ecjzb2mkB0VhIT+YpUKL73hUv/Q+z5kFgZ9uwNCYueHdOvG4VpyCnNp8OtnLPbuz
nRXd+uETZChh2jnlXTy4bhgPatijelLLbJ1DX9kPv8wHLmo536GuvWqOnP4BqFPA
rl/vG2nyYs7zNsh7m++1LOBCpoocEoVkPI5r6nVSp67lndEpsvdA0Dx1g98rK8Qr
PG3mVn4ZHONf2zLrVAa5RpkCuxgIH0YW5p7tdT80fYFIr4bMIDYpK3bWgQ4iJcT+
69FjO3PPy6KW8h2txTMj5Qduf8bLTHoiJ7+eJmQm+pZjq9PVuva0x8ppmBVTUg+2
LQH8pFVQH4o5cXme0dq815dXDOJgElZEOSwPEZxWZq0o7yvksmvPJQzSCgxGhTCS
9ErZsgJZj/JpTpzopN6vfsdkY1G691zH/gPC9yczCkXMQCRKiEO5K1IpiRy+UsBn
UcWaPQ59Si10GBtFA2ZoYXLTS9echmS+5t1MpW0H3qJQ9xKeFfCaeZrn9RZXqh4H
cDmVvjDZ37ENcViz1UhrpWc4DwBp1lLb8cKYEK0i+PLvUnFH6f3suWZN2tLj4W/6
bmy1FlHDAEXuDyO5cRG3eRtAouxpwxCzNmRPgomk3jpfGhJ27l7LPRqWFDk9oJ/O
xUOHvhjNgmHnSMWwcoujsKChAriGn7pg/Nnr7mG65fCMDM+RmMcdgwkcZnJpBU0h
VQLp8cx6HZULgybbLY58NW438aReoKb0JrCc8QtEEpkVkQLdI3tHF3qHt0nVJ03e
hW2oakgvn0/XuqZzpeHmoDVMsHlNH2aBG7UsURK/YZJnepco7rOe/0qS/JDaQS6D
BfsR+NJJqX67++lnPNPj9m6L7eo6poQaNauvjQdy2asolQKNxzYoiQpVr9MpUMXR
v0/wn3QYQbJ1fpAdocDdS1QpHuC/shipz2IvJOCLMShvb1T70uRHDgVtdoBkU6OP
9M98jw16auupQihoTVSFOPr5lNfFBl4c9hE8XNSFM6qD72SWG9YZNK9hQ3DJnFKk
5SC5yZeZd640V6tf+HPcepD63xVfJlYkUcsro6vpy7oZw4lHCfGnWoqXBCy2gNyR
7JAP/WjUt/i3uZwSkhcMEBqUaj9Sn481iw8+UOnH/JcKv74eLRv0qdiwpgczIk6i
xSzBQ8iv8OVeWyZyWEksAw2q5PSO0B0lgUeEJfKK2Y7OqH4JWjx1h9qWUD/L8A7/
IxGV8jQax5U9AjRXtjbhl6IJGf9A6y+khCyFNIDqL0kLSrath2OiXUBrvrW+wMcq
0/8ZHHCNWudRwvWzDaH7Iic9jJO45VQLVfBlCNGMSW/6a9vHkN+U7i+XWnpZCsFv
PoklPWf1GQfA4iE7BNzZWUq4TIZPq+QE5/pRxm+o4YHJ28OyBZSY5/axuehzij2S
92xvZD2f180GCsK01HpNDcvIZ3eKqjMx8XFDuJqxq/xYSOcCQzaughqe9Oi2ok0S
qr1u21Bky8498Rsf4vOr0VFWrHSxOLsqbfv6jPFP2chUw0BePJzCTkOgpfOhdCWG
Vk5/i6zDpGoG0Jj0fPkGcmSRj07XFC6DbOEItBz6FpbHf0JvUAQp8NjzzeZ47wX+
Hde8Tk3phqGm90ikrMpV3LiN3XJn+jOL0vkL5HKkRUB1KyzOZVMwPN3cmDfUNYQh
svkrbuycEZtO+1Qb09Fsz7qIfBmQbMic4p9t/7jjn8BbELzN4wqZ4ayY17FCXuiQ
+V9V1eNjSfWHrvbtLNtdeOsC0pxw7LTupg3uapU56rZk8b03rXzFKyi6HN9xTUdm
ghsekppoxJHwm9WxKrRnEMKyyJ51cqXcLKuwGNi0RtcORRyIfVQTCkY8iednOdRS
jTsE2fmO/xvPq08duHoLBsPw50qePkJcnqMwycDOCcKjArsKsG+zyfGArlCijQ+p
DRaJxrRQrREVCFFHLnXEt9H9lxYFGQlyr00xewJuAAHMUdkoOKKCmvuv8VAOUFBf
Il4+wzSWIzX37Ll5ivNOMGPkgBp9lp5HlvTCBARy0hzCZIhIWQIxeAkSb3dSRpu0
GVpAa5ZK/S3ttYCNFkkDLzYrULawAEhgXw3fam3iEegLn3mMqfFxhLJ82jtwq8o7
3rxKNB3u6SArOKzOdK6osWXVVxvU6mkY5Q6cHYcjBuC5bUeDaB+W4wg5ldZKsKVn
4YUnOn51WXRhI1sj/Gz6nQu/qkr1pcKdwr2Pxv9QxHEvnUP5vK1I5pZSIGov6Jyx
IXDUTppV8A47Ik0A8nv0dSQlwEtQa4zlAu+XSbvdxOZRtZ6owMyb95dFeC4DX8C8
2EH9T8jQm0JgFySjBtRls7ZXQFn0mvpGp9H7ztj5vc7YoxNCxup+6myfQDUBz9Tk
+HYEicxoTRr8FgG+PkelLJTTswTBs6rOu8GB+6X2/RLuTRst09Mk8OlcgxTntCzL
Nms0IjYcacSskvevmgTzBM2ixoMKmrDyGIa6Ck1byPnOlJLVP1xNwP6zQTyfaGY8
+Fp+RFZCpar72Hf07cRjB8/u09xgHkt0R8SDan0J5QFbLTwkLVHA1Q8P7TE3em4J
L2ZbGSUGEvnxGKlRiAvLHo6goWZRj79CnVmODXjjS1nxdH/PN6hyrOrIKjkWdqPl
sgu+NZFnPJVts0rwg8xRyH2UCZdaihlODnIliP79R1B8bGqeloPV1Vp1D+CIqsNU
b/AXUIgkaqmfh2zb6NNEsL9815RxpVI5TUG6jio36mNHeFm40PUPdXSqtN7VgrtY
TBliw+MMeZJSJe/q/AxoeFVbczB20+LW0R1IT5wFPlCo7BbbenN8o8My4Kc8ZCsk
zZlPco8a/UMkWzWMcEKFiUDrLdg0FDKWZz4/5yV0EKqMsd3OYikxijheDjkgRQxi
TbYQYoYbWKz9qy7ZPVGqjRiueVsqTjZNUo0KXOAIyPHhjzFOw0q+hpxUQd0FDX0s
BlyP1Dyx3RzkLEcDm4VnoC/ETIeFrAIBpgXkytEDWzby/yfAODhZ6tGPquqaPI05
nds4V0bikE5B5NVoHXjfvT4qBuNDJm13eAQy0Hrdif724iQatNzuchGhfkKxKA9J
9B8ufMcecjfbbiQdMTMNa0v6A6Pp1VTkb0g9j8Xe18jPQU9gPBkMFPCMJftZkm9R
PrHO8+iqt0sHYs086vOO4CxZX4q8Ie2rV8VOjiknxoNAXequ9HrOORymP9IY4r9m
KG2fsObvid+fN0AwGGZOm+EIo/eq/4sNmhuRNSiKywMXxk5NxTacZW0nkXtjSanW
yvMla5o5z+vbbRLsYhsPf1P8NOI60JusBWmXl+Mdrvyo8HIV3g5hw11Lvx/4APcl
WIXpiPvwrx/kXi+C8S/9q63+/Gf7KlH7U2320q2EdNj3onPQHwq0ARes9pz6MCFD
a2CEizIVwJBwVYoI8pwBBrhllOXShpy5LS/a5btCQd4zGjZHIpsWqFVOruqO7Hvv
GY40iRZNSkz7R0ZCWu4lbePAhvXlK7cz9R2iZrDV6TO5h9LJbWn2L2RgPs9azXg9
q8H4DIMH3qVijE0Ly8ldTWzIYPei1ZTH5aAUud2jfkNyGJGXNPXeb/LshZdlxHjw
GRJ0K4Al7j3Rqso4TWj9DjhKGCV0UMJ+kTkiHO4BV+UZhxR/QWxFjxpfoZOc8msj
4V05h10T9UXcilJiwUvfrxI+gbrP1xi2o0ahH21rQ52GihmMe2uNkKyA0kcgZjg5
Ibk60UXxFzuNd3ctJUSDwyQdGah+dvZBYUCsoUgohAXf42KolkiGB1CWaZxSINaJ
FGHyhClnWdkN8aM/EGK1ijERsm5sM6Yta0dGQUbY9uHH/3yQ6Vp/xLK5wvT1AKT2
fB6iCbX25g37xXn7FAW5zm7UuSbEqD9kwm8wXPBEmYqtSvotHdMsrrgBWCSC3hWv
7CDh1zwnnVBIeO+zxIROzp3mjpg0v3UByXR7YjW+IvR1Gyl1FPXdpZnpBWXmSaDT
Bgad8iGyVA0uJEyz2fbIj5+Lboh5FK8cKOIdWPl5n+iZq3M5kt9JT8IaKqYiy/s9
bwqIZinSt1+nUWpNwuse8A==
`pragma protect end_protected
