// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F2LxgrZilxhKqVRCGB1DxvpwsDk/4Ng9ku/sf7E0Lml9P3O8X1s77/YaXZw2hmYb
KDmBMGlmxMkUgUfXyXe1AVZzJps8PjAyqIA08YDqP8l3enTbZ+S08egvzIbI3c6H
OuobpMVb0UxgbzKkpGov5BMqL8QluaJRoIA+TB/VGxo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 59200)
rVNKScCrDtg31RmfQjRpvGBM/87YoApaUjoTra3k2QbbDmIx4Ua1rDKsdDb47N7N
EVukmZWSuBv8DJ1tInF4vD5t3Pw7fr6oNKsifgSmUf9+hM0Zdg0CfWqmPJ7bcfyk
fnK9zHjVhxi+LWXOoht+XVj7HtO50fcUubshGnaq5Rcu3yeJepc/fur+vNY/Rgpc
hO2tBhSMWm+/qxU4LYzi60T0W4w06ST+TcvTPDDHLtcQp/NS5KZSfI5U7xegu0OP
qdSbno1p8ieBpDL3a4aaMcnoPTnwS5ZCesmqP6STQpmIInUvdkWM6T3u2xtnxiPi
7w6sELjWr6ymXU7wuPLENYKnG57P9vV8vJiIGzfgdhaafNXZziNB6CbCMdHYMDbx
j2DWGKkIntgdJGPdM9XPYtrdqt3YwHVeXwxVCKU6B2//GDXdhf3a3HPXOtOEI4+a
f/I7NAQMRDArA2/hzv06humPd2sFk4nwYCHwSwtCoabezsK5pAaDK26SBqyCMaTc
MrUIZFdwx7as/ePbdPn/3WUT3mGx9X+8CldnCjA0LQxYxkVtCpBo6vEnc3ZdFnuK
S5G/Kg0c/+7Yitm1zMKXlnQWMuJprRJJ45JN/czBEshfqoDaXdbpwRABtFl8VFxv
k0Siu9DbiMdhAJfF7kP5gSYTiLcYG8jG3CRWlF0hrJbLc7eY/bdShJq+W5Zzpgdf
7JXqOwsIXbh+Hghx4wTMGDxOWdT0l6/J22rXeeyajzTsQ6aatZ3356px4yuVRYUD
SINbE32eDutLISc11pPvAtd80V88L/d3ZdUp5hxG6nS3mo55WmsQr6hMT8YfvRXC
vwJL/8D+o+MP08WboQc821RGkbVE5a9KnD2v9uylaA3Owk2Pd28w6UpaRsgjuNYm
C5v24S1/zmcZvxYYoY/hb8bkyvt6bWa/8pp3FuNZoObp5QdnVk5XJLZHkYlSDZIV
wQaEE7PPGH5jAl+Nzq7/g+3BB3sZxgEJzKN+4LWLHSewp/EkvpW/staJuBczMtxE
k54ztpxU8kKl7WvaUGZv+goiNnHj0vG4VtSoWNKzSi4uey9V9lj6ZMq2BZuRpReW
Y4tfBVDdTbBjAleWex7s50m/TWk0a+HdSeJhZys0nC9xz7g54JEN56kievF0+f6n
LtV28EVB8gryw7ygMwRh6hBg8Xx/uyoDHu6egRXOfP2FCtUgvwJRwfSHdNOYQjhY
5a+Tb2fdVBwFKVqJpARI7vRXNKHQZps4BbrVjYK5TcXF1aES2WlyjfU35frDD3Le
bC1tqMjpqg2s3v8lcUxwUmsUKj81lFy2hVgA4CjD+wWxhQTO4GV2fYniRf/0u43Q
nGlTx/+X4s5TnD6160c8/KQVNHL/x9gBsDJ4RkDwnwgCPXx173odqRgvbulbZUVR
V4iv/T8RbWjVxegWfoxVXnclPQMHdS2GbZ4Ov1ZaRwL0Z77vFLvf4dYRe+0ZHsQ8
NOc5lvPu5OrB9OOXMJXIU3TAE1FZrhJGNW4VUgAWoNDRS/AejSEiuhjYaEiNZ8CN
Sd7/v+zj0BUFh6acPbD3vYqdLintO1cNh+8IZLRVhgrsNYUdoXe6qTDKPjWg0NsD
+OTdPkYnEsBtdkZ3pODmYIxe0PZcL9Gh+s3uNjBgH3PWx7Y8iyY9BxVSAwl34/Mb
Eqeu8RXtpY1tB4lRBDmPPYaaPjE2UvF7PprE6GkkMjYF4veQMm8O+SDHrwBgBPqs
Gi7aIM5zTQAsERskpYo8RnJhvbTdlWQpHDF6YGffqyEX8hOksIPJdxGpI9XJp3zs
gT2NxwgEOMNYuJWhlTDdaq2rFYnMSnO+k7ybTr9ewpg17qxrMIdXR+ZTCit/wUi7
tydIeuQe6kJt6ND84Yb7KZbpUu5UmzuBEmCUTUmPNZY02yBqik78y4kWjtAHGnm1
6CHmZeA4WmEY+XHdtzYjqOs3FGwlHG/zuysVHj8HnK0fVJHccEooiIwBf4opvkM+
M8XGdwF5uk16JizrJlmaocpkinfynSzT9TK6efa8tCvqJU0FDocNuiNBQ7YUdNOS
cSFjmVdiM3rhwll/VHuZirFz8mX3cLz1PDxcJ5X1vDFF5p4nd7T0wpOsL1Vj0ynf
eguVB8ixSAIRmyr89ij5EEyCNO9RmiSN7ijCKzywS4E/2WKUHVeEiAfETJ77soPJ
DQlPTT+2PfF63aCDnlF4uKvii+ur3jzNU/EeA3Mg/OEKJY+Kr4T/ytLUMx4Ce6oI
lx9dek/FGw2vKQy36ZSg/nLMZAeHrAG7sO29dcqY40aqclI64rriPFgbgY7+eFVd
s2FFD2KcUAiH/rteC3P2cC+6Wkd9m3AKePLAtjjiasRs51M0NbZowCMDT/6Sx6Ub
rh7RAydvCpcD4bHnTz67goLbpFdcdlRSkgN/lW6F5FrgRmasvUOQCVjvBjWhKMpO
4TnNuWTOfFnXzAfW23FiRj4u2inb4Ld5x/5e4OdDUo19yrkWJsUgMGZ/VfoMmKWs
CrSdfkxWzJDetGntUQloROrO0q4mTF96onv3dEmKnEN83UdayxoDK4ILHwSJHcK2
0cFqaxm15Bwd6VNRAclT75kHM3jUPqq9Z0dBY/RglZ6Y49FSlPd4tIqKyfwjlCmd
JnMqrssY+et6dQP5RJmeeTSMzbBu1oktIpGFXNiwWrG6Ux3+rfHL57BH0oyiVxEW
sdMjXGXgPfl0/QNhNbqjkSe6yWArKC5pojhAmb4rb3y1PIk8x6N4Iace8w0LxMLr
63M2mgxLpGgDeuLeHxdPjxhoo6a3JGWrIF5NjHkZZRMkIb+YjiFBe6TfMlpxdpcj
jxvIlz4moeBQU6perp/uR6H6Kj0GHKWjE0ldKP4LaYqsccC4hjdrryvNrnhoW8GH
nJNi3gessFspK0VVQfht2b5um92X/j5DndGI3HeD0cKEie361FVf4rzNxcDjUC9h
OCKUOfximJs3JQs+3pB2Q3ZoCosy8CrhcqeSfiXKFtOrSSO6RvWGuzuppK8kH8NM
WxB3YJt+MBtFlGC39O2UPJjNbY6lFmjVesoo3d9voAwBHlNDnwrnHcqsMag3kYMu
8vv6HB11HHZA/XqJvSy8zV606nM4FUh26K2zKnO638YFppej1bY0AS1Np42ZI9R3
r3vzX/IGEJEHOxQwpPMTlYbBpUbffqW3wLO85QD+0MKOmzi19q7mxsuOZZttEkC2
AByi1QBACREYcWsd18za+kO094+4QdbZzU3jjlx8sLkoik836CrpHgnOP9hmTNor
flDPISe93sXDLKque/HClujneDbaMy9kmmjPO7xj5r9N7KIzgJhiGTRqDi3ejBX3
ym+5VsHH8mF0pPiaWj/jXn7/rdb0wTYEkRq1YUUm8C4UpHlfZ/LmSA1DoCfdpdw2
hm1kLeh7eHWoINeXKTIEUQm0ynbXexOeZMrPIJxvrc5d8QbyHOYp03saMG9S7Szm
NUDjUJoS8H8nseoob4ATZDuKFKU3puxw1qCeGM5Sh0kR5FTNa7hsN3Ezxn+ImVAz
nRYd3JKOFwVFWNiur/CxSVD0gvo17Ayj4N3dFGlGsW3lQ9PF5qqZuI93quEmxWSc
8TBgkwqf95TLiYyqzENQux4G9cid7rBUt0VI8ZvnzWU68nGdpboghsuCHKR2KgwI
5AOAkm/mfF/3TtHrWi4YvmK0PKPReJSe2xhK0CSHpFMng7h25vWg3pGNFqlBDWGT
l4bQ0CDs9I4smnn8K8vFBFppUMqsVK+hvf3D+QQShPaO0tyqZfUIo7sYi7oZ/8M1
+yuF1czss98GYP+f5vYgh417ZMe4s63Z6qzsNPSY3yB2NXVvuPLPOqJWV0IPEvMT
/E5jQxRiUN33Z08tx7viBwe2IshRkG5WDyPGFzRj4BP73XxBjiu6FGlhc1rVwkFT
Pv2XvUP5XnHmVLIPBi1206B8NF7YC4vYfl7n1Atj1r/bETgqozssfVrEunz9mmxd
DuyBSmNclkObatswvAxKlsbXpuD0/g68PXdecQu+Tcue06KZ/TQhe7bRshzUMvar
eOulGa4yJgg4xBFvVyHPT0ANRQe7tYiyLVUrU+iT3NNOgtS+mtO+kVSvlPv5Ho9n
UElZWy43mKRA8Vi3xSanV46DRf5JwU3ZFTroLlm3IqOHMjK6iNTp3qCfm9LBhNhP
HdTXrVtFviAVz5Pq7dyWsdftHLYTdT3Z1ix8kmpo68kBkQ1BvlQ1cIqZjmKfXEUy
s3iksxg6spYAcCn1kL2lhwWGQ0MnV4Jl+dOhkU4jUN/sp1+oqGPHchGIDNwFngNR
PnoZyy2V+TLFgt8HnJYc+h9MNquCo2xkwZcr4nOFLR3hm1jPOl0ilt9HoKhE2NgS
qd6Iuu0G5ICBkfH1+MeRK757wg9DjymuojG7WSwIPXthR1jlUJTY0LEsXccICkBt
3yvTXc62z6/sZii7tatfmJ3aVNYVPSff4Qhpy3fKe/G8XWi8I3xK91knU5qVun5K
+sXMMClA3PXTxPnLYn1IgQe65N7ZG5QRrqNgREqKbcTUqO79/0GBUhgC1TsCrBZV
Dn/34YhbgqguMntIhNXOYRv5mPfzge/DvZOPAqHWPiXYFdJ03p6CR4I1gaAU+Div
eOlMW7hT3x38L7gfgUurLOvX6DGcRi7Fd/cphzTRJZ8pKqsO0UKLcrIiVMhNSVS4
+DLL1p1HH1sZ/JVszutv6AGEVDCi2ufHeWLDopZDk/fl5KSduKKADfJyZMH4PLhQ
BL48x270A4KbSzWtc1+IRmPuMNpEMjh4ik/NH8m88BCaLU29q3REj+4gW6wpgLe8
4I+Mb9xsAmSAk+3ViAwAf6Zoxl/pwwFRBJCtScdP6jd8GSaFwwbsPQ0FCC9z+Z6c
5X6G9xeU6+MT0QJwLt5kOy3Tl1/dRYbF9hreICMeN3eFmtzbyqRZboWjwFnkHtxa
nswxfG3oYDhIOIWlaOKlX3Z9MLwrXtfgJljeQoqGbJk/7OhJGKo2QZCbHg9DY9Jd
pQB6swPNynVA5ktWEvHU1xbOLZERmwY6B122zcRJqUeM7RKSptD6bCnMQumWplZk
QivUQuGaRJ2X8uQfYw83rRsV97RYo6edFr7HFV6Ebd7FTy1VrMQLdAgoP07YICzZ
omUBKmXodwW28Anm4anUNPMgdBRvDssYqkwl+7J5AGyONE7qKSW69MhiIlNfsxAl
FfHedANVwkeF0NVLjO0PUobskSTyMr6iwOPkvzSeTxVyxt73aIMJhqArxTVd0be1
OuzJzB6YgxYVEcWXvIcPrgQ7sSFSX11TTS0WXBx2pEYeJ2jxhCb1SxI91bAM2BFI
0G/F4R5FMe4bKF+o8APIyhwDIP3M3v+Qv25sU4bche8VfJIoguv6TYsj7DLj5gzg
N6zE9SrOTo7EeS/IFbu+BfjPZI6KFKI+Xb8RvG38HNTjM02LyUdHrVjKXa/BZC+0
SaIxIAZubM2PsSc3XXgo0H7iBqm2E6peFrtInJSgVA+vA7IKjQWkdWhZhbnqrKzW
Nipw8wu92KVqB+j3fBQNm2q6oIdgwUzguGO12h+htfYUFVpnBpOLt/NwwSpkdtq5
QfC+p1T1u93q3BnKKmpPBumEpS09vjg/hC5yaO6ApxYDaNfZvA/rItNa2Xacwr+v
xqQHD41rap3eBq9Ehlj7HwE2Vb9YLnFLt8mzt4qtlAGVSHf/dhskr2scjiPVNQH6
T1qmTgtn510qj2nGaApRlniFmH8vHCTcUCo258WnHA77lhwXqueFSQneR243FYlF
VugMsyWl1ho9xensZi6jmjPwA2gXuBZXtELGNrKN1jEvgyZOQE4FUOo0QhA4d5Hz
y5NGFX9Gq075M+TRvkuk9d4RG+jnACCVw7w48JGMZdSSvGctoTHuvD1DA0Zhhbmb
XW1UyAZILLhDmbFt3MgbcA2Q+odzc85+GTFDfCASLd85c1BVCV2DJ+yZosO5yRXy
Qs753ouBMDXTANGyijJWoonxaI+x7TLxG7HbX0NksNA//qEqJlgW/OxKyAewAXnp
YXMn7dlaFi4fGvDJKqDokQz9OKKsWL+O01cbP+mKjg0Z2V7OvVXZJX9VI8JY3mWr
0STKYdpX/WSWaKDm0U5RJty3h2F4NInJsibucs7mDqLcO9ilPSa3KKUzcrlETJSF
ml2GksMhIrEq/gYHDyyklQcROp3o2gwbeZhVtmvYRUNbWFS9VI+b85m2cZn7A3qX
6YKl0aACZRc6CR6VRr6Y15SJmuX6gii8jX7M2bJ9xpZrKOIbU4EgbiyGfpLh+GCE
523FsN7JVXAdOFIMIUKkUinYwfWoYcB0bieA8R3f4P79qigHQ6GzqQVArGM7eRMu
zqneOq2C7INFbvAmKRRV2+j0ClvmL5Fztri4im3ONyfIGxEZ7wSVU0/bFryBs6Kf
LS0k660iCIG8vLRLmTJlaQA1xcoLiG6OhkEB3t+R9Z1WQcbBWlZxQW54MHG3YbUS
p4wkCD2M70DKPputMv/9akJ6ndtglCTqUe712uwul0xjpyCcmpE1cF5NvVK7w3EU
3eK6rQ4N1BfMZtSfc4LaDyl0EAbHarpKrEEze/0/Rauxss4tnE3D3dh6YHB0sAzy
ukWVbU7pAk0xnY6+6zHlKXtyDlKPnjQVHPr+9ExJpHaak1S8ArAFHWsxGPUh1DoZ
8NhfalaPmbHJaFYjmtHoVGDTRIHv+7vhMDmwL+Duk0hmRgKBFF49JJ5D9XI4GRuj
1HJgFB53QyPRAgwPPAfY1FqtYo2s95g+59ispx7FiUn6nKr6Y7YwMvS7+orBTO6s
m9dOUEO8SUpn/JF+wlZSHQEN+na1rjlpirPl8SxJD/tuOINC8seQBdmypwYeC5q9
ICdVaBO/6KoeN1nk8i9YmvPbpd6oxtUKAGMV1gdZSouSIDv5ylSJKn6dIFaCoO/u
j3AziRF4MLZI6X46lgb2S/aqnFwocQTApCkv1WnFLxBkjNsRmJFFaUfyVuUOU7/I
IgaE02FYaESooyGBRKbeq6VJ6mwVsUrwirMiO4tby0XAWLkN9mPLUsJLz3mizqyC
UfifXvewUzq04y3m6WH5grF2uJYS2hyxGfUzD/upc1E/0ZqJwAKwVLwMq+vwoj9/
PWwdCgLtVHeYAlGT+CDKsXkXRXOchknjjN9pzZhNxD6KusvvQrXEXfa+5tuEFXO5
kLQcI6LbVVULiEklyoOExVtQvuDtKOd8HeVt3ekqlH7eN0zJqt0urhIPy4S6cvOK
Q2TTynH94H263QrQy2v2OOQ8iqm68gRhJ4c1iaq9uPx8eNvhxTEeGQsM6u0aRVL7
i7Lbrlf6mLCHyQwLt14ofb72I9Tn8gzdk2LQlN8junxC3/iLsmQMoMjdpw10gKLD
LhAg0Bfdi67Y01+RXsk5Nc3TeqKXQPJw15U+RhEeZ5x1xZ8NskEaktaAdWjk8StD
V+2GKTcKhegWIH5KASPQwYWd3OxOer29ZIBWHYiGOeqVb98AGV8/ug+IcgUZpwu4
gydHgOmAnMEG2Yh3jC9F64n+/frKQfzWwswkPPyIGWCymXbtdHzr8uIk6qoHJgA9
7nXaYYKPW3znf01nW9OwRR1Q7B98Dl9nscSYvTZ7hIjg46nPtX50ZrRzywgumN7i
+WHCGkx5sBFhrYGQQdhEp4JUq/9qLLNXAnppmLNuHcLVu/6+R1Kz1gPMHrKIpPHz
tnI74eOKF31sXDk6fOuTXt1ay47W9JHdFOUu+4b3wge5HvnEFbr6gWhz6nN9oTmb
3k1YkRXskr6SWDBn0l130URpcZEnYtB5CBOXPm6Ntccinpo5R++rurb4gBLvrcr1
ZLLRag3XitTAILfayZJoyz6MVh4E696jGOvCXwOta6KGnmT5rGVjblPUned2/G6i
F2+eELhvSseTBU7sH7V2QJL16t4I5vjt9j60e/bOeeSLZKwbqf4ANT36ZTFzlwbM
uXzgHi1jDJMRZQ57E9phVd9dTMtu0bZLrcCU0lgIs+tDKqCBN+O8DxVphHmD9D8s
Rc5Yyi3MHblDimB95Zrzx3xbLIrO0nTDEo5rDMfSZ3RrxKSgR4n/2k+a/2mr01XR
9zbGVhurNtUoA0KCPUY5OSfbcsQeIpoTbP3VaSG3NG/ao06Gx19+oAYagIQgCcSx
NrzDzWZ3vg7HnILO+PHu2Sa/W2dqB4UyGCSiyz/Juv4F8LTCqA8uWaf3IAkNqS7h
kbL+gxqlBjGs9KG78WfJLlZ4LhmsQ2C85lP6vN2fkIrBnNW87EyWSgNN3yIeVWu1
Igo+VQOGCzqcjaPflVgUmS3/p99fR6yjgz1RAH0tGDnAKeNFpIeG8S96rNsl6BFq
WS2+5i6PzIEQ5+LGgpFxgH86GNaMqqtym88U5j1Jsgrq11VKvBxRyBnNx9kJT6Xo
G+tv+r2FrBNGkQ2wqwyEbMpWoKIDM6yX4sIoMPahU4HZcK9M5UXJhKABx1Dl/d0I
HApL732MwZiatq/4+AOKzJ/P+DDHmdPq7suaj1RD7/AHfVQ6JRQxJH1I2meDzRHQ
VehmC2FvDuyVetd7PtzwT/gipNIxGSJzFR6enayw4MJZDNL+B2lXTBj0x9UL2OoU
OIDyV+JROrokCcsq9+jQt8uGs+q19ugVWH45b1j/JAGtQj308IxZ8jhNfK4cgwRP
dbsa+A31XeiwQ1ZYPSLjd1Eg3gQccIfbdyaTFQ64F6oi/wkuFb7pVRtOJ9+wP3xt
LFEaDiF0jfylB8mOyYhHNOJ1yObjUrjQGgSuJM/gjqC6pSyeTqlf4A+izOAVuxUc
NgpWow8O0OECRAds0YGx2yaHRJIHNn1g1QhylBPeZC1WTL92o1AvTXGZZRMDihyP
DqowfeyIbCI1O2L8pkMwjB8c3f5RvfA27ztpy93LOU6CjidG8CniqBmVV9t37DEM
8bgIJK7dIJRYFwr0a451f9XwG9F3iEBoaXeF58JU0YraK2hrEFB77jnfiysBcBFS
rMDBmW/HkdDetJKjmHakmThqMR1ZYt0ZnEChOyUuQxxm/YwWSs7tfiJTNLfrcaWA
lWks34CVRa7j1DRXchLGx7ctR93Usdjp090Fheq0+u/k3xsyUrkFAekKCgmlAFY4
YLBMZUHaGJMi0qSKuPii7U8WqQvCQGtOLA+g5CS50/JuAFNvp74Mu1+9Do+esVs4
+pDbVDXbw9pvBKY5mkSBq7INTBFG5ud84aTpu4AEsXLz3+BP+gUcXsld7+C0h4x1
TQzHIOp908EJdZaED8ibvfV/4CP/c5YlO1q/wAGYraapQ/kS9O7lq1PNLKytUNHs
dmNNYr1K7BWDBRsdEFiDZkUiiu8/h2yKAQKm/LUISpXsAoLisqlQNeqgV9lMWgt5
TpD7DnYdkWKqI0EfCz+iuhIRIR4KvcbxNtc8wRRmHUyEvrLOjvYMxOtFliolo35z
Qm8fgndkw0J9I8CevARYP5uWTfkTbz/CW1wFDuZxojBztQdP3YrLuEZ5cYxYtHCP
I0ml2DgQmb0x0CpFXqgnDdNQjgYdAEnziF4gN8ui0+eup3KxeQ9bOxjRb9pff2Ay
rwCBY+Lp9OKyOvNW+p/FOEF+/FnB+hxZ3K/xlT6SoD0LMfPd5u8zkMdoTJLjee+Y
VrDlQ6umMQiuviXy77pXa4jZ3+6SceNfjvYZe8m68YNULzlHsZKxT5k0ENRNhc9R
Kxoz2HJ3r3npwiKae1xvXsJcA3xY82o1JP3SzbOfHj7RnIV4Ol0xfR2gv6htI9l6
7nOP5lkBN41Ys91LNSLPpiFq+kGZc2adE6/5CGRkzRkSNKRyFvkUUCGIEB1B2KL7
rapG9SY+rG/RSj7mtXfxwRt+OQQQM2JYtSrxZRsuAdxaD8ZyVpKFEqvmVJsi02cz
RSZSypDazir2K731tf/8T/cO26ZGWOm8rlCwL2crRfMiYSkzOctBplCh2kma2ilx
bTFqYFSR5VkTxwUYDZXXYgs1w7rqvTDdg0cBMMB4F1C6HmYAHvgUyvNDiD67VUHO
EZ1Q593anSi75UxkMRSMqPquOsBZ4/wPIkY52eg4d3NvIS8hOr13H48ijuJGkCUW
jDZGi9r1B+W/jZiprDWHCy1k7MnZV4HaS1TVXJbJ86baRHBpVHwAK5HUtEd2ntFS
grWhxtFTXn+0id1TsqKVfVfYJd1Zc56zAIQMiNMUvTkKrC2Go8euIGLQUpJjZexx
ULNHy62+fmzCmffVzYlPT6KQlb3l+4t6x3YahDQPCQEBlLwOfB3S6GpSxwYvRs3c
KGCEaPi7g7ezz7bxHmgWGX0B8r/LbCDLbhgP6MsehOJKFKfW+1PomkEhK9TSRwBD
EWqdDkaeZ3YLkKcX3COlqHBFQbEKsl16JIMm5803du0VTU8sLadJy9whFqjo9v45
oelzmYYUsDGcVNZEVyEz2bz5jDVMXJTf5C0S1Y5CzUFn8juDwJvyYHpyTEISkp4t
ld83IF3kvkmb58ocQUma/wj1fSHxiRl9O3JY2ZuEI4cSFNNWSMDTh9/Hzf/D6Jzx
mfbMak/HYHgcHVZCI/UV6ZsTcLWjwy6dlOB2gFmwyhCES3I6O744LPY9PUKSvUB8
7dgL7IyeVGitjCh2RtEchyCMtAgvpEZ9ZUY9gQ7BRVpW9f9tpLIxkSGwH8lhbv3z
oMq/Km1Xf7THQ3DmWZICeaMzk/FjLYtjcyRpzmPFgpVUEg9IUPRBsXhvVDz0pSwY
sQ/5f4ghaas8kmNfJbWngmclIYIefx8ACMIQzXi7DojBVmGunB0/4TFSzV49skn3
ZRiG4fl60SQ9LDcdxWFEaQlycAqucu6hzDRywNledQsPly0UK1vUl5iK0Fc6pE/Z
FqPRZKUURa84WyE1BsN9Vopzxy8kNthXeCB04NqIm7E3LPTdXSADWt4h64M4XT5c
x0pmBMUtmGnZn3iqeX9+AkSHDdxzQVWzaGijC3xGL61ENzARFFt1VsWRPTQYeVJl
1kTT4YlZ7waVogSw3ykPmxvc2BtapHOOoc/VjJHRLRmrDhssgFcb+NpbYTi2AWcR
cRlynUQBhAtGtGKaazlrY8cOXsVThv4ILiMs7FPeDOEWJhF/RsUPtvnEpyMZBmPa
tS/gLgrqSAaGcJAbRCMiPjn/YF1bAzzTwA8Z2O1+LCwYG+PbOt9GpHdWFzHKhHmf
06y8FhlFTlUPGdEGeS6MGTc08M8D46IwUeXLDp6+xkH7HVZ6kCx0dnXb/LLoVZCK
JtTDcwhLSwWhKA8UJNnOvFfmvBN0XzgyFoDl6H5s6Fmjs8ljZ/TsdVqv3aN0xR01
L8/PzySM43vUF+whqhdFTdeI9LpOTmNky4mOL7Y6IJdZBvkOStIFFpUrt6uYBIp7
3PNfZjALma7IPqO1QNQfpv24Wnkq48S9dcxYJjDJNxKOsBsgbjx92xjcQ5hxBJPU
CexCTPfHuHk/CBJABjx2UtTyeTt+lOgfjeWqcQeSfMyjhlX2jn9nWk1eYV0S4bx+
BOk02RzM0CfZ6HrqOJf4srXgImRXkOlVF/zPX8QWndR4Yay5c8JWRqK+4mh5tC+Q
vF3lTwyP1cZfmUyPIn7x694tlDi0+GSfBTebDhjwyYshowlawmK66cLSp82tWuIT
NGn1rSHhgCV8mXgPEhV0YXUtYOVAl5G0uvbaAT3pTDEzr2v1xC0K9GO67Y6Bc2ad
i32sLwhqSAIuLksReoG16QM2J+ADphHYZdaY8gEXVpi3eAG3VtkcUbhPRFJf+juc
uPXR22QDTtn+kLjTltcEqUPelM+9nqUpP61bzopP8r746/sP1F9hpu7KQK1STvwW
NoIF7fflDp/5bx5VOqPPdzTpWi40P5FydfY7/FgwZMoOt/gpzN3qRF/GbbY77Qvw
LfX8BWzHHSPvEBDn2vwefdRzqiMSIOR4wvO48LYmzy9PBKv0+w/8YUn4/2wuRp4F
MekizY+Yde0X4gmahtPV2Lzxw9sbLvf1fesBrl5bSLqcHq6nWrLBbdci6mOjVKTh
JA5VOuQqpvZxezI5xS0l416eklVq/rqiqoHweQb9GkBi4+mf/h1ABq6UqBJzLWba
/IyDude57htWXFNR2e4uwiVQz8prsXMTzA8VcdA1wbxnfQmnTgYoGDUgHkfBfK+y
wRUJ9P26YhmB2CgP0XoT18OoCyvID4qOYohz6kX9dM1eZ/GhGQuT7VW4uLyNK3FW
4MebSz/Xzq+XB/n8Cvo8orhC/P8z1k7tNiIgtl97Uuur+eCUHyNBfFns8VnF4BZ2
wT4+Bp891yH5xGH3YccuocndHD22IJNGnFWN6RhZMN74hsywqm1QKyYd/bSsGVyL
9/qIIitoK97edmOKQjwKXA6mDMYTQLAcEq8bKksfDmcWyqxNKYRzXQoaaPl1BwcQ
azympmdIuPgRJh1y1LOgTwjGm9SlJnhVEyT/77Is+eXZvDuVHIFk62zdp65ZhRtF
i9P2TsTzDa/n5IkVCtEeFFdI0D7CKM5aFf/SXBhlzrABYkG6Linj5usEbvNxACHZ
hYhwiZr1c5o9dwVU1HMpzJtpi47qPODU0fLG+b3rYmKNMHA1aftWri0UwhMnyQ0F
zrFjz+7cVb0K+6fHcoveVdVfgA7RbVbC4g7t7foIxF0HHzS5j43SoXcmRgBtk4Yx
OB1a4v5eF+VWupt7QtrqraIuH0pVQqLkybcnRHM06GJWI6aeaZ9NsE5iLYZKLbTS
Xuq0O+L3JTpAw7ppakcpUXvJDcUc2ACMIpigHYUdFkCqysqA2SmLadby3dqLPTeH
Bt7wJkVEM1TiKLR1nE1NFKSub+8DYhEM+DF1uOJPlWY4tmX1aGYYSJ1qQ5+Dczc4
tY40XkgWRk92N+gUEWqPe1QbIctqAHFr9rCyf0Hy9HBYV+g1MVTEsX3T0ntnRHGI
J+/qme6chrSJoccCE/kABT8E+cvkeVbGT2ORRzMEJbLex0sGsxqsGw3aSVGXnWdN
ErjNfPrKjVB8xUZw0iggv20fkjDoi6ETzW3iS6VTX5SKXoz9kxvYZV4rElRCJWgX
ceVJE9kl43g73AC+kPwLqmoP5hemRI4J4B3/VCJELUCW1yZ1LYAS9m3jd6uYIeuH
e68mDCVTGECDhzLFraJJAiIHpv0KJjdE3OqWS5O2sPqMLHZz5BWr5464uRgxvodR
bNZp2QrxDWmy2Q/DUUTsc9VqGIHt1LkxuHiA34GR2cBVgaByRAdBk91g/FFeZEkN
chOpaLcLb8csrJcAHFguciPTi/A8LsEmYrf9eQEf2w2SBUTEhVr2vJ632OUhYYwQ
3OGWSCVw48iZTLOIZx0Q2nzax9Vs+SvBZVjg8Ufl351IsnguPFHnH9eggza6w6iB
acilIZGgO3xgGANUASi6xv16eiVLoldaZi7cWBhfetF49R9urs2Eotz+SrJJOBjA
UgLZaMX7Zvw+qxUqYtGnCjjafj5IDCCS6IT4zXJtzO6NNt7MyMVymMioDoY3IfHX
eiOvbL1je+UQXrjEztAF4mXfrKBdt2mfONVyC9WXGhZmZ8d+WQQBWztxEZDjX4Ki
hgtg3ryn15rVWVMZ576A4fjSt+igRjKW7n/x1mX+TtvemZZkmbkTr3+yWJ/7pGjB
baDRe49ZJgtKaC20hMJqbDmryU0wb+Sm2ODIOEkC8r4s3UsY4l7O4ddt3wLagEdS
fWumkpKg/Q78SqttoiEQKEjYKG2OCL87xU++aHohcLroQt80iHhR37wGAXmuLFQo
obKB7vAOaQ3OOxS5Nv3Kl4xblYH3gyxErjy8jNFvESOr/Vxl++LzLXffRMrezgFZ
hUyhqoivGvkLtyAJYLrhAGU6uIEM9/MMz9e7qNIzMReI+3+sTE6b+eLSlWxsXbOD
BCkDMSjOBiOjtslfbjMojLkvgKKNGeVVgTq7GiCK3IFDWtdQgHlubqQ/5+/IDHOl
+oWK2l5a+XKbGc6YZPsyiwgAp2WaQiZPdoBlpwZzGqLt7oF8zRPjlbavqYZ+Dnpd
rMZNpeH18LXVQkHFGF+njoSxrQcNxTrVauUDVWi8MxLMoJtA7XqShCtx6uDpiQQy
+uUY7PZbWdRxtiVz6shwvKRJOVslrSC/Wc86u/lKU4KTjn4mGUxkNRwJo6rCJB0p
RClXIb0h8Wx4qgZZA2y+aA1qAU57xlJG6eiJwGnTrllVCDgTJ1wclh7U/Mgjzt4j
mGQnManaTb4vVjOSwVPL4rIe6+IPA/b66taddwUjucEQKexCxVedJ/pYdQeZHukB
E/vz72ehgOmzA001qaQ2DEHDn01caZoZarQqLpXQdgdIHiQRXj1In+MDUvxlQV0Z
3xWMbMNfJ/uO5yIlpwBpt3mQH1lmp2FvmB6RJZzPAC1FU3BzA6i5EdNW3xMn7wI0
obmXyG1MAXBNpMgXtSV1aEBA0VH8AsALhD5etu5HINVwKMfvLosWWbFRsMiD01ls
U9OAYA9aIYs6sL1CW7WRCyKl2ZYtOun/4nXQkzZ5LLP+zNCPWeCSR22GAyvquLaP
X2+KNxUedPEkxCK6CoOBZH2RF1n288bsupjqrrmN/nNIJAXAuQ+ndaqrMiRsc8yB
dQTyjAWqR7Q9hV2uSKG+lGnW8a4UBVOLhlLO8yHrmN/h5MK0xF+MWR+MTKKn42FO
f81zwkFRraJg9AFX3vqDZDnn9CKvyKJlskmASEkhoENNY1wFx5JpcmyvhWtcVZ/L
1PvBAlpmEDvc21DWdzk1nwMsiF++NCiUb2gMgvwvD0jI9+vtrH0Qdggth46G6skI
Mv7xMebauUyxNkh/AlrvKX/wM+Njfa7gXnantFLC2UuBoT523wE9DdtYKqS2o14L
Wel3IwLCcKAtnZ2C4hT43rETdfPmFqy00lkqe0Ezvz0kZK6A8FLWiBG4bDZBsNR/
5JFZRJcyQ8W51C0fC9sERNVPQLZvtuRjgxwOmSQoRzkZRM3GG9qZcUbh90F0JSdq
/Gtti1vahFOFJs1p27YKxNyoSMiYv51x/xUnsJCxIRD/9KUIYd8ECa8MS9p1Zbum
oIYU7OwnBxuxqM6sCmFEUl66o/A4yrpawwGDasCqHnOS8Qli38gp4PdtExgHM/Bs
gbbiu1lt7hu8JPdJZvbA4ExcGCbYj46aYYdILzsm4JuEMptcR83CdONpkWTLbZQP
v681Z0Q/i0qVzzPfCdRN8aSjHKsE3VafWEtFmuMIdhsZNIOqXoP8kwolxpLsLgpK
5KrWick2SyEeswnWWDAWt/lyML6sXm0kB6db8yYCTOWQb16bLP29tUyYWUf03zZ9
sdgQDpl+ZK4HcCsXB0tuMkoxmFUPsSdyXi6x4RpX54UaRXtphu5ab4JxfqaIYvSp
jzxrTu8NvMQ57P+HbvJMohzElyskizt810AQPNzAiYRG+iwxWvf5Wz95ZvtzNRRj
T3wLzym/k2/qL8O+ydbJv3zsVEGflpZk/lwFIhH2iJ94dhgxAvvOwKcG9g8wUYMy
I81BGJX1/N4nHUo7CN68LxqKoTiZHcojtItf7KPuL+U7BBlluJDfZm1z4MipjTID
8IGoyVNVDZ238rO6tA3HVbhbQ9HGMk1EM+bhPBmuMXeSSyg3ROevkse0uXkFSYIr
A9Xywuv+CuI9viiRdh6rTlHCPnpK7+19AxiU0k1SHtjFuPduaIH408NgQouylZ6P
1YMuIKPQ+6mcyRZNH62Qmj8VlQh7CwMLU2mcmClFrBWwUKkORY2HbI9mloB/AkjV
Tg2L0FvbS5zNt4/6/QpaQZajF5cKgkaLanQBYA0iZjtySboD1dwIHfxqcOxcF/jC
sgMXSc5FMeSTlzInB88UKdupoEDjZZFBt96HdJiRJRVlHo9UBOTZcsPlosvzpeNl
2gEC79sxdnCwDqK75awqfwL9l2vHdkL3/BK+Dg2fiBd4gcN/csoCXFZnBWscMYoF
yHfumR0FK8zGuostYx+ep7oQzf7/7iN+KleQlX8K/rM3Kt4mKoJz47dFqX5P3oK1
2yugoigU9CrOWpjst5Cd3UmdfazlTQ9wELelI7WpIkTW2QQFuyiLwnagrK/cWlNv
/nUAPaPcrrvwOyxpTb4Qe5VDRJXBhpY/pMIUjtFsmUc9BEFUgpKx1n5kFSfgZGVG
76894snmTtY1D6wUdX2WThaABmE+9Zg5NPKZHU1DwGiQFEmyO2MXUpOYqo1Wgipu
MCEtA0yu4yXB2pYWboacbPPtV406oXGiqkaCdvHK/TyC78MTs0mb2Jtiq67VTQiO
80tBk7t1w7YcY5d5QbFhDvZiScbwdZoitQ1Z0Khsu7mgA86J9HdczKa2bTYYMVQN
sCTPtzv+rmk8V2nOE3LmAcmpduBfL0KaIb6/nviPDSOwsEtyOtM+v+ZLgknNkjPI
nYKUvAtFfmiwtg/ftEU5vcY+UsYrjmQtmLOyIbfssxdZqGhqyUX5/3O9FBFfyCZn
XscH90CPIeRBxNZTioi0yvs1dlJ1jJuup3EDidH2uQeHxQ00kk6TY+/9t3/3+oJR
pAQEpbl8w3qSzKicDa8ka+rvQYXdh6BXO40Y4+QW1OEIV0cX4mw04yJ/NuUR9jUI
REKt+WnBQxFfDGpH1aNUVIFx2cz2iKHU26Cr+6geAYLdYASPcMe2NSlqRtIqyICw
aHTOwO2iFXGzIlC3MW2NZexLChBXoG/vhZ3d6YHhIipNaZ4VEmRtCD5K3cgyfzCC
ltfJiyK/DjIfTCxpbifsJy2Sbngh/mcg5OHgkNFrHhyLqY/Nqpsu1qgpij7BZgow
9LyPy67l9vsf8/DMvwj/53tThtQBOfroMuWZwPl9bFJ1QrrT+jX48Du3CDAjiv1Z
yshQowf+w3PhrHv3k0aoSHpf9IXYzjcnGlPb7kcCqgYx6LX2p6I5RV+KiGiZq05E
MU4LpvnCWXYMXQIgX8rEpUzQDPRmtR9Jz/tRju+BN/VoYpd79juNVkf+842yUW76
zV5u4LRIpPt+BRXOHQfBUitFUlQuS4WYc9WpN/y4inPA3AxE9Gkm1Ayf/qTZ0iyS
+MUXZW3dNKkCE60Na0+6qJQnvZhyEiNdbHQBVsXsyics9WHAQAxITRMN7Dmzper2
DeiS4tqwp6sAhHhLxG0S36pCnLB/E2jPPOlxq4mhXguUEJGj21Kwjcq2halDC2ty
cit7chEWDeAvir2y0GT/8v6xD+MFJkeNIC0HNQnRAPZT11UDW9R/CWi7OxX7AGWX
mRJUEZQqWS2M1uGVV40iZb7BeH4UOrysq5MGIZgtLSBH+sknZSBVx9ndqgum+Cjn
0I9w16cKbpdjas+lfFtqFy3gg4SG7DpTuiHbm0Vb7pDyjOXJ+eoaCb9hH0ko3NBR
0GJtes99qlK7d+E3ewxJJKbh9PhzywX72r7eRJV16+UwxPb9cKAc0/nL5C29TvhA
PexoN/4cD7QVse1C/kqzKD/qESUxHJU4eDKQyt9VhKuJt90F/0A+S9vEfdU270Q2
vyP1yy4kDPWszYAHYD2RW2NoL2Tkln2dGVfu/6oZAXHAiA3Br+sSDxZPjyrijywD
XYNIA/L7TBuoFKR8ctFKzHFjInRYROLuqAqy0T9ahjotdW3yj7tQW+AqBnFMD8pI
Dur8gbYmWPNa7xux05oV4AKn8SoEXcuGgdV63lVLfQM35kapcGawOxN+qwHvZmz6
5hnBMyNFzZ500EyAA/voxsj3JseZMWY24EndgEn1X5XZ/n+tLlPv5kWhLernutp0
YBJMf850r+CxkHgLO/nFk/yEolqaLIBKwS6gJzQ8a3ubYBrQTwzawg3OL73HfXQK
a584kzy3op8MkaD5lNjKj6BAyj1oX66VFn0C/VV/j2pIxteAzo6ixtZXAXGmS6M6
jmrFwl94wlCs2GN6cAiaZ8nqVdUhrEY+R3NsElAYINEnF7XkvsNHjYr6LCZYQ6dY
cG1nxTmHELjeQOW8lAVNZpX5UaPTRd/6ohW7+lFRq/Wp7im9pKovdap27PotTgkY
SpqdHG2ld1p5FPhhy+WZG0+nTJWeuKJLBC7ZC8eOpp9xyzTsjtQNZEcfukyMy7zm
bzw1IWeEw3+dqKqC6bamuvamqndSd8t7/PFJG055OwW4aRngazTLzJLrDz2oYyT7
tro/AxLJcrtoCePbXdxJ9EV+8w6S1il+bUPHjbztnfs+xydSMFOnVe+WO3LsGKtZ
aYdS11JYWtXXWkq6VXYZoeU+qIcpMcC1nzze3jePBMd48Q1AdqvYLfvcK1jnZds6
ys7XZLZZxKePCDrcjDx5KJwLdefco8nhyVVVAibYKW2IiI0g5Dnh8qG3SqhcgFSa
7j+LjhQArYrpaQ3j73yPpPCprkD/YBr7alLFpjJfmbMjF8lMIj2NebdcIL7XP6bK
sdEOL4QahDxZeonGboNE0kUr86Cz8+lZM2EPIRi9JYZ0W4twl2A+dopiWswvkLJI
f/550ScnaZNlrA0cAO8ZEdmyJ533RdxgiKpgJXsqkuYQLuW46+Wpz/InUR3qyCMB
Txkw5eogniKHleokFo/mQ5az59e/GbKgVoerpj4eYpLI7DqyMyWYDrCcUnXyv17r
Ew5e0NxzFLcuO+FjFkN5yJJuFGbvzd1cyQwsEuuU4z7XTESQTtInh4tF6yI/KCJ4
SOQlfP5iJHr4/1hbx5uq/B3nELbK9I6csFX/P5+uoCKPqylZg0w4DvN7FG1c9QrA
hksatbjtcR8FlLUtmiwM0hSzlk5CeWgAAkicIQQ5xhb8ayQ3mzrOlodb8NO4Nsdf
dZqwyC4mG38lbR3uA1NXcBQ4NAZHVuEKNGvKtA9BvbGGysUmE3swpWnTJr9pNY5T
Dgo6KKPiUs04VEb8lyHk4OkbpBwO+4dkcYd0t9qKfUkh5IWKoSSuzbu9hYa+yIy3
3eQ/yd34ECPjgDGwHSqDPODR3ek7SzJ86L+jqvTa95NsjVjY2MsKpscRzak6S+Nc
51EFmpN4iAPUf6m6JjiEQHzlFCakYArPOGI6M7I85ac9iY5FNnVui7DJDbGcP5IW
Eclmrw7sv8Pa99FJei3R9cj5Qa3RKk0ksRrWLSGjPRLedPwMunhSYAXDISLNPgJk
9ZzRp0f7bV/lyMGg4JdtDwzqHbqazP/ocTH8HHMFz+0LMZJgb8IGmglHNw39uYLz
bvnhoLoJo6InXZE8Qm++J8Z2HrP2Ti9msbduILDmhFgkHbfNWhaD6Gxjy+wb5ygh
1nwdXb08jpecLEwy04/a8oWz0Q9VLNCWeakGHIGcEYLl7gvMxFV9o8gFdm5vZc2+
NwBAoYZLy+jWUIVRnq06frzmE7yDasFLxKN0lXtSNupoOIbuYJv62I8clKHGFrOD
vh4JXgPBadNgWzbsWJ3p+If/yrHz99hbZUGw1hbEejh2Y3Kb7FWfHH8wbvHahcAQ
HtVrvtGaUuFBwcwjsnF2ODU3o19nyj/x45nlAtt9vNal8BXwxptQ2H7KoHKkoBqr
HfMGIYckR1VlqNQObdsP5qWxfVYS49eisc3SA3Fcd2PJRlNJFizaCLHHPvQz3tIv
xl/lypNeIyXaAs+GE/wkWylUQTVBKMP/4oZYUcOgELZwCkkqjHGwCKTY4WT/iULY
V5q7sR0jzI6fscHOMdy1ZVZiiOZfu7KtZEm1n/YnEH8flp3ISOaF7ECOOLrVFNbD
Lbb/jY3GSe+C265DCFat3czpyaRCj4lpjdBcGOPw1sCyukWXbpAKUQk146kntix6
1YLBvnLvZ3Ys8MOJ/b/PM3InqMUj8JClDkB+VHxtxjvwmEnKElJoa40WLbeuiw1R
INj/QnUPuDwoP+5vc2LK5FnzUMmJtdKyZdRcleyYzBwyg0ACqvCMBES5do19HiKb
6ClcTCd9S4zlBXSK9m/UG2DF4j+9hw6ohsUhN+G+ooqzCH7WjbisjkUHq7FkeSUk
l1C9VhmfBVaPoYhJRc72JPPv6S6Yg51DHO4y4otkYL+vhClNf0DuPQDc8q1Oc8Xb
CnfH/bv3nzyuFWUjpsAmuPcOkrjgtIJ/fpmPbe7ezvTjGUkRXHdgO5JownzgdyUM
ED9OQkCaTHdNMPTOvgu19RQgsEt61oA3HORY0lna6XrC2FCm2vNbXgepmdl+z7WU
VK93dfz+iS6wV/6X3wqFgvVPBctojvTWslQL/uEw/OseP7dMaNWRedbLOlFEVnD0
I6e3yDIjVgz+/woX5Gx+gyYtbvyQVz2mmf51ubMFG9NNfpLQHi3ZQk/FCh4niKfw
pAcF0oKTOLmIXtV2T3mmgHGiQF/wcGpllxbm6xZKVY6Yv/v4krHsak9PmAEevRCA
In96OYfDO5bsB1IF1kSjIPubqv/0vht9mnqrsykncJ5EwyXRzqqNerkGFfSMrkzj
DRcMxYfBsEvgaamMXSwAmbmdOa6i4mWd1r18YTKGExM7LVU64DobdGmuRqJT187R
xI5FtSUjdBU3ysXRwOpOUNknz+tUMxBGnchM/YFz01zHr8ItzbxK966nszTjDRW7
tPJDix7Hd1bwLgAIRyQ4P6Hp4Zr9/8oNbSV3CNjPU4gVu7f1Ou8u1CmYWWrVXksT
/GVu7D+R8gvDrsQFrCLgV24wlChK19jgecJ9ol7OmZUgYyLs3fRrZJYbtMKG91IE
deYRy1DYV7QWDOy51Z2a8EVwkI4beIhnWjFeJ8KYxrmmvzcI2xUIoXwN1eu8ZHoL
NFBfeW4ytoYT0IpRJv7eSD+kMZFrPpIztfwtMez2Ob/MEMPqEQd65LSkR9X02iqz
wguXhTrh3e91ASclu47C9PZSTQ8cxxvetTvOkuDST2hXMmp2xP+j5yxL0MZ888qM
8doXRu/xgopO5HpdKKPy8ehybOGOeThTW2cFzFkVnqVL64xw2d0MX9ECUrHtNV+r
6wTwxp3Q5TOUMqVrqmZaS8S4KpaNz4v8j2oxbUcEhInljKt5XcZDRnM/YyXl3giG
fUhZ1avH5a26ef7ctX0PYaLBvZtE6v1K1zsqroeEglMN8u71t0kFcgrAli8+YMky
/i5x62BbaF6n2wAr5+sYLdDyS7AwW/jXDpBLUN9IDEeWlc5hiFD1jv75q75XcwxH
ZRrBJpy6BmJBaFXLOIe738AMMDtbSUg2D6E9tj/O0NRLcu6/wWRIBVeVgY/OdChK
F2UFLj+OEdh8hjDS/oJPdTW3Wlg4CwaTmrJ9XTUVFEDOC03bBnvQc9f1vu+GrwXV
AKO6Wn7/osQIuwgnxf0SI7GfRt2c91Rst2vIot9fKqX/NNspLTSjtybPjq/vVgFy
BCNtaq1iXhQBRNst4dGajklzIktenb8pbZEy6MpDCKiC5c4EMhLStv7ME5mxPhiH
AcCpsFMVMik4l6mU5tmA+Tqy5IU3fNUTDMYWfzw96k4xY/mkWRs2fn0i2snuaEQi
lBfETdJuE2Tri/GKfGCQQ5FmlBIlZg5VHpHfqWDHT/jlX3gnFrjD7BRWln/cVmoE
nm3SRc8ldgtKVjaO1qxiiyAQRLX4bmhniBh5xecPNIvea5MQFy+SCAphrj87eDRW
0efdUeJZm9GZ7ZXopRmSdobcBSVx+0GsnGUpr9e6/DAFjDScR2whlCBGM/CE1B00
uW6N4V0fjRJbfnQSkBZNwotnLVw/2MKGR/NU1YeQiEwSfpXPDzGQHwm0TnOYnUgG
vSh9GXN9zSr+wJ9fiHhWJFRlMfI81nM7BGMl6vlsoT+V5aKS2WUm1zEel8u1ckp5
w/TfRiPkddFtzhrhMX7DIJemBJ2i946UdKno8OZmeJezDb4YCO+XRhEUnpR6DKEY
BT22AB/L4lIgK5cFQOhlBro9+6NeSyP3yN/FraCVkv1bdhQKFLeevZLbp/EgK6eN
Gu7vLYVCPo0NlpE2R+b9IQI8fioKlrdFqfEgGGRjWYNvGd2uiuB4yVkj3HD2YLpX
k18xFeaGPoW0WUJ+wBItbYMaNvoqlZKnTgTaqHZjANNeZKw14UtldPJaL4h9uqUQ
yevmag8GgdYzJS1MZDyBhvKTOF5+qh730gtEm/PD6aV7Oe8xqWIHEq8a9PuMGdzO
/gJyY5seLeZmHsk5jNWWPYZ+ZYlauQpSWkcyC4OvQR9CXC2GqgUkzWCyEcqd2G+X
qo1nnk8RhRfGO0W7VarypwTur4I9aYxXE1i2dTWKkKenfEx9KbD3FPt87K7i92sG
lGgK2sN9ZsxGbwBR1hzcHVPGmu9UYwy+9gfVz1QspihiqKEmmwjxMq4OpWF1oyRG
00yWZPSLTfFIKltCsgxRCBXvU4YLiw/g87tcWkK9GzZZBuj2MeiJ1DUB1x2fdetT
vrp5cWDZvkjKMXc5w67qjN9gTep6XTJgJ1RPQCFW4mcNUn0gCkfAGnY2y/FKlV2X
2fCwR04nWpnXezfnaY3t1shtKIv/s9CjYdRH4PTc269DXHjmvHrSQA+Sc9U1TwGz
akCb1icIVZRQjZEO+NAv2tHcwm7ZQDBBAV9XjEPzIVXWJJSfkOiRKx506azAi9RJ
q4K4Rh4hCz2DgBCK/dgPXY5/GI1UpR2LR2vj8H3ZFi1R8qioINMhmDYGpKNprSSR
kDNjL5L48KpG23fdGg2Maq7DObNZ3de2tzWn36/kqHi4lS1syvgXQyysJHHHixJZ
CPecbKoAUc226kcUOc7EQbgEWB+7IUr2+7lkWQlDYyXDIOXKKsWF7Bkv8r/d03Pj
lQ6rRD4iO4pafcJT9U0SaMkiX2sGKJvudoXutlvvaTC7AkYmGgA85++YnAlxc6S0
in05OIdg86066RN6Mgu0Ti8+o9ox0KiReFNW0jImi4kbdf/NfhLGD9wTkV/1YXrW
ny/6vLf8jeCKmGndeHxoZ5+uLtI298gBN9ThDn0RFD4fLuwoWwZab0bdAP5IOeBR
n7Fy+vkWclZ82TfCFcGMgvsvtY/EXQ5j7GUMv6/7Hv5aMO4uEDx7IjJWANWkZoBW
zZRl58GFqfTChuWlpuHdVk8ukfdK2Hd/uRDX++MaIRtC0FVvu5DvveWu7kUQi7u3
sEy4mjGfPPD7Ks/gte2ZHpQnNSPtm2KG9+NSv7utGb/IrIrjjBR8LwyU2oIAaMAF
oNKJkNbUm3Ok3hIQDVNbcF/6Kwxphal77zu8BTAH1hO8QU9wM39DssX/RtpJY2KH
JcKNSZ5fxMx6rM1f3AfOCQ2vpoTpJnB8CEyGPAaFo8nYZQOu70obmHFyEJGTFoQZ
ibY/26S8s6hT4Jy5P+IkS1FIWCkR0gKb7I53qFp170+4uB0429LPzov2QedSJ6oD
C3hIPbtCyepEIw0o4Id0cG002GID6jyUM6jNkHFsdGZHAgNEc1hu/iQwbLtRE1+F
AcGtyNQ5u1hnH1mAHBT9tHrJVO6/1h34ysHW6aOIpgfuBELh5xGwhrw0uPZ6eC3q
rBD3OdXfSoAM4ZcxuqysVF93szILACQSenvTDR8hp39pId3vol0TU4qxBvFTyuEU
H2HNdsNSkJ9ptiWv3oRn49aBNtJ9O7aqfjkP87UKk1P4HDU4IiLyaLDc8IRbxOyP
46F3kj/5RHmQBv8MjR8JYlbPb3NLkMsFvVxi0Jb1YPDxd04+Jc9PuiU+DRnGTmK6
wnNyRzsb3wU0cqg4NthNA0QYstCly2aEgEcTc0tiiClGac5ihA/6O4Zor+aOesW7
KjMsgfws6BExfrFDxgXfURIGPmjQBJB6DFx6ep8H32ZaoIZp1Vaw9RWMbJR6ZkMW
ttQWEP6+8HM9LYB5UgVaQqDctvNKOtVz0qX/4h9sNNQa+wJA7nH/AsCQdp0Xm9Vh
G1RDPpNEbG5ajFOZ30/8p9hdhZ7yQUXuwBwwlkvwT54TUZpq3tTUaXzuFBK11cST
cBNDLZpEypntGorHuEPBYYQwirYudMLyUCuE7d00pUB/2oOXjlH2fIuKjvPKqMZS
mvxmam2+pFMygeADL2SGV5WWYU4bXt/oG+wZ3wpsodwCKrT/q8dkvR7M4LmKOvtC
q01/JXjkiNQEsc8XrhuzoYqs25lrLvG1hD3hvfWy9XlPPn5osKf3MkvwqBdyonG1
IARMbSyyCCYiieCk9LHcG78AiRoc33Uy9UA91YTkLnLKUxvRItkYqo49jeJdNWX7
hUdxVNsf8EN8vQ2Vb0gDehTWAB5/QoYOAreUynpJ4MYuEfUTNMnPRadHyfkJklU4
gb/y0Qgo4yiIaEv9XVLoXi+QZdP76B9tsX96BTvUBY7JrEkdztRinu1fsKnLuqYM
D4+KMnGAIEZkyUctw2jOqJNbg1G9zWIgFoWhd/Ay0oTMRoJh+TkLrZ+p+aRZSP6v
A3X9ZFl7HfolJxKnWGUslmawogKogo5suZk2JOj/IwhtqQyJrr7vrwF4H8GZLK+V
jw3tUxclYU9TTeQ2p3qEQoilj/ojKR0oKSCYI+1owyxYYPRHkhIjDg8BnSDn4eXv
SSNkV4nDYGmCwZ7VjUoRGifS7ba0FVAnoa3nEGLBpLx4HjLOl9/s/ffAi6t9SduO
VATciSdlk3EXd8yKFvliaG8XO8wZWIet+75aDfjGOezHRCVQmDVCOEbBZIQmjz3g
V0M5YCJLqtjR/WePui62jBMAlPcck7x6ro7aSEVWAq2onjkh4k6PvPyuperd36tY
19RBsAZXLSTKfsFoLdxu+cdgJB0TOcTsElLJ90hRn1zo4Q2qHklCpw/vO9s0fnhd
vXK/RJpeS26BNNxcYKgqAQk8beqTvpRHUqqYboY+GX2/dWmM93mJXXLNSsqTCRnz
VP64gI2ZGhvDrP4MEZYCNN0KdaYe9XXTt4BVQKSQMKBlkcVCNU0/F/7s77hMog/n
JBvHCi6gfRWlunSpp30ON0ZJ2ok0TzVIsrQvSd31Fu//QuOW0HZm9hwqPSNtYxiv
LPNJmQDman9cS6+mDb5ICEUEPCu2QgKjnTWpzIdKunjtVQ2CwkARTJD8UKGIEJ6e
IpJjiUPQhq52pAR2NXLwlmYU5PkDOzkRYymFt119EfK/xVBdg76UPtgJVQw3goGn
XcyGzueKOmUuYsPCemieK54oYo3TK+8J0w5UBEFLQoPDjJLeJvuTzNA1kMrG/43/
eRV+apalPq2sPjr8PFa+2CR/yqbsVg6E8b8NUeRcocA1fBKIGZiamemgvHZ0hYzE
wxkJMtgl22bbQYE907OhpanqNyUwUpNSPzuMfUXGQE9hm6mNICSjcRYrFuGzgkAj
nOTaah+bm+j5p9BznX3TAaUWKWdnkczwaeKCnCm13O68ayfpNKYh1yoyQGzxuSqA
ULwUBiaVONymO3/viSPosLgwAFu1qhe1Nur8KSGo0DwrlylD6rl5xVBDp/nhXBls
D3vbEW7yMKoOJVRZLjQNyUz5SuEvA8IQ03gMnrRtgKRRSN+CaxTY5Wt0O+M9Emh4
FRlfQSO0a3XO9SvY2lysn8noUJc0HpSVHsrlXaewKHx87Swvo0iZvt5sYnmufFQ3
WXuKZVJnnQRfIGGr/rSFPZ33AD10/2l12FwtiN/CulX6uamfRyrIDIB+AA0iGt5D
Ub+2M/iXiUl3RvMqy84+87CA6EjfseSVxaCY0k6iwmXLckTT5yv7JxgZUUTuxYg8
F44q5SZWBDCmKQV3WNxN9nsWJgvlNqaFo+I4u+DU+LUUHfnIP+f5m0Qfa+J6pMYJ
k/HG/tvX+44LoadYbLWXFS0zPmFLGhFe7hJVLOhOHUguekCUaf/11qtpD2YxxCb7
bz8M5t+5gI2rdkUr7kqPhTFvV76w+dB/r6ETT0biBoTm+ljrjCpP0c049/rfJPuD
EIf1nWlYeXeOrtoXxiWC6igsfaEs0ba7Nz4qpzxsZeVitQbM0pxbLb9le4KNWdam
8bTXjHO6rc+/Ade7SkSQLXgka53NZoE5pyH+RVcwSp/smz891p0wuZBcgrJ+p7/f
aq33yS+fjzwgyRefW3uatLBtjQd0YnWYPP2iNCo0y96KDibehMI2baFHZkTarDZw
Ult6MIfHaNV15xs2jqoBLDUK56EVgAk/GuCswmij5AZufCZzcWqHP/Wsh8tzlWaw
EwUfY6UK7ioGhohmt2kRZwMlPUrLjl9X+XF8sHkY1U22UWm/BpPcFoMh2MOD1dBq
7Ua3tIoKp197GwdSYuawEURB2NVfnWRPm8E3rVtsn7esAI3NHa53rM0dwkNgHtnR
ROMCovbJvXyTnOpcNBS1xXTroKEH7CTIUxo6yckIErozc9Af9yTgbC1pgiQ9OKNw
Nnt+hPM3WxasnTrPVPkDQfMq4a6o8CMV6zLQMZ6Mz9yvUvVXLeEG/QcyvHWUVBDc
A/OOi4PMWuQ4JvEFdnDti0qXKfN+QNmWVoMRih2mg+xSBDw6GQ44y7lAU0TMe2j8
DsF+4N1b1zZ0YORr8KUvcT4b6aeKE2lfn6Ab47AE8RqNUWnN+dc1dY5mneSpkUxv
rZnqy9bo/5XTpAitQtIUbz7/DU+w20mU5aPCLGd/4G+ZprBGlrYNUcGN0HnoPJOb
9gj5yOhKNJoCus3IobkwWVS9ssn6PCaA1Kk+YY6yPZODDnGZNux/BXES4h9Yp5Eh
h4B8p1HPhX1ydXbZdIZuDyKBDB4s2O/mugj2d4KnRfGy9Scxr9otXtoS/O9Nr/3Z
D5Nbt/yq6RdrIhDy94Nu/BpYbB5BOVgZ4FUjR5ftuLnVoO4DN3Z+eEClKuf2lrUc
xbNmUuQ2TytDTqtX5Q+zo2CDaE+BPz7E/7uRNOS16dwD7+pL//S9K5vXpEqab5c+
sPQl7B7dHLEvd6W1KoRoIV1Z1T5ZOjhdDBQQk333n5g8d3SncLKGFyk8uri32J82
fBRgAmjT8WZhe0XJGo3atCYN5/P3EHS49CQD8U1W4Vy/E6tXtQWBr/ITztt9LPj3
k2KICUQ1b6jLJgOiGTYyeep+IHv02RmbwAz9okR8Ebk26sBDg3ftrN9Ws/BLLD09
fLEyn6KyTwa21d0Zmd+SbJ2fG5cnvLQ6ZQW2u2ThqZfswb6zOLYgdhyQYI7IEpG6
gLW6U4OD7+sk6JW9IDVyJxW2djr701HCLXbKeZ7kN6hZtArQRbejd2qjVlovW3ao
vf/sEWfoT7L0xnOtHUyv9SMWJErIeLNGW54aMFd/KX/0z+VLfyVEpQV7krY/zKuV
3KE8TC0c3sMbUVuj+GZ6A/JFFO604rqiFdGWKpFjaZq3ADMYEytKkSJFgYgaAJI6
2zsj4BjybZaDekVTjTnUCMTc1vDKH7cXX/DHVLoI6BrKxeo4CYDJSyjIMhLa6J/7
pSwAVOoXAqtn2Ear+cbsHGNN22qgA7qV6rYgR5PG5zlb5nhBw7JdvU1MWVOURzxr
Iw/zux5QaIriUoWokMFY4q9vAPmqMlBwfDzCdquaZybl+lGWr/G7qDvzdxuvR1Ro
uJS5UswGu30unkFZwu3UW2W68R1TAJeeb42sA+dx2aErd11x+N01kD3eBsyyIriz
rgViSDCGB6/iRyOiwF6RBAWUpA1Ewv1RIf9M8A70/IBbbHg2H0njsoigkGXwiHOO
3y07Ryo6dvGbn6UsD38SZ0jvHoVQGfBZ1eix5uY6Tmxl+PgAIkoNM7pb+/+92PbM
qbrppRWg5UJl4DzOjw9KcK/9G8/REyJVCbhdS9d+RisygRcc7AHxdeAztdNyKsZu
aUr9AJ+Stl8xpodGxdNR1uSUZ2ZiOFCw1VSYaQPtcG+2/cztqbEw+PPDIuZd1GU0
MOtNNtotUVK5RX98sHwsj9qo5NNdIqIFDAsXUWF4/AFWg6fe1H5OiFWKlEnPcaBc
pL5SJECHpw2BepZsp01a4y0y0q+lwXPLyOt9hOGFGgghYqRIG0OAdE0XGpFE5mgs
McuX9gQh+DUTJajUE5uyEmJsMBABCvFj+If1ONOeRwmBUiC5UARS/75UdWvaIUjl
oPrYoocVhINjIvmzr1mC1rKPUNluy1jbEkEsDsgIguwG5QwE6j/EdV8OG+zsx1AD
9JfOjr4rZVDzxCWtAycojcR2FAtEeqDqCzU/Re+QSSdgT7+yIaan9geGhRcRfDaP
7IaBSLe9H4mlkx8XCRpalgspKd5/6B/89v7qQ9duBZPHKDa+qkp3M9+Qa8UXB/zU
egETH1oD75JYS8Fi6Nd+JcCw9dORgLeC/Si5L+tCaZsP2sWUGKCfqJxiSd9Voj0+
iRxRX2qcZcgvZJVBBKTLmX6CUllievURCxSi3uzvKbyfk7Rwhn1p9tGfUZSmoukN
L8UMY/iXFrR6kgpHIPvlhzlTUBfS4X4SUGUvJclAUxEkw6CuH6vVXvlF/Upvhno9
EF9SViHPMSQqbiEqqGKNnj71XtQ4S8K1AHbDjXslmi+BHUpwPgMN6TK29E+fCdFZ
vm+NuHK+3y+IcWqEbwOiHnSaOH0cwXF2w9nMAq85n825i3NHCCjcgv5SJ1nHhpNW
hwQbOiYbDhyTuoQVgbq4UhN59BdVGVMHvQGgg9jky0qxhRcwNm7qkSJIngtBcgYg
56f8bZnNyS7F+sCEW43wUkIj7pggb/WYRVNRcznG09KOkTJX1/SdrWNwqGckl8VL
ZjKpbUiG/0KGNyHDkPxYRd/JqzXtd/OR9QxtN1R/DmmTJqA6sJsFFuj9EcbcGB6S
qIPGdt/y/RD2JTMeAf1jGZWwDKPEJaRfPrgXNrfBucphqMGThWqPCQbd9n+LLj5p
aavD3b2RMq15q7zq49GtQ7pd5QQGuuSFLKINUNyrzFy+jHjpQRPk9a04rfdwmftL
XSx/Kr/bpRjOrubp/ZqW/seBeMJM+NzFqraroYkVnK802j0lfomuUQOTIzQdc0Xk
2qtviuK+xNgNb0sYrWmf6XWb1cE2nUgGfWxpgxt2KsoGfiLvYq+Pi/PgjSMJTTHL
EZEpfrJ/mFzXgp2pOcKjIHzGUOj4g9UVW2qvXvV0NoX/tehqxWd8EmNEM3TuAdkL
X3HfrAKuKCYhOiHoYaRGAW/ovO9WQZdYC7wJMs7ItJKuHwxYuYII22f74mYFoVAK
bkVaQZfUVEcy7cs+2JtZDOn8RAkoR26qTfrsDBE8XX3ffEVKcu/Bs9ladyjMNh3o
gl0W+rYd2wy2y4iwSpHvzTWeWV9S0JpKapzE03IhuD/UzuOkYN++mF8HIFlNYKil
V8UJtgZDQ26n7EOAN2lW2sUMBKt13wld9seOWtfsPSDfHy4Qnk3EOflzUki8Kczt
Uy6jhEsiFijnk54GkWPtqFAgA4Srj8ph1pM8mUmCuTpsuXKFura7pbF0fwgYlCvZ
nEkaz1eZ40mFrtIPgyu+EuNK3/RBUL8L5lKPEaxzvlg+5ZrHbgSDq2BA4NkJoOD5
FklF5j2eSWhGQm9XlfAKGKAIOnUHW3FWrjKakc2huNeO4wKEU+AD4kynf1wYkhDW
J57+lR5nAZZu2fDt/bd6yeqJlSlowA6ofadgEnB+LlzIBREWIiUHrRZzSicTSLrh
vg4Ry/MZFJN2YzM2Z+SPCExoVcwUaLr009dPzpwaxjp5UwRRoHUiPZ0hP7t1qhNH
26iyzWqy86BUbvo789ChRXOqOCwS7083hkwUG6wnB1vZz0TXxngrKJ9W4r6ojKbL
SAeUr9IACLsnH5mK/9lEcz69AaLHzFGU849VX9Nc26bEQ/G6pVaNea8FYzF2y8rs
F/RVxYnRB/BeKlpfqIk1sfoVMzRQ3HFH/kXwYlKXlEdI95YDQFKSjHWHnk1AnCcl
5RQfm+n+MPKYi7CPEP9DUcBpUUEo2bcalKd5BV0ADMxW/Fivdp0OrGjncvieJvq0
9GXsepkQ972V7NcLwkIB1yNGBD0TUoDhfaQQnzAOsSxZVA3TamKtefewJnh2R4G8
YSemZMlZsGRwqR207xxK0IOm4uvQwXn4acKZLfeLvop9W9eM3gAZy/LjRoASVkpm
5og9B7z9+HX3q2qfbKDq1lHe9yNAFpaZqCfXeNKG2Q+K/pMtgegAAkIC5MYE0VEm
ji4jdLMlfDZwrX08rkbIy32By7an5iYeWiXRbG6IiP28Xjz9ttfcpBqE8wQGlUea
n+x5ap7eqDEdpty2tUkcrWKGs96farz0c7hUHUD7lrhmLMeknGISocE1hbZkM5Z9
DTg5a9tOmZUbsMQKpgT76vS03Zjgp9VonFQ7Lzc7ZL5L+PS7Y9olwjQyzHOVFcvc
faNz8jo68APVnogG8yOEKNu7PoGSYz3s4aiFQxEwwM9xePIVYicfEK8FEIkKrLaY
h+koHudnJ5FgpWgqn48BdG9CmEepcHP12liWoTT28RmHdhjyBaCjoV5VrXgmGem3
cTdrSN30uMyHYSDZHIJ9mWaYQZkA/BPQbJIJh9s9eIBhVWXSxtJEwChpPr5oiEcV
mSyw1ZqxpNEHQVfEDo3LUZygYPlXj4ed6mdnjJV+T73jojkrbh/zwasFx2XshBCO
dd+YClKqeaufMoKcZLa+V7B2OooBBZzQJCEiySFnNmybxSyCE5aKoYej3U5S/rGd
QP8yGkZ9PwobhICP6v3/X0Q/RbMpxBe2oHA4KUitLpUwRqtRNSaJsNb2VVvb7uFv
Z+s6tNxL0xXO27JiX33Hr9MUMTO3GLis4WaOUwceTjJFHyTNmtAv8qIkS95q/An3
7QaMAe7SWgL1gAwqt7V+1YXHM3ebnTADdhtUA3WnafiZg/jqvVmoYFOe7QhIasiQ
33acenWt0GKEGZE9iVdqW+bHbX822HNdRighqJQQ07d+Gs9o1KWO2CBCnxnHDI6R
cdKMl+qUzjA3rQ4fxXONioDkAsoRM+c44H1RTmTz8TYNUswjO5+lBifkAg+vtbu9
8t5wOF28xaXCU/gDFlO1pB/Rde/3fqOUihVGbXBAlfzQ0C7OyIqvaJ4xL1pxJWNC
2SuVsaIIqt+5s7t6ETljWx0s/WXy8Y/1RdDi6RasPIIl6Yf5TueLGTO4G7oW4hb1
/XsnVy02R+SpwUa9lJPa6kWK1X1DTXs+jnMV823pE8T+g0nLscybjS5ePF0HH6rL
0KqdbVC2gRiX71djueCnL/Xgb9e27ZY/8EVVEjDgeNEiJOkPEv7y+Ds9rc0DBtko
18EE3sC97shYg29J6a/1+ddL9ZaIwsY/Z5v+UQjwp92GXpGdID61ox/d4gpVBu/X
9cbtSw803WNxbQadotsWOnNx3dqrEBj5ZSeShKsbqXYLN1Q6Ei7qfkWeDzj525GG
anvy32Rn46NbYLGjmS3i4npbj0Zy85Hjr9yLzUQc2aN4nt/uApRH2vEjp3OySJsw
08AJPnDHUxLnuC+YGgOyRpGHGVXpp4UHW8xlOz2UhhAGzfQWji83LQawkyK7Vk76
v7N35Zowv63oPmB9C/ipNHOkxaXmo2GiiZvoaWmvkbGX5oS552NwY3OME2oNxXNj
Lvy8Fao/ZkwFa4h0P9YesDwcFgvCTGCOAd75yilRsBl6G1/9XH5VGAvTGcwhWhfy
nCeJOSuM4+aZDOdIYsV70zsrjfLIz1VT61Qhh3Yw+WoVhGz7gd1j+LMoFnrkEeHo
urT7t9cYjD1VNmNTe8kzGM2gwUKHcuSMHjhLItDtFlzvv91RH6QL3Woi7vZjaZsu
q5BiBvzN6tQE+SbEbYPVpPl33/cc22tndjbc3GzHxZhRB3SDYURCRCHnT9pRX1ZQ
2SJyLq4TXu0kvOr0JQLycpjQk94b8WasLpQQtPSIICW7IhHaFqEdrRw4ay8sMjy1
bl/hnmIDgIpXF/w/zenzaqME4eSK5ab5E0hVxX0jx2t07TXLqMywwjUygVsU1356
WCZdaIDkIlDXPEV1XClNuaM8/UmCqs4WDQPWSxbHjze1Xvs/Q0siz5WfJZ/pxpN8
SNbeyi4ILTVAmnl9X8Kz0YreMOHxT7SgX+zDFEXgAq4wwyh1fEOcW0ihJ9ZBcs6j
VRubps+Tfl4m+Gg+DUFwTW3ef0q5vRcAGaS7zYiGedmdeToXusygLPczeCX304GP
311BbwRi5pj2Tx71SEoxNi8RDbjAlxyfjb4LKrWOJKGiH1IEkvjjQ2QvSUzTXBNK
aU/9LBoPtPGVnUYakz3wfW1WE2ABy4rI6FNWMb8OgO53aLZubDLY2oIjoMiI5ZEW
3eK1QKatsDHgNS9A3EHOT0EWQrzDvD7b1x80k6GxbBnuF8H5gHn5BKhIZF59ub7F
3IVCBH44NcJ5dTWvp87aaMpz/FjyowX5O68puhoxeWkcgxzjFh6vUu41pcpg8bRy
TiIuZlSFZm712blz7CVbGkzeolCYwK8eUtpwtVuSuEqZTfTVyty+0XtbeqwAKQQl
16CVeaLxYUFCn0uMiNm/2VFdczFetZcU112/bKQZ+UovxDypHvE5ppvAt5VSaEHs
L4SbAzhyg4CK19HecKdmsb9zROajcZkIXXIbfEcblJVXs4By7vu0jH/C0phATNh3
WLuFoyjH22/VxipuPhGfXJvGeBa17kuWFcMCEbkF19M8ZjYU+IFrS/i8ly+Rybec
sOUnze6mi51G9+RVqhffOGAS8fYGwIcnYlHEhGNZRCsLvm3HosJlm6aEHfoShTnm
TDncqbODee+HA/3UMVl/dQYisN/i6o8VS3zJ6aM1IWU4Hkrd5r/h21TXP8s/Q4ad
Krw2bbhe3DL3Njnx/SoJWNoz8lA18Dmq4y6w2B8XBwjTDSoc0UgTeqq58GeczFLI
GVJooNl70Tv4KndV0q4veD6FVWMu8RtQdMBIWW1334G54pLP7Xx3sr6nqNnTwU0A
v+U6yw7Ef94tuy5HlcueWZLJfeltgIXutjNi2beOk+aVYb/YaDfmPomrCOll4Vwp
TMEIAWItlJqHxV0vDecSjwTdnYACcyGLTZ16VrbuXvJUh0E7XkJ4Xprx74C7hTy2
CBgbFP7rQcnKxu4KCabCL36q3MX7tKpYF3opvvM1q2c2kCY9F8VEzlB7gjd5R4If
oA5/APHaLuZfLsIfxrBg0isXdkKmegYk883OQuDs3L6szCSYKv7v3kr8aRGcecPk
aoX4SJi7MWjRjR+GLlq77GJE8+G2axvegTMUt4NBvlDiXC/TX5AOiK/+M27LISoT
Wa9D31OBiAJbxRTQCmXUGnonRZyC8G16/s0bCuNg0xwZB/EDHH0rHcxKjgCraWbw
Nt2Hn9XJpf2zdArL2gJruemdhVcApnTVo2UlgTLwOFfogBMEnCh+gSF65NLhwuOW
k8gG2Pp8PA3MKdro6q7pXwT+TlgmZmSurIePntiLPkNArmv0WLU04CeEczsA0hgY
Z3qrto2mUYLzgG99h/zPQZ9QPnfjCZiDBlrTfrFt1OEtSKvLt9mBtVr/Yglmiata
JNSG82rJv5DhM5ioWGAmW5HGqfLh/duHb21H4X1TJuAefWsIp1ExkaBv3rHIvafM
R94yXpuK4e0iBnx6KxRbJ1rpSL/lZoXJgK9QK+L4A6B7y/Bgq60ijSWscno2ZpKI
QyWA7W8eEnY2jGcb7VmtcqPtPeGxRXLPuXVxJWjEw/Q5YTfwMsrQxOfFwzHOaHf9
vzoVSGQDWmbQu5Xe68IJSzwVYhLDGt2TWXkw2c6wHvIoB/biAaXUR7Ifz5Uj/59X
n8aiYY/vrnB06Iw6v5iq41R2kse7her0Gt0ifcrKf8Z56CE9M/fNgH7aPmK5BSML
kwc5WU7kEes2B22o8vAO0GP9rkWNz8mf+bKdq3SyVkXNztaD15qR0mpQPeC9r6YT
4rL4wG9P4qy/g4673FNnIgPJuS/aaKFU2eNLchwu/QQf+pk8PZU6mw1HRldhmnWv
SyotxZGBFQbuJLScBYwtZJGrl6iN4s+fOu9FDKTfndjPNVNZYqpfkJJLHle/dOHp
ectDWBa9gjglhgKtE7EKs/F6iBa+6oJ9NPvaiPugwGr6V0wKp9kb4cV+cex5WLD1
vb4hjPDnOIygiNUprkjEJ0XgYnJyYB3X5ZLa5JHiJ9qvojLf7mxro/R07GU7dGNN
W6KnI8E7+lRtn2d1YklP8BX2pxWkfzfq6OW6n9gHWF/V4IrblVIHIkPfOXJV2Zw8
+ynXtjCJe9bYC+zlsXyRteoN22kYRvjKKoYpsGTpuKtAgs6GfDROQOwy8qTuY0aM
4FVbY8lRhiZdK/e+wvKh+kBbQGiuGrvnur04vYUYfIibJ9aTBGhCdvAxARBdfBy2
VNgWjZxWhIsAxNPYTQ7Vbmq78IHQsJyk4+wddsW/1vp1nqaWnGbq/GbkAczQTco3
gz+kWHeZ5A66QzBMbdq0hVMoDN/JDTeeXDRZl79hSex6VBDghzdMsuNQx/auaQEG
yOhrFouunpdJDUTTm76riiJiOV5gsRrrb9m+faxLvfp9+wKb/p3rkW9oH6nDYhZG
k/FHdzFIX3Ar/Uqw3S6CcJzaiRmH1ZAO6pzNSM6TlAmrzfS0Up/f+BKXKDuh1Wn5
l4hlBWhkudGap9wq3Gd6X1R4h6q6oOeFYV1DxtEHl0RKP1jt1RNk2rZveESVydro
ztnJGQaMWQJQKmXncPJEdL3mtBZYgkOL1DGp/lB1dlHavGqZJaSh3B0hUqQuqLYo
N0S2abYeGEVoyjPwvij+Raynmz53ffLLoo8d2VN+27v6ClauDo+aMXOAm2nIiMvD
i8+EExPobYuuYAd3KNnbc+kIRwCQ4BC81hkmcvy1dOAoKMfDBO9HPEx+d2Z5ZBjZ
mZ4b3t2A2bGHevzKXnmNm2f5ZlmdE6o7cGWvR1IhytmRSxEfAGI9MW86CgLYcetr
Agx8gcMqds1qCWpXCUnK0y4xowBxtC3kQsgV6txeFHiP+5iMqOYggTn9bQ0dmvLp
BgIQzPGrEqIy5FjsBl1FLHOcXAwMBFgHSWp3UpNTmFtJMlRGpB/6YO0L1A8lAxqy
Hyf19yX3/xUMdDysLPxsktBfQZD7gCtpcOzcTLzYcv2QL2Elsb2ccp6x9rY9ckMD
b+G4jseg95as4iL4t/6/p6M6yU+sj5JwhfaWZ7MZuOPDTNTfyE2Zw3d9SrucMgQ1
/afqL84Fd6JMxywYhV2srw4uavMSzZsd2SwPT9HP7WBzTIdruvUqQTND23ummS7C
HPs9kCQmoxbpbfwcZsjUYkUqOkQ3nk52lRShYsl7onZZtKBf/gfwJwEHxkEXjzqV
aNKVa4erytuSO/B0FPwM6Tw3mE1tV6umVPP66zXtMIIOgSH7ddnM/dte2kcjcqQ6
5rpvnNomukBdb2Iu0LZXaCAkhv2lAbiDHJGZBruXmemJCHZ6DNrzia3QsroRM8Qh
F2adiO5FwItCggkiEyYXeaFnrhEVNcuJVsAboPugUgV1h5ZeEcfOCPnLZD8rbWWt
PZh5R3LVQXJJQ42O1+XXBpDx8WNPsez2SkRAlZTlTm6kgqYWkvTKdsU+n4O9ixgP
SPUKEZ5eMUOcc029KXzgtIQVysKaiE8uRhIgAdHvDAL/k/zY0QilIzkIvF9uWMs7
u8Tkzb/paosQJS9gWhmAwSvZGRFaFOfPljC+0S3G4qP3LZlEf8UpP49waZjeofyo
ytBkCYfnPp1wlKOPHcFZrR3urA1Bs0NLgHnvnbr5aGbrSn9cFH1bnTosMhdEq7K4
tUfQuKL4CFRqq2vOyISydpoU+FYZYeJtrAX28haE5RRdfI4KEldDNq9KEEcp2L1y
AmgF4rL0iz+r6nVJJ9Dy9LLrKb6JUnDrYXgJN/GJ209N4mcwhubt4ifYaxGgEy0A
IjCKE/okHXH4+eELPQM2DDSmoD9SsddBTrPa4MHxIjWM05A3BOl53+wM+gAEDWea
/s1jBpWwrbCrXBiBYqY2lxkOxh80eCNdJ49fXyEoI/s0P5tuY9An+x1J/JPA16Bn
PIzPKBLvqsJUFndzhXbt7AJAhLeSt8aLH6CdEkBcgH4XHuLoWgdZCK1bN5WcgkaN
9FLsHSZXjAPxxV2VI48AqPm9ylEp71MbhQnEqVNn84y90AaFDHacsueEEIqBqVi+
TWaTigI2QZJexOis9OwGsIP+XwuVI9lYmz56ZB/ulmrhZ7s8XokD6H/ZQArBLTlR
oJriTtolrsLAtFv7zuf7x2i8g0IRB5dR4Ac46gL3MEr0lurGFttWER7zWV2IGYi7
Hb1A8l5m1pih+uQK4yXoetBLTHxD2XGH59iPRj5JEV0b4ktQhIQgKEOHeLhD26lZ
vD3jjFxDvv07zU8MwYKWGGad8JjZOJKXr4qEDm5K3R+tzqjQu4SeOJ4wYu9AIFD8
5bOuZLGX89ZVlQXcc+04Yo3VVCv/Ox4quNEYVzb+27/pMxU+8eI6w8ZluDPR7Hv8
WCunubNhXP6yEkbfYvHrMQNqs37yy7Erz2tl9LdG5oxuQSvmKxazfYeT7ttV79um
xT426JieRbZ6OossdEZetYl7TY17HdTJZBgxZZ6e1gK5uncm5wPuZceBvNw/jn33
f6bA2RytRcoV4AagqhLma4QtfxpLB8hwX7ggn1seOVizvRBzjUtRhF/94MfJ6M20
0f3SvcB0gcmUAqz2hX2mrQdJ+q9SQZ91kCm8AyzLxhW1S+f1jmFT/422OH+e6ppf
Tz98tn3AlqDPI9LWdQVdGml1OscRH4wc03FDqAuLR+PXwE0PTLMNB2ymavMCGkyh
uNRSPOX0u9x0hBXrBKo0Ts7NnPD3XdY9A4KUOGjNNSHH6LSt96pl98pXR2K0wNpN
iXV8uwYZ1dIB546MsKOAKhFPFVHSwguu769yJt4W2EPICSTNKv8Xl558fkEz/8fR
85gOvYIPrNV3Yzqp0l7D8ul4v6jB7WgiJ2+kM7TpRo9alYccl92KOV/sQLR2Zvs+
ij2bsCnstJRi3REUZgBbJ6H6XjXoJt+cNEMp6vV8o+ZfACwfUb9OWAfg85tNUo2B
uAaGF+eSel9wpzVNe0m0+LHgvolaqq3zDGZ/beLiuL6LbNqvQEo3OXn6ddqvW3g8
0USMoVJOJ8F38Ioi+lBdYjA8NCfooEiJCK6srEy1xrQI1r9Js65DZ7q0zDkICiUh
OpUSqc7ncgRZKUwq79w5cBMrWkriNDa9r8F8cZaMDhPTV7bt7wJa6JrtpQ01qwb/
UesrPQEd5R5PoQk302HQJ5Es1kWY+/KtzsdOK/QijENcEQHdUQ8XJ2b/BR43cMVL
uB17ztMQ7S89EiOQKNn9uTlao4dyEG0RT+UEANkC5LdhrkLMeaVKMaTOQOpOQoI3
AeUYU8R+Tc0XVEcs2lgstDBodBZelCAiMdD81is6ykfQdaU0mdlGy+r0Mx1IXvnD
puCPQ6l461QXSOPyQAOUzKw4KY2K+Aoa3qDuTlDyNf6sHbcyCb7757co4ESs2KUE
MHQrFYzf3077EPsN93VBeB3KffwyVzX4vZdLJZ6W5Lr2WYSQ5piVysTy2jMQQCKR
G5T1BRyw4+v4m3lSxlDFKLOH5umDO+sUpKlbQnJTI47It1v2ldAtxmWGueqz1j3X
7dBfpIzGJ0EEbVdyQQPiiwUPnUM92ac59VdB5pL2+h/+N33llDby+b8kbFP/yeH+
s1zN8S0Dn1n0+LTZkm4b6TK4y6YtgS0crSyMnnQKZZx4k4a8Gi2hCxR9Ab1fMNjx
l8PfFZf1OvpTZwlAyrXe4V9n/pik86fSAi5CITOjkf2mQQDy3i2mugG2qXyuSRgc
S/ARFQx77iopY+bSxdXrs86rtJRHLLorNOiAChu6Q+ZsAIFznJQmkg/WkTf7u8RY
lc2iJ8A2CJxPQwpfloUhbJEiVKiug/giT66aX5+yRHwvH5AfleQ4NHV86u1JuTlW
mF5e0JeEZOExYyM5LF3+MIsZXBYw6e4+Z6st6bLHBwxZ3Iwygorn92jF0FQBUHWU
kSwTc7G8oXp6RymuwJ3a4+5hWRN1a8y7L1lmvJWetWAfSgZCRLuzWcyVzrhBH30f
igR116FJNVedx7hISasE3nG5IZc3qfQVj4x4aLoPouPb2FXfvvyEaND8C1SeWWaV
sWeGPrSBIdSrdV9XW6Jc3FRa//qz+6FDqiTBmxHRtqkSQ0XtaqtY3OwThekxRyJl
xu40VVm4pkP9WJWbi522BfLtWhyRjvg5eSIFQlPblEvQiHmbRqM0p48SmtiWB2Y0
hpm430Bjb0W0HUQqF0moohKxAwuok2GkOnmnXIOOBWduWuDNdtsoYPM7RNDUk5+R
gVcgxIMOBYY6mvPBycUqvf8v5tV+SXO0BdOl+BhfC+QEYcy/tmsdh5Kg3vFh5IRE
5/ax2ZrtUqtCrt9eExkGdLv/Q5hT7W4BzJbPyC+IEMWrZFhusK3EdHrmUtDPLbSE
PE6fq3V9QOKEOq1CWqMziSsyRxoMwNP+y8j5fb8bpfczcqcL/othQVfL5/Zk48SZ
Zr7NpdGo6xql2oFLhd3hXuHZJIiljhuCHky93fHpcMi0Ry+A6LmYdAuW+i+tgOV+
TRu6gcKGUi9q77of/mX3fLf2EZG7BHoLkwYW/OadmKanXRwRGCxlhvk/C/NAgJQb
hwv4XAoSK384BRivL+nncJ+b2FLnQuqDVpJMSHUZObI4gaKC1Nm95d2k+ly50eFJ
nDclBNkJOEacQUmjTMoALBVZoS9rtCC2Cp2qBolM8gfEMzz4KEQszJJSH9TQEt16
IBySWRHbpQ6sLlZfa/RFK0ZFgGBYn6wuA/X/it0618PkfSA7IOpjue29CiIvcXii
sufinvYaselJXcy1gCJVfXmZx0eH5CG8owa4/b+h4bWBXUy0Z22cMpyPOZ/23eHX
B3nrqHl3STkK5sHrxCvTc4dgXnHrDDnRy9MpPJYnXUCmJfEa4NdMns4PXutvvOj9
vb2yUZNXtmBUyqGiK1Br/qdhcS/jaCjboH/UQm8OFCDzRMD2/TLjl0ytcX+DUpb5
xRDSKQBBviDYuNgHiJCdsm0mhJhTdNETUQ6LpOhTKqKh7skrhU4xqEAURnf9UQNW
ynABi1KY06QoHvaMX12w2uykwDsk2Edi8X8XJYFxy0ZuFeBnBtnkgAHkjqs6eA4O
JEnbyGgg/V6r1Qmr+5d3lVGhExAiMNy6evjPAZ5SXqppvVJK+c5ulPZiPG4rqa4y
OwPbYxgsX4K5jHQCrMQa+Scfi+nqV3XA9i5d8LKMO3TJw+FRQukHCRVDgL17bsSd
8vudfKtndNRz/TzeDlvJVUM3Irpu+WawoDw6KH+8M5wPnMC/L6iczUM3/ZgEtdO1
myHmjEz94oxGseZ70OQQk7tkYHQXvRIj1OLle0Gvuho7l81EM32lylIPR6xXJc9V
EzbP0KfeWY7VkHh9fljQHh5n0AUAC4+Q1JORZJi7Pjle5BoqqksjV2RbxWNsbDcK
FqgXh82wKIE9peMrU9dZmbFSiyEX7APOE858olZxGIvKC5bpfxYcHy8N30iraIHb
Yf5vk7PXEdvwGlZOdgTeJwcqQaFChFDslg1eDNSbDZKu7K7zfH9fJ0fvyX2u2m34
bPZOxY+oT+jYSca1FjSU4dQilEg+B+HawOHJvFqtEDZTETEO0fMo0XZQ7sbLR0RL
D+0v4W5NOuos0DLpsOgLaQO+g8yLNMPA+KANA7v2CEsXYSxuppQ/njRO6Wimmzs7
MmbMyZ2RlWRDJlDAdO97Ub85b2svCQku5Te5vhhANQHYgcVyJgkOnMdX/z+KylDu
B2o6vFfUxi/H5NpRdcZN+yv87I2W7d5TmwlTyM1k+5fe0Vu06W8i2catfcspuRY7
XQrg+h4wITCgbd+deKNfgyjByxIdVcgThYgTvFrNmmWaIxoligGgz9aI8rfNtUtl
St2xuq7ktximt3XMNeQ+mLs7ANrQPE+dSc8kb27Fz2cyiUYmXvpO0Ox79PWsKx+m
K2/vebYsn6hT+ArGLBWaFLvOg7AvB6moLf08YJsTAxabtwBOaZOt7ahB1NCNlngc
7xS9AzrR6XJzqJ4VUD96CQi3yawVGT5/PYtEQfy0SXTH2itZtwsz4E9j6R6G5AK4
XgRsE4TJcRGSqzf/7OPFFMtCXCPsXEEvGf3MIecyGDgmf2tHnbwHtKoSp5W5HnZA
j6ObMZ80RAQdEnm8bqTwJgdOR6YXttC1lm1zm+fNZhCsMjU2ZqRSRL4L4J1zd0Lz
VLmePJyWlQDM2XPJ2YUsU0Sv5SesJkVXH4B6B2VzXmJrOfdCAI3KYVnRy0dzyzeS
vVZ5qYkvbJxX2MrnaeBNqUkNyxJ+dE4/O/r4RlFSxo3pihvvf8NpVnA8A8HovCGS
lvRThy80OHYHPxR72OJI1eOuBGcBlYYmXgG/yZ2pUULhcB6mb/E9Knk6bRV3HY1K
jNYLRiCLwDeAeyaSiaNOX/r8J79aDSJyQzUXQpekh3CAIXTl6NOncjOpVdxN9eWj
Ap8jwFMMcqA8zE6oqzNAeZ6eOIlWlVjmDJsSmMC3/FgHUyb0+kka5RxyKZ+nApZH
7oKBfyz7cfGqc3NlhibaqZJ2Xz2BRgbjJYiJEmKcG7CzkRQrJBuN3NC60MfV/408
x9KDYLTfN+KpJVxRWu6bC1EmK3R1Of70Vt/zBzOu+GVZ/LmbJ0mYoyZOrgrWTaCg
8+0xX6lbRtJdXqnN5nf9oVzSrFXMLrN9+wpXdN88EE4ZaVUWuccfiA0Aa3LHpJKJ
q5DWbRZz36jgsu+ovieTO9TafO4PMkOoOETXWWP+/wUgYaIly9sArUhClNVtHDMN
L4vJksi4BbQP4vQgw9NMMJCihS0zztljKJU663m4+mR3U5F9RZjfc4Zsc+wVo1hN
pgKxkbiw6caaCkBeJntpzhocv3pzKP9egbSB8awbMKRdXVoCFAj6hWWcUXqxcomT
kn8LWiaCH+6C/H3ONAZ0m9OKzufn0/ety02SC6T0+He2WnkNs1b61bhC1yt4pgfp
vtDYzq+J05b1CeEItbFY0FMWUzFv28BvV/HazsrsWDG7YtAwkx4IrOa3BKLdFgWU
nlbmnTvecPfjp+udgrwl0lG+1v5u7un0dcTEZdx1qYGASfkdEe4ty5SX4QFMuDFI
PxN8i0J9sOSFh8E/hVrw6kK2MwfqbM23Yln/eiGetkWK1XO27mbvj2f7w/QgkBGI
71TpT1qyY8riVaXg6HOCk++grJDO/7QXfyAqzeKpCUaun82MdC/v2j1eXfjQX7H1
e34f1ENTTGlmke51v/iqL+pPG74IRqORsomgHaq6ZX2kvQrDn5XZIO5PFG26tyGK
m5h6BGwdoHANXlDiZFvbR7uD3aCmQEErXL6VoBDX3soWU8AXSPvPTzDX6IOVSV7m
XfGejQvssyO09FFa+aItvl5g+V/4KbnP5dIBiLfwy53/cBKsmj15aXhGaRVX0iWQ
027rBZb+6/Y9qsQmRmPZa9d+ItubR8FKL/Z+MxpmV/oY7+cXDa8rxEdFsNk3IH8x
6KsgzQQj6wtu8mLdnSe5Etn/kr4lp2IO941IBKuq7id50S5RwinMFOiJm3CSHaaX
D0h+drWUoQNe7e8vVQEIifWHBYjIZSdXrT1kuqC2mDtLhE7vEGNtV/nxtHJ/tRp6
O7Pn7hye36nauQTyOj28FHFXrw+JgG3/w2CAw+JVb0rAr2oVHDj2qrUkal3OPOC+
2VwtNFP68sFHTSwjSZT49wyDQqFMc6pFukQNavRKe7vQTKbx5xFSgGkvomtrtYi6
eg+hA4K4PYcsQG76fQPWovn5v/YLf/mBupwc1/NMqv2oYjgEh0n78rJh/uNBlFs/
CqWENGEcWTHRq7j4aNGMFcdbMpPEIyC6NY2s++i11RBaoEiEfvrPdNpVbqem7rBk
74rLMPjZzv0D67/y/QxFvss5irOrXBLB4ft3iJYK7AKhBbQKF4WigX4P8kdcVj1c
O3HTw5Up2rM7rMmN/hZqx0yR7borTOJql88Sf/ysSJIZyqBdPhKcnwsL3OTKdu53
bgpcE8FjUG0AV5QOCpI1xJCluNcDQ+KRXHynfOKXOHVx7B4faU/tDMKag4bAb274
tFXPP2XN2Ppm3KcRYP9gPriLjIF5LsJb1ZVCuFO57NcQxfogcPfS1MLuqJXvD8md
WeNs1hblaTjMOo/jLsEK4uiVw0v1B8FzBPzVjvXlVcRDDmmA9WxqcfjXYiqkW6te
J7KFCv6f9hNLAEKm/FgLVfT+zhZZHMqzf7mkc0cQA15HCGVAd2J/oVcgVGReikH5
kqvG0iJg0+VvcpW+D9o5PQLJf62v54tHPhKvAxq+bTKT7skT8WppEHNr/hqq0vjb
ksKwDgxnm9XxoZmGkaDUBc+2lbj2ptDXwPeNexsHTZ8biBIkW6lfHzvqpJEMlZOI
0DEDGdkvaF8Yipom/cJetILj1GK+4ervrHL83r6svedXAhvH8FAtypGNfbLUVY0p
RMYykjvtu9gQTwZetCCJZAAThv3+Saewu8uQTMTpsdvjc+q3bQKVAz5vwOQMzRn+
5yP5V96LVKGH4uv4qO8iXZH9O1GDMxreTe+fRthZ/0CiuL0WcJBoJOGzAWzw7eUv
HuI0wedTXFQaYtyzjAQf19BCeTGLiyBHlHseMfXvlbR/Nilxdu/k9/EgsMIb+C87
7jfAUnwc8UUU4JYSifgXPtBOUiPOfwQsSUQoF7fsXlcO0uMUIZLkdZUYo8Y8qwqd
tM2IJl62vbxJqXPP8LSFgrbJX5IaREx9Hb8tuZzRBkNvwNYCU7d7Q3SiICSY4E0M
z/vRSVRBuKLJwYPWU2hpFmzJfCGCIRvXBz8jPs61jeNsOhqcq4eQtfuwXrJktNj4
pcnGsb2SjdpjdmQXj4OacIoYhHiZy02xBzAokofloI/pj32ZjanVAECSgW6ONoRS
Wx8ueJ5gfmhVjOlJ97YjO1fkFfE3r6T743WpmyNOlZ+J0/+jUgTA08RdyMUeiH6j
Yy+LAKF+R8WgkW73xbjnS8wHyFUS2X79A81N/9u2w/mFAirk+Z8bpeLRb2MuqgMS
hMOKyWaFksFSH00IKhnMbynrBa2O+V+oUJb2GtoV8YLt+C+U+3U0OvIp+d+sQCd8
/tkvniu5j6THU/uXLQ0Y8deiRsjh7RMgEOr5vfIdaexesHc3kXBEF2F5WbiHS2k1
u1L0R3otdRaqDKS9rmE0RZ2DUo5bWtTdHd+jxrfqu8Cs2pZ9mS+Oy1KBmZR98Fkj
fWRjyhF/iTJm3Z3yyXPknJBg+TwW/6F4m7fzVvtfEGw+Neo1qEUuVjiUF6XXhnWB
n8Oe7qNTskqeH7YDP4nZVOHWtQETNBpVDIyvTBtrpI4gDldFy+oPf2xlKXB38lgh
1VGl4e3AlzP1qIB07OqSAiW27jQk3Qft/J09gPG00knhTQpHR3Mr1z9nfidiBzss
qatpe2snXuZdPF2GGYNvmmN/v/SuudxXWYhbHF+Og705G2/NxejqVL5eZMpvBRgB
LmRH6c5a4UOqFub/LAfPhVswEmZ8GYW3n2bXajUCWJjZ8OI5tmUEzB4Lekg1925t
TnrgmLssYLLXZaABfNiCwBYDD2pDY5C33MLf3r6GS8ZkdMNav0sQDDSBmWeim5r2
X7uXdIgHqB0N3n+wTyWGCNK+zw9VKetIqMx0frKjhAFTLgGWbmLZgynht1KtkXpP
KkTtbm4qY6sXvZI54zh8FqeSOrdzb3+FXRKfl0LPaA/TMG5pNC2U6gZauifwRIKH
59TSkDQoj7LRRUbBFHk9CY2IlB+c1lbmxNEB+oRWEHKgDrhMBUOZQZTy7Khwuf8V
XITG3BkFi8pCsn2QfYq23eYOZUz7jdEFeSJhWe3HoY2WNkKIXfwzzaUoKnUaI6kI
9972saOOods3a1fLCKaLYzSGZyMfQMbZ0FGEvjdEjNmkQ1NImrZweNNt4F0BbCxM
Ul/bpKsIlO0a2ca/oCrVH3hR31ZBhF5p2S6ccquSLhr1m38xhkRQQc5NcEV0ZLLx
XozbHb9uHk5ODRbSHxPhQs/SJVZZBhOuLVHU5pG2KKxRGVzK+QEXLINYzOxQIG+e
nUqFg2ViKc1JfXJIQTqJdR2kBVR65Rk1Mo98P2itG8sDB3W5z7H1eM0olemIS+KX
P5HLKwX07NKhEy/hmJyx770TMywclxqHm/sWMurkmniZMlfqwRMqO4lLL0IAzd89
JiLYtI6lnQEjIUYmN7ZYzD1MuwbgWqar/7eLv0oIGtkOfNeRxq7t0plXRwTCb+O6
+3rRhU8AEGClUS9Fp0waK9OhN0mchvT0WSkPcZqoNJRELr8f0ui8HY8TI5bMHDEV
xNbFjH/PAsE9xauIPled5WEl2b+gmA6yUoQfUcGULYetLWApvCUwX73yquHTOiuy
kuGqhZIMcGOIwpi4GpnxiZ8JQtEjh6roZXroYlBzJj/zS1qOL2p5hdPhtIe6qp6b
AoYSA/5/J5mZYWTC4jR3B4nnDIa4byZZrPDcoaAHGNr7NLp5z84F5SAt0eDfhyEu
mqDampWwN78FDAOSLH8+A+1edNteXSkqhJ4Cloa0PCt90BaxOsCumDzEV5Sc6W5r
aVL+2/jA0XuTBL+wac5qqRrtWK7boEOM5wvWbLI4g9laVemihBs3X4RDMsfY9LPx
QX1gjHCSJyMdHMcAIi9siPEk8Yd/Cx9BCVJ8kMaUT9XJDg/AcH9UcpH0YEPqZvqK
8NL+DM/sw5YzqTN74dXioyQo7AnIaz66D6lAihWrg+jiC7ousFjn5rFRRNgsZQJq
5zeZAekFhQggR88SlH4tM8RxMZ9Zm0bqreX+EqOQyQL1CJFz4iKuRiMsDwvdxiQK
8p6tXM+1P9Iui+XwuTY6jrC43r6DIDmYpObnncsg7VP5i96ZVcBN56rx2s43Mdmm
7468S2wloVxZ6JGrfOKG3YIPsgz3oqxWOFyhwR5grXf/QxyvOiUgWyk8ciF+CVAH
QNAmGCB1+9FeMfNdMKRYLJjZTIWv8EREg1kQHh6jq33O5k1mD9B7oRw6PaHWrSDR
63J3Llr2lw8EKqCyVDmHuyi+siPfTa7uXB1qTwgVra/0iTNeLIAI89lB8TeS9xvU
S67aoP4AvSDUHSAR1ZJJOz30zBc8+Q73T+XHbTX6sFetutQk/0MnYjGglRfyEHxk
QF0eGpiODcnL39e9QSavd8ANPyL7IWZ3BQf8amvs0u8PeFVJoLOhOYmIe4SsYYFB
l8JfnM/x1dUaaTOy/BRsJqRHX0HI7uezIhM14c3e70EKUlJtL6uKt1KJIC33fV6P
s+3VQpm3IFHVFypVcLVHnbbu7mzGSvG36KAue7EpBDyxI1ziEizDKPbwMQGCx7Uf
pGgj2TqdWCe5qNUbV9k+B/fPX9X8ZwGU69Q2ycWFKC10e86X/rCDqKaYoHf6QIBr
Vyg2CKWhi+1LmNlHq3a62NxSGRcG1A2C7EuAbD1CqLu0iuLPbocYIAoMvF7n/+MG
d4u0ZPOQaB80UmhsTcXSVZItcON81t+kwgctui6YP4FEs5cmY0P3d31VY+DZ0tl+
xENtnEzegspHOMKIi+cPnVG5tyYj2t3GJVPHWCSJgvN7koc1BTYHn8/92ZeD2cTi
iOX7n45ZiAg1ykIUd2cAn2504sHw8jxGcmD0sCffHW8sLgdnLk2PjjH6PYTT9cQd
xlwLRf6COCRyYz1AdLRaMAeWB503HiQ8g4zzo4WrsGgKzfrlqGgvH4+lX/2z8dFI
R1pKBPslM9HkTUcHtDdJ59XBk1mWQ6jQajotacLOSkUf9sLf0g/7Eb6Xls9pHXFe
htrP+A/KKWAiM5X9M5qqdkkTCwJeMmlCuYxMy3JLflqSibrekUOeF7TL1o9cPktE
+pzksGowkPjq5FSwYUKL7M26CCkiYNIg+oRoq3TMuDl2kpgJAY9yJlxK5FQkwLmY
ukklOwQNnfwjCsOvjpG48yKffx9/7F4U2xyYvlxw6nqt+XWXhGPP07RHcxtEwNiS
AtyHjXUvHo8o9UclszltL1aFLWdNri4aRN487A1XLhELs/kNCVUwnERfQSPM6QXl
MulsfaeuzHIdFf+xnj4Ynbqg3AuVkY4CjQAgx9LzDqWaFBiZwG/miMeUnjrpNVbw
hCNNZIwiPQfnYLJwJ4pf8T1UdZ0IG98y23czgsmtYMvCZXL2+5gIuC/1sO1yBbMt
doXT1EB9IXH1c5iqd03wr9iFKso8Fa3BXO9QT0qAaJ8q2NiOwoHHi+arbmL1fOux
8HCeW2drg/T2j1ICPze3Ft1AEMSZeEfDEsZpiwhw6OuNMeTFWZmYQJ0a46eCNE7z
IpfZp7DqJZ/Fdq6+qOgJ0V9iZ8ScO6/o80/bzJ/8RFC8n32d+h9cy3uqhqkr6rJx
mnYxq9qT5jKZ1U4PotqfRLIjLsLyy2OHiTu6xubz7AtYNxVBnl0bP2LVYfy+gqOS
03d6/UpE6xUdKLGobU6o0XL4s+l6RdZib5t3mPQe57w4HR7kggUukvgWMvPu3rP1
4fwFTtq29tKuvN6wKo+RHMOGoXRJXDhnmdm+fqIv1/4tnrcoDLgRkgDJNzX3ldZU
v+gAVqplWYUhnfMAOL6W2e06aaWlETF1JI9ngLoWxw7vjj0WfjMbod40BTH1E1J+
3rtMkmfFNXxHu42Z5SFhoDdu9nWfHiuT1Utwkjdasq55wKdnA7AW4Ki/6zcsJQHR
I9M7n/T+hS0AiezPOWB0ORVCDIjK4lKIe5wDzOP26f6gdkQ9V5aicsxBjg/JGhRy
oRIBtjIQenFDyFY4yMpXmeGStWnQRdCjZKsaknEQRv4pQMZIRxCI72H7ejF+exfT
yzUujMK9yn92qoYDM7K0s3CembJ0QSIjlIsCPFtJY+Ff36nkGPhUNkVFT/IAqMVM
/H+3VdAxI/NyBIABVR3pC43OehcTpU/QK/hq+J2mwRQJfEedM0olAFqkqqQf2his
K3jn5GrIZx6ZfnumbvuTkptHSRnog254YxcYAui30y4HBlue4n7Bjj2X09iXzSoN
949mAMLG1+/OhCj9PkrJxrtxO6NzpEDpoyKWh7H9UV2+mPmHyPRGHSQfSHjXvHmI
LXOaNh6wlkGb6IB0bysvgwtcIQK89EdWJp5vZDZp6NYf4EShm8agkgcTCE2fkPCl
UkixsjCfY8t5Edx/tTtKTvj3CKxMLyaNa3u4+BX4nPwvNtW2CZbd4WPj35R005ct
h5S9YzA56BcKdZLsqyY5TZpLOZlivBI5DkZESFRzCExT5CbXtS15WuVRxZk+87k2
Xc7/AaBkFm/1iEL1Tf3oJpHwx0mSJqeDWZgkdnk5r4k2wmhCf/RaLiqRor4EUSNx
Dnfy06EtH0jmxQNe7U4uwoerLCyBkoBkyomKAiv2hAE8JstEgniKoXhGzki9NUr4
6YylkeSWscq+KwFYPBbBjyB1Cd3s2zxjlGWQEwYM3YK0XOCzxeGPZf2uDxziBm90
c6TzikZt1YfcUHuEL2VV8rFwrZHYW8oh+wCpHM9ipWoMupwE/ckhksAwI5FP/1UT
beqoNk6/GYBq9WKHwqHmy5ZwozMYvD73yj8CBIPwLhDMtKmKSL0DlejWthYuom7T
dNsTKgvMPZiF5InqUa/iWemmVz967TcbnCGtn2N1Xz0CXJuOy4VCSVs5xB9ate+5
dnWrM8PRaV5foITuVLFnnVAR+3nR9rwi9271oL4aWkjcdd920KK1/VPPdDHUbILJ
igu4arUR8xOO8R8SD11GHP/SLlX8zxaAFSp6pfDUhYF0dJMVcQ8cu4Dyh15uGnoe
S0Bmlt0OzLukmAZsc2hIde09Qpw9iChz9qZvYnwZnKhhB2j9klhD2Q++WTWpQENa
wJWJ8ckytoY07uqDFPerO9JNTFI4e4bIWi7xAmTn9RRiWFs+obF2Tbb/XNRJPPB/
ipU3fMxVc8fYQqDCWl/EmN4KIe2VFB3s9VgawxWR/Ld92TccKzi51ikmiUbQqLaI
I+Q887lezTJuX+wMtwzcNP8b7FkOdNTFlFJiE6FLZ07c87we32RVQcCgs2GGb9Yb
lyZelHzutXZx0j5gx7Kc1anRc37FtvT84HQDL5AQa0jJP48gzJMVv5ezcbaeqM9w
hlGNrQgQwdyvjjndyomsynro7exKcqxBNqKbSGhMwt49QfORKLwEfMF26bRTm5rl
ZqOSC+Th6UMzbEQAd/IoIra7sSwd/c/vH+hBClgMewz9WaXQAz9YpBwHXH1VnkBN
iEeq4gsQlWxoiyYwpzas4TQZYqW6uiW9D9JAIXlkN+uQmjCF93sJ871V1e3oZbmt
krgR53+COGaPEkl2OnwQLLk9eOCpI8s5ooePwwf5OGP2HmkVGv3tk5CPYIF4FP6U
kFvFxIDOY/Ftux9D+b+x62doD9ggAYTUIRfjYBgx3cYv3/ki+l/jVH1d/uKDcPss
tXPmuat06rY8iQqeLnBNAgiePHgdc9IexZIBZQHUYbi9q3PDSjR+7NLW8IQ8QMaz
n8jrgBJdLL6gjgyuMJqsEZD31cyAGCGWHXHwkocGDy2aW+P7z6E5w9gcsU5suhr+
fwWdrLV7Q+Pa30ypIV6++cb+2UKl9NPK08pqjxxc4SvfAPtd0yuKf/W/TJrN/R7u
Q5dCJ1M528RKpvwYZAsR4kus6TkxK5iVspR+35KT06wWXn9wnjNYsweBabJ7TpP+
jOCX7dnkLW99K1AL0tIGnDPiDkzRUJVWfWT9ju2PQZZeV91SyfqfFWzxxbGt8n0/
6888OxZzyfvgjAKxToyQO0oRpUwXhiipNdzpRs4WYqe2q27V7Vmssj6e+YTcFX5z
YBZuzyFXZMeH0mh/xod1NaBI6lmX2fOPu5a8LKTAzJWOfL/Zb79NFy/+C+N2Enc5
p8XU9DvXdHlhVPMH2lYsC/c2qJX/h6mJ5ATmO21McqtVl2kVK+Tlr3N2vDlBbYKD
j34xC64+M4hHYD26FXhJzgAqEoYYyLqyAt2TkdrrpREq2HV1zRzGjvJ4mN+7vZrB
+t0SGXf3jgwmmAtNKZlTu4P0yERfia/U/sUkQ0QwOsEsEQtUcVnEvIdbl7quvnVX
qTggyF3oEFypSewWhC4jKO1VMQbRPMFBsgy8m0Y72/ySFsJ/o7wFecMzIj5Dt2Gt
kAd4sNfZBBGvYe2ZblMQAqf/74uBnp6ZVxUw9o2ltXMwe5ATGa03HUXZblKHKG6q
lPVrqpFLzM8MCxlgaRMXElZ+kF5LFsYXxw/q3EwIrq/V8ziYxglX/QEn3ReL0Gt8
qZDfq8TYS3sw0ETghH2nRnfKcHkUkkMPAFOoNX2G7H/4g/zdHiNkICfc7VqP1YyO
X2HpfgJH4GkhQK7ZCJMUHgJFOShwMGRv7CnHC+S7XxBIBx1jqqFmygDrulJMZREL
lb6bqnKcf424kpg8yFjlKNOEW2Ud36tZ3fnYuzIuAzYf7qtCVBMRRDH3EKOxaimz
/UIFcVGhd2A8c0oWQimzf3AHlXy25xLhJJ/GYuLlwjlJbObIc/cFB9jGSXTNYq8b
cZDePh8gX0/BMA7aAG1iSeYtkHO+PdzWm/tjRTmkT1DmXTVXlWLr33DqtheGsB16
lzsIgrsyDxBezNj29KAgothmPPq70ZfAol9EIj+VaWcrqa8hC4HUoXyhtm3tmFx9
KpcBbPf+5PSozpFb91A4nyuLEV109DGGx7nqSHstv8pvIV/JpMOPDFaorvSYA6xb
s0OZXt4qCG9AFCUqUwBUspnGQ4pP5/Ds3im6+mNyrnCmGGbSo+cqRaT58PiwKUq7
z83NRELvS8OodevkmAu2zd6bDzZVzNjk2muJfmv/QJ0qIMKaAEJouiBX31DwImOD
f9T+Vus5ST0AZGEvhUnwOpbQrR8lI5PgTSjJ3wmpK/erE4dyrqnoaUEGM2U0p0sk
7/+5fDACtiiTNNlmBWf3EItp6WBp6w1Hee4CnouIZHj0UzaPGAL7fy9ikLTVizJx
kTlAt1yoYIosJOxN24A95JiTpN0HZ852VFAIvsWTH7kcwLTwR4aAm+u4flthQ277
PhxgmPpt6F1eH/IFZ+n2HC4uOzgfKyVzeM5uGEYBrg3WCkvvTqcvrhWvzUcqmUKR
peP+RZxIyfSSUZpC95Re05DnFBEzGAcm+6WpitzwO8BQqMfNZ/eZUqwy20lXy60m
15vzZAvcmpXe/K9zwzNDqM7gtmEnXX9lspHHb4cmWpQVzwxxREd91ocTbrAxPfii
p+XWN3Q3LFY9SK9h7z1gCq8qeA3DgPd4kT0qwPd/VyELzpytZvQX2Nk3qSqjkhQB
a3/AkiGUlwEY2DVQcslPz10a76GeWQCO0UYPBLzD8SFpcd4KOGqz2GDC919jKKuq
vIugnZKplSRr+IbmSO43Pw89yLJjTYo82c5+bAnzi55vf96UxxLKl0hJxTdyHWXi
p2/+pADDFKKry8QNv6Oio/e98SbLQXr483tg4jVb1Mm8XjMbu2Q12cMn2nODgS7X
pprD3TMVmSljg7xIO2qxa+fXaHO8qXnFV69aLFP7zsnqwxJP+zBNXmrb4awMyGfw
EBN45Q6Y5hsGqsvOAkgDGeDRv7PKuDVX0HChGe3tPUwIFSkEX2nbOBMRA5hhkwa9
CGGMDTMNPajuOX6SkDrSTNd8TswHHp0+pPHSzj33s70sjrL9VAKsjEjqfSjq/CPn
IiSS8N7o3fo3EUZzXcmSPGj6W8SIso7JEJWyTCY2UBbcMfoY69w6JCWSKhwRbeuT
g/xgV8KjXpspaCNLyhib3L/6KKn91RX6rwRrWBIZ5eqrSYlXsmNDz3h0TFnEe6OF
n5cF277S8jwnb86w8iA+NuaUK3QL9xrmKZVoYLuYkRHAhM6V83cu/0SaFMnlqV1t
TBulCte45ffKudfjdJtYdAHofYljW/FZMsRtt1TGvkOsJP9wnAUMeS6x80pAp5FO
Cum5+BRB6wne3zaEPw8x/ttu+d+TCcv79exF09DMI0oolIKfDc1qI6kzX3CRkVSl
LFrn3DF6hifvZQo5aO5EOLjrR8MrRn7lvbFgaABzKm2IzOeLo04Q2i9UUhD0Tpvv
efbTi7TGkypfvIxAvgr/HmM4jECvfMtF+EqK1wG3tMfjqij/vK3hKMnLWSQaX4Ms
Ti07yMYaZI+SH6ruDxDnx3x/QhjRsBZGcO83JYD2L1lAOaOnZisj8Gv9Gg+SX776
+xxfPWzQUhaGO2sk4YEPPPUUT/lTyrUpDbYGGV6p1XOH6IN67VPwH3GaEngHfT66
ssO52YGgs/Mdzvi1ycDeQ8LCyfvYw30Q1geVOH06olhKnqp3ESpzPgxOUpS1c8TL
EQo3tx9n93E+YrAgb1Gy6g0RTTKxeP8pTA1p3ktPAtUewMJHEWK6YEmyTtqwt9wf
mZ5OE2iP4hy4bnE3m08+mNfQMh+fI1XnUe5UxF2LYPYTmLmOHtMMLGAb7blAvcuU
f2m1dXX0sF12sHi5oJfN+Cm+xmkYIpelUGzbU/Sa5fxCb1tep8dAD6nA6dNr5Fhf
b7Hxn5yqQSLIrkU0JH7k7iLypQRe061WPui7K9usIskcWOpxUM+g3At+SLMnrHC1
KJeIMBdYB0/QEA8RdJ3Ib0fOnXbFTJ1MkxhjoCx470bJeiXORVeH61ZFlpQosWzV
PClKoC67Pebw/4nlv1v3KCCgVWq2ViHJTKlGaqPuleyYQV10QYXyJ4AdkeBxeVEo
t59M/AErYSi4CitoVi0alzB+r6a3FBVjuZMf8wT9DMdm7DYoDEPA/1qdqbxlq3uY
AMXkqvesGQXjHhNNXxxdvtWrUGhCn1nwdxLDx6FgmSUBIfOQZfiHfULBxKTewlyB
f5amvgoOvnWVh4DfpGnnwkxGL/mnQlLD9ec6LUlsLlU7kAp3YEgB75muOR/GEB0q
6HfK3RWqhDRC0FBy9dFmdr8LqTsyIAnBFS80FQlfloMiS0Fzn0YfJngbupaOLJUN
EPNMeza0J4pJx6HgzBoH6TJwsczCz01c7T9lH7SaHvjtQ8DoRK3LZQm7PkRTwrqG
RfXYpkt25urN5E0ipPoQ3DeS5SC0/tVeOXmqblAdkWu1up1L5e8YetUrsz0rFdL/
yFnQOzTsWxc49mi1gVb4GqL2iHbHgqOfMDzgDBNai1NQAYhJQhAzCHkDFCzStzYd
2OgxnVsWEokChdbUTFKslHYgoToP6M0xva3mOgGo0z6dt0t5rSOrvhzY4AYYYr4A
HaR/JoMjgQ5Epiz6qww5NgUzfUG9kHUUOySQH4SfAQE4zpyh+PQH+pbuthZblYAv
EF5Oos39ch1MDVdKGyzWBS2VJgdZKpvuNSI3bFE+ZHLJx9wwGAz39hTXVTvGztnG
zuCPZLFSvw8BZkewPHf7BpLd7EPtGFfUiGQwnZ6cs2XkhYyrLJUqTHq8KBSs4+/d
tzOcM8TO0htuX2Pq43Q/vSlg++ARev6V2S7jh+4KG7KWAtS1pjurbUQbaSdFbcse
xuINRdFTCTLqnoDDg8I1e3NJHxzf5K57aHEYHz/kK0rdKo7a+W7hAAjaawf/n8V8
NGedgrP2hlLb2+cUNklgVebFOUMaiV/acEeOGElEon2X7W/xEDjMu3hs0WgI8rzy
Y950HWxsvOlYjOseOs0LGI3vV5Ujrb3c929eoWHl48bBqBxLrpIDftUnL9yHE04+
s8ybVpUFenJvEjT9yiSOQtKMbGRs2V8zWyTYtHO8E2kl161EdiLOdJNd1tLBeMPD
sAp1qpDPaYqW2rblvjZ8+nwYKEFBxg0Ceqpz+Mzg6L/pUHfzcJuM6wbw3CbdycIJ
9+o3CvXTECiaiBlfBPtDfrytWmuIxa64A85ImxURIr8ikCur/p1CzmdrYLfhmoWj
D44f1YSRX9P/flBhXp+u6+2i4lIZwxJI/epRWOGczkO8fcVPBPK2hX6uyfU12+t9
ibcvImYPBpGLazDDNpbDTUjHDowR98aDWgjtMAwTHype+ec3m+Zy00AUlo8K0I1o
5hthXEAa9KCd3smEQFfenDWXIzX5YBnVElb2nuJQ1HKlMW1tHGU8/pitiH1r7u1E
IduKyijPJenJBDu8JlWE+RaNYMRDDwfgos0zesFAfuSswxuIig/e2pnAcYxWs8CQ
/ycuEBznRm0YzZF2YIW3tiCVDl/5JOzOC7kVkWy0mw8xWUchcgJtzYNzneOK0fnD
nQKibM992cDJyFuvvpnbHDEoKcsd8BtkeypuPT3OAHpVQaVO1hvQn8axDBRwjIP5
ruWwPBQrDqusB4DippuwgSX0VIzqnHDpOIDXa6MA109Ki6CtVlahzM2U6NpuFmkU
NkJkhVAKetRHTcxNmRL5laUKZvA43mPW8G20QLNkoWifs6ckVPAof9CU1fLYQ0Ox
RYa+71sFF8Mn+vdR74X73btgKsvRC/4wsFrfU2HqQNjgHTVH6t8kfTTm4kw2HDdu
vNiuPjTIu6osBxhQnvxthfEu1QfD5Nn/kmPE4oRRPrHf0GqcvvI45Ygov+TkrQ1v
EFLGRyKKropM8A6Nrsad1R4ijSlSM8txAxcJ34a51O6Y3Mce5129a5pAj9Q1UknE
C0KZbx0c7gQ2TQZGvnZtSC31oqni+ka9qtiis/VUJ/1eYxCuXg+5Lh8zzPYtBqjV
vqF5MWhRYqacOoQ/23Z8mkOTPQNevWr/1qXT/fvQJxjSYq+bjOc4uS/10jKP6JSd
0HdxMeQcfWO3qNsHbCjnqwA+pge/MEa6AzpN2CHtxauzIRDNMJAHwWVBo5jbRXRk
nnE5O0fq8RQY/GnwGHbge/IPKjn+PxGrwtV+pDwHMAD30sHoLrXqVpwDK+h1g5Ng
YwShMx5Y1GyisrH964IeQByOhy6Eq+VBFqo4YIoGn3bEUWs0AgpC0fnRRaq/PPTB
KpCbEH11dRmlvMsdHg2o+YZQ9JyinyQykyHuZ1JZEScz3RwEOoLjVEFgge4sMTJL
9V3hXUeK8MRa0kBkc7eFN/d8Fo/86MKH0pd63g7bIdc2oFSQUzibFpB7oF9eIuus
CGDE9tT85opIXHmFs45Qm7lczywCgPhx5Nu9rnQ66zPZwTnMerJX/Z3HixCWxBG5
yhVBJ+rlw6aBrrQPx9GM7v7N/MGcHfilj8t0esqHUqBC8scO52dgJ14QyWecNUMD
MVwrJAKx8L8kp/EGGhICkxJKzSR+uDdXu4+BdqnMAHi/z5P0UUuRmcEIqmYTc2z2
W6ig36ZGt5ohH8NNKyvlYVlks0ubB2MTJYisex0WfX3TnraJ3+E+NNWxxTSJqVcG
e7POH1ijkjLhntXqj2SE93kkKYQozuMHAzLSA50G4oCNLeySRJ92tkTmlJEpP35x
jlVS77bVcjhKsnczETOwr6D7k4lLeX6QEAeqGLHvVatAVesCTX2mAfvHdAuGmYc/
3Xf5n0IPW/mvuC9qOT4U/tbNd/MfXUMTgPKlQPQ41a94g1yL9z9CJVEUg/C1IRNJ
mKivUOhX24PiJzVoQRfEmliSwDvTHcLhHtvtGk7Z62o3//XygNzOmMaRVMc/znSn
dfBoXcUZ3JoFKM12Y3YDw411MwotMyIQQtJ73yh4tFainqSVgpdyd+i5dFwknVKq
rCudyuaz+axyz+9nL8EuCg5L6oSFA5oX9th3hPFb+1KF2Mt18s+EQCefv2+QJeF0
RIuvSRk9Df+3chMIVNnr13LXeuDxmGyPaXGhs28LVBQHcFcBBppcA9UI+pC+kJeP
9hVrniEsPbeCFGzgsziArD9uuAjgk7zqKK5uKnNytE2/EFs7PQj9hl9jnqL3gT3h
xA0J+AIatBYtqX+c2gktgsTZE6ILrKbEl6heOpMqFHeRO9HmSIKpWVJtByJdx2l7
RbO6IvuEAKsjU+vkKfeV2Dy+PrT544MBoA4D6BLz1u9wVMBr+AWzlPiEyEk4wUqu
ntQvLYDqXw/m6chO+hfdbqZpnQiAWKx7pQaqwWKfg4nvKj84lOFJU7ZyUZUEPppG
shEW05Xm/jV6Hxjaj3rzyMbv07NF9DcVIIV2XROYZVTAPzXYi4YzJWhXuVP1Bscm
JQvq5qaidWpRHH06JeCWBy1Y44ML/lcfeTmEe2RXdXJ5YTKnygPRBgggUi8sMx6u
gMIzP7PeGDoCm6k9MMxjqJ2ce091EAQhjqvxHiWUImn59wyZYtGytR87FPrA72jr
fh5ItVAWLOQI3E8u+Kg7fO9A5mOpf8vX0h2uAMKhkOb9nwAUf3lQWd+Hdyq0EvkT
/bCb/6ovFXyL/4hPXsHJvWn7i7rA4ZRRCEiUAt7huBJ7YPheKVTiJwk2gaCM7EqH
868Pft3apdpe0EILVmigPlMdUJHEYc8U7mnnr604mW15xwWSKkrao/XOfSXrelJR
HY09HTtwgkcIv80E4qujIGgHTV1hfNoc3xLRWAEMc5efZCwuIye4qeOMRoPqlAMt
uZeVALOmWI38SbaK5Ht142arv/TFnR+UuY0CrB+tRJS6+BCIae0jl18+1srC3YVu
A8eFxXhzAxGGW9cgMls9hk3nSO8EZkVhI/pLajSmquVB6AjCTTsDHfeZkjvD7WQX
iY9IEq4/VvVgweWdaxhX32oBKlI7UtOPb8k2z1jZreg/LjB7U9EkuWnuyqXEvnib
Fj52EQcbzdqj6wZENB8Nc3pVtutpbjml04X3R1SRaykkF4AfOPb2pKPsOpxoxIeA
GWi0fj8Hd7pk+exrocP4zUCXjakfkr0Q2URtNyFfpisSjzdyUxwfan19pxNLoaie
4r8qE0jsfzxn+UqmeMtFlU+GHt2+JtT7TX7ACTpoZGIADu084dni7+u8GGr4Cvj2
qEYNs/cReh2V+pZSDfFkrzVphv05KXZXQ+ouc43eZxiSEtcexFwnIHtsNDaUsBsd
qsrOVmV8diSJmO1agTjvaY7NzRKibih5XNaWyweFNBJCdFSHmtURhHE8WNedA3e1
7sNkC5fSIYom5KHGYNcwH1TYGkzS44iWCXRIRN/nvHd7GpoVo9hkJ7mbZdTrgb8z
Ab5JnMBPIJiS1mWbKBCmI3et5SyvYaDVAPmxsWIHdcvqNS2jwYNBkYfLq7Dmi1FD
gS3WlkJlCHcyerYCHxpq6mTX6a9B3foabtmFpvs6cZJKohqY9KJGvPrsrn52Wr19
aK8AM6t9Z2rQNe0TezMEgv40hux8q1KZ4XbCCcPt0rxwAyBG5ksvS7ofXte2WD1w
+PM6oJAOzst7YSU8UGxxIqrpHlFF+PO3siXUW1RcG9+R/LiyHtEuOR9Js50kwzad
u2hGA5bzHLGRqvk4jNPuDP6u5ezBpeWV1TJjlsLdel3fLfVDJTLQTlG+LW0+mG2l
aoYq2fv1p1xTAwstbeUhCxieLzRHFCzXTCss1/02eRYnXSe/EZouNZ9nKFYH7EgM
KowTLIO2Vs5HhsS/N1oll3Xi5DHx0O62NYkOpeQgouCvY+WnXXSgnindqsyEvPFh
dGVAdV2J1ZgwScafggn4m25Hrxx06vMCt69UyIhXvVGOUb5LVT1bwngYaQ7Gawly
61zF9vH/iVS4oEbBDyhAP6LjGM0fyM785nVxr9h+5vwEy5E+gEQzGeOUTf0mL67N
aDkmOyxdkxVBuiYxFjXZoSrUXxUiEms6Av3c+rLW0YxyCo/7+I/UTSHpohMV3lYN
ep2KuhqTCXGa4Ws7E7ywvdon+T9hJuvR4AqRrUIj77ZoItiue5/R7KnhfLAsVEJt
GGG6mWdJehQ3ud9DvN4LYSInnVqlZbz85LQxpUEkfqEoOj+HHCcn7LIxCulx1b7I
o7F++lM2Lm5QQruRyA0NP3PL9ZNoXOieHg+oKCZ6J+yoO/rIpychOx/v2ahtc3cT
2k7qc7LCljOuJudiQICt9dBym0BI1OiazgaMkSGw0CTYrilwOLMRWRa4DcYpIkUN
k42rrRz1gkNR2ugd/HO/4uGDB9rZSO3YSFrOH9zUzdRQdrE2OvPfVJ4N+Q7C/1Jj
0+P48je8Npx68OUAWcFYK6tkI0NxRILUHHXv3Yj52uzKivZEjB03NASMV9o2P4on
M/jYdte9o9FT/qFeKsHRk31Ap9Iop1qjskKv1W+w+gGVOVt2feyrDQ0TeuS/dPLz
hFAKeeEWZ7G8OW2ty8k8t+FN3m9iIzaeKINGnXZ906Hgeas1GaE3oCzfn1N6B6KO
1ut2j1Tw68xdVER/2yOxEEiJDosOl/CVdTMmsJMU90EnNRdPBsbnzaBqn7dgHID2
Sooxww+WBKtfLimUwdORZdJ/vvchfO4DRfzeKHqMOXODyvktUPGvGvyuvF1QAE5M
k5o4GACyp0vG869KWZxwBRnaPCxpRRFTRzeRt9kjZtMSGv36Zbu4nTfD/olYxvfx
RJpBh20ZIAoyNVFV9QpBEtU/fou4R2Uai0W7FAYn/tNy7YEUuRbvuIkMURE6MYNk
9V2gQIe9Motvo6kpgAhHOmd6y/bnKpzrxnMwYQBTGbbj1iDgAuKFNHfJzDT9D3vT
Km27H+KszkeVkkOHJQUiwnw7h5ETnbC7CQrn12douOnhN3+mgMSE1mY8RZV8ArWV
neP1OwBT5oQ/yZ1goZ6pEA7Uumth9sIjmTP8gGK50b4ksGs/wJtcnnVqtKtjpUPS
k/aLs3Ky6xeoi/CiYqgKDsCwiru4uOMRo8/vwCVJmy/V3wGhR732VVu394VVhFbO
2vadizri5/zvyjZ0igUkMq7cOSbFbB6jNVNEFxT44HPvfVJkthkajrdd+4nYqGVu
cptn3RttJ22/LfvAlcYoOewNGz/34Qij9VWl1ufbvLncdpEWqjKV64H5AJPG8Aty
/o+/Y74tCFBGAaC5qmN5U9AyeuMMzVpye/v9BIFS7m6c2LG/PtScfCgD7hU3YLC2
8rKbtUGIM4oH9S9aCbK4fTiI+wVOSiikJw5J2VmsRwZhTT4mw24EMWmSCJ9jwG88
+iijvymmjplTM0+m6L8OLABEIOWi6H67onfWkpMMtKCDSS4yxN8c1wr/LDvA+JNJ
+tRFKyOMviM3fdQMiLV+ww9UaJhbiu3uwUP6A2HDRf3A6j7WaNwu5WRRyStBZuQO
luEvIkH8bsaiKl6cYyjB5viGfOcjYGV+TPF7GKW69APPJD+t2xEHAhFJWz7gqJfl
mZZ6Ust/eQI93lpRY04wDguVr6mSmAuUobEEe7yciNQ8+5LkBcSLcU4E1guJT7jG
/mdas1LDCvPUi5RHCFxrHFwnh6KpLMstPoAvpggaQOJ73cazrj6tKnTDoPRkGDzB
D9SD81j8oDlSQqrPWcesfPMfYtQbPn1bGfqSRdpKxKPmpSiP0o4Aqqh/LOkxMYOm
A8NSsUUSKg6eDTw448eFAS6l4DEErq0hgfbrAhk2NXJ57Ts7VNgfYfGwxLCJjqLz
Rg8wgHeRdwmvRDuWtFGYQ27rziebfsWkLU9+Gg4UMtgMpEfQfzoocKqze0rq45EG
o5wOYowq+3jbkOxuEnlTa/2dVnW4EMcTgizjF93OYKWgEOFdNHJyqq9PDoBdBCWh
qOqQxZ8R9PwIAXXjUUUixJl9EXx+wcIlHU3uUyNHnEOtvpNmCQnl3wcj/0xpOJK3
FtEPt3rTkdNNBNo/pF+qHgMvh6Kbm9ckQX4HPFdK/LU74k62OPgFQaNOnlcnCN4g
MGmMtqDdH+Yv45nIyu2GPs03cwr67tM/a2lZylOX2HeFuDd7hXKzZt5SwvHcGDsv
0i5n5M/SssCQqaC8O07M22e/nyFnlc4DB76siB6UW1puAdmlvS9sDXr6HcAq4s+y
72PBJu+06kDtv7URVAcvDsZglzRUDzG3bfVUzCGp+TcRamBLh+eoquG1ICg7pibZ
ecsnVWjIHiS+CxMIIAhS6NKSYaKRKR4IPGv4iFb4SCoCYz5UyxtAdT4X0vwChMup
R/GWywtamvbCyXZPYfIGyGp8Kfr614AKWQXGHXHJtqdA8q1qunBryaosX9m3OPar
iRrVbkIRcAzzF7K7vBfHkOMpPERNd558W3zNZQxxemOqoIlbs6mAXSG1K4ZDX9kO
3Ckd+fziNW9yXy8+DpUkcoIJExoCpSnVX+ez7bE+kXwyAlosm+E6m9kLNMdxcfoU
6oJzScfm89Sgik9ZdW4gRqj4bzw5Nsb12uTaloyZ+72hckv7BgQ8/CfeZvjb65mF
PY3qToKnDIIzKae+T94LZV2MspBZ20nFrWlS+mDzQe3z/qdYaswnknalU8ncwUJE
l9hZQvixBZxZGQIKT77vOYnJSO1CVXv5iT/7fgNyqpSzf/zcQ7UXLuWH5qUGvSW5
y4gMHPenFeDqyqFrm6+M8aRuSPT+tu2Jk54trhVo5v3QNC6E3IUXp94QL2VeUEFD
WYhCYB22Q4ZKUKsNt9HPJAMWdU/ZZdMOEQnjyH+WdG8BuBv9kul5jZcYm4rrmUVF
oUmtkZbX0oVR0QKey+Okp/zoRuO8ulcak2m5pW1J+ebHFSaXhxxKYqp3fBcFES0k
cGVB6/LpHmJb3FnYpMIr/HEqtQ9rxQSHiHJ0MTwijdn/gF+u4m3tfoDUzO/YHNe/
Ryb1bcMpfCzp5Ued/8tRhx5A8EVDl2Ep7CsdtFl0R+heAlxvE4vCbf39Nql30tat
gSNImcseLbLJklm4BFL9QNxjbnel6JmBNtbgOrSBZpN9KFy6WHzAtKMZrz2C/geF
eEc3uWPhRi2xsyo/vMnByX/UXhReuN73hY6uAVsQ4fFTq1NZ4++hP+Sj9TLxHYIr
+LrgGqZ3Tk8AKnbqojqJrrW1C/g4HB6XRRzBOm3n0veMVZZCuB0KyptZNK5N/3tp
/qc9VXKmcoPWMj8xuVpj5TbS82vS1eR5boaBin+w7OsziHFK4pgTYmL8SpTF9O1m
y65l4swzy63XBo3N7/UL5kNm2n8PdjJzMfyPU6UlL6a6d+M1lbbzBU+KaAuE3rEg
KmDNxsXLUhBxn9HGTRmAUdw5NHzR9OjRD9iNq6UT6ssrwjsOGKWh3krxaAUuIHTV
3aKp+2K9m0YQJMkNimJslSDFd1VffoJ4as5un2dPqqcKpAytH5lJKhOOOM/Q7o8w
k7cBQR9CWEqp/KSSFKG9L3VFRN+qcmSIsSj8/4GN7pJgUlJgextx/sK2EjLCbR7K
A3CBp/dJEasj4Fe5xXlgEKLQfsLWmB8d6+D5EFG3b91CG05wQTRNnlhxhOa5A1LO
IinM9sNLuMIUDYsklRTncAxSTVfD5rPtcSu3Qr1G5KdaY1izZzroMzT6n6+6I95D
hxWNT+i7YhRSPHRmBG96KZfXGoJQuoNQRyuLEBGqgkPKSGk1mjI1+r2sjZ6iWeDA
datoD+VobGxHRz/zNrS0+Ma+hdBoKgDoOeDdblD0iNgLEGc/X4YGZmIeo0dzumiV
IpbR3qaMCXtH7JCTIPl2EHKCBqbc/bNC5DK/RUJSETNldzbq8lETZekrOM0UzFIf
jV18qiS8QqT+TfQtLQSlR+//iSZ4T79kZECvIB363/4wVVOqnk5lLOtnKF0Gk9/Y
GxN8fs3cZAOsU3i9VVnnz0s0mlskRSH2+WmAZDvI1znrMMlkaFwpiZtcAnnnz/DG
R6wQ2l2YsQR7j6Pphln7mZLFMkFXm89pXvGpFx8l+VbPnF2zEXgK9DllTDq+b4Ty
JbbrWJigjtiqed8Q4Th3c+vaJ/LgHt/eJJwKbQLr8IjiKC8UZrcFsRxsQrvusNJ8
FE8nrOQ15JtKTPYWwkZxE6kKKQRQGx/eKeBp+bix1wd++F2RnmHchoHRrBrBFW94
wYvyWnev8vU0ZAl9RxwhaYASywRXel9YIJJWlt+efXxrh5oywt1XT3tPPxo5P3Mc
NDCfBrmonAM6eoiLWkzXlDOKtf+/DCsXc9YPWy2uGwqMOMqXRCGFcbyu6sjKseu4
BHcgjKRsVAx0dq/FX8B7fYsurHq3OhkfUtWk5IaWYmvNlI9xKaBtjPVRh1jk3cMv
UBd3LxfAUo/FseVWWqIBXrv474qEbgoWaTPf6lAFO+pii2MlxVECBE78gIYyVWeK
5zNl6G8oSufh9f82sRbvKqlCc0W3q2pjCJQYEGduDO16oCp4MkfY9INiXJgVUF26
GFkaHiGd5MiLF45Ll/4pgzwR1GjqZsAEEZWvrNHANXeLWggkNAR1LlHJzeo37wRT
K2bBiRL+RbdB5rr3YBz58G2QEGbHuCqKw2RybRruaA/DiosmATCbv7vTIOM0iXu3
PVcLH4QOD0uNRPCcDr/9RgKAXh2whnDVO7g3aoyNfFWA3zWJMtXh8tCvDPBFtjFe
VBc2NuwUpZuVP2QfHX0oHorraScqrv+EPi1NxUeQ/UmmY+wJUtMLcr7BndZPBlD8
2mbnf+l/R1qXngSLwgf2Ua/tNQpCbHthabtgNn5FBg5RU2sJX16FCtHqLdp1ilcq
FImkPDQMMVmXWSTtfp25nJ1nW3pb8NLB2DEPoTmtmCIedUcgbQJPGokKTcn2VtB+
r1PlWFo8AcC2JxVhdiNcDCPdQQVKAaQJqJ3MRf7HHojdPS1bTWEYFzc90KU/UMfa
XJDV6eq2MdeBPa49TK4TubN4mACttzjOVY7c9dGJ6j4JSTMgEiCXz8BVsBHgQJkk
nAXr4OzwKxZeLdkY51l6hH6O+isXRCEvaTyunt0FFzM9JpXiO4bxapjnniB/hrBl
Rpb8SA/DwbypfJA3fG0z0B6TEfJDHVB/OSDG8B4KG9qI4Uj++Uhat5SZWQrqkVPH
QslF9HZk4+SZOfT4jWiYcGySud9jW+1y4kOsxl1r5v3+4N1pwI3CmuRPdJ+xZ0pA
zGmyJRGMnZHN4FZG1i0Lq9ovabEMdDseBC9XJgvaUsO3ln7Ke2ODCj9I8oiVOOAc
SWMAmblCT+pXx5OwSYWnXiIYr5eUJ5yk2FbEow5avqdbjwou9LAIGTPZF7Wfkili
EFl6zo4bSem0nJ5VGQRHvVLjHXVYCPJepUqwSpVIbVEUnNVsIxsagJB95fFoaHe+
kZNpA2DG6beiX0wIZ3WohfxCLJY+G/ga6E75Bpe8vAY3p6AyP2Iakvd05lmNSIdN
kxA6KdrRz7hCKyfq/lKs4LsvemTmjxKoZddfL51J33sDGJdBjuA065I4GeOcY1lo
ojEPq1VVDrkBv97vZQzfJ0jmoICmDRzX+ZVXWWw1RY8r3cdPpu74wU3gRDyvK9AF
Kyr+hVyqBy/AxhwQuWMZBAplC/RqFqr1Gun3T46RpHjMUBoiX9wil6HeY7RXfv71
3KYbMYNZrh1VK5qsaurB+uMYaPggyAp03sk0Ay9kL5NeR5117SpjyR+4coLl5CvA
M9OsPdHnGewNs+JO08Rt5ttuJ+5ynZbX2AI0x3DJ1L/xWa2Ifcs8Lq13tfViQg6N
SEdjEHIIf3HEnn+2bHyvLU+9PHObXb07xd6zEPkqC92agB/hILB8a2/cl21O+pvy
xGucutkmzDiavmClfODfzUlpooqllh1vp50bEQYxYtnu/aedvo2OhWFOaVGrWVdO
brE0aI2399I7Ad6Czo/Pl6gbb1Gddn/CKQNarOz9ZKHJbjR5hUq/NjZW5FKTVLWz
yDeZ8i11fLpQgylLEgUMZO1xSDZx2owgpFkIJ1876ErnotYjOkrYnZ0wxnLrLFKO
7Qh0UPkB+gtApR+AWdNUuJ9JvFWjsl5ngC58CbVtg3/Z5h3rm2m8XfNZeuaeu4iT
9ih5fPhwqrRVyj636EbUxxjF5yc1EgG+74MUB80blLxbSL3WUAVeIdCcHhcJQeiF
C5zTPhLdRfEvwkIw8P745dQcXBMtcXaiv+/r47Sj0DncgP8YdxrZJu+0JBhWpWa5
s3woibhEOkdzInH3oNTMckknrl3Sci7TLBWvG7mjtI6gizQAULQdpxLrVfi+/1TK
2H+n+qxKiOCojXoDJsQMB0iO273D6roftIFWDgLqOeSCyDwOQLWPYvQ1IdQN4KI+
k4mUm1EQTsdPNpjzzqCDl/wJ7V2OGx5rKItn0ap3oe3CZ9w7F0beYy01/7UtbxBf
JwfvbfuWPnalLfBvj3sh2fBBsIlRNLKl8eaAIfjIJOMtsKVzwTQjIinzWtBXKpYA
SGojdy1WregR4R39SyZXzWfXUvEXwokM2wxozRegFZDOgMAMpRPUN/pL0cAFbWyY
z3YsbGDtW0YAfrHdbiPqhjA/cPUq84vgSzBxqOQor9Cfh301b18T52+OCtwaJgaA
oDKb2ST/zX7ZVS+nZkk/OpoffW36nLdNGMgHDcORPBRzkP4lL+uH52PvfRxDtnQz
B5bpEAanG+tCBkK8TK3scMEE3wWhkiFwjQNKDx2unE2XiIjt1lWNxvru63yrSywr
XD32Earu7VWrdhBm1Bi7tTN4XJJ46Mfddq2gLQmFaS0f4wfTclX7F8+jZBQqX+eN
uPsGhu4rAtNMtpzitW2e9GOEdSFjN4kWfldL/wPi0bPTAAR58L29QFx0s7FpAZyP
7a7yqa01l3fY7rQbtbzX+zxC/GvLgTU8K8AhNS6MWrZj78USnsrPKmshS5b4B70Y
oK2CVx4LwhXq/c2YQU8CBMYlB8sVU7RdK59CRNU7dKuqXWObfguLti6OMSqn3FgM
GHVihUgFN/MQc5AjXQn4ho5TKxAOrPLHT7c6BiP1lBso/drCznWEOlS9AHtDUWFB
tXY4BVL2Li/LQvhpFBlc2rtgenM8p/Tog6FJJ4LPr984TDZSqVdU95e+uChdULjt
SAypAFuEyMpQT0JFiYFxU32UWNaN6hMRUBcKhxYAZqrudv4JhBAYPC1EngSskKPZ
zKbbnIJwtAFujhMtbnqaZQDaKhTczeHgGbodV7jAf815npT0IfDB0/FwIGNMJcJ2
0tM1wOMRVDUFDd84WiAImxUGp9l3sY/8+ku8LCaH9FFtlqPxn10+m1Ag3dRTWLTv
gPVrAjPSfJWVpcPUABNKUBNRd9gDv7MWlFMD1v/WjmRLYb9Gwz9970JLm8OJz99m
kPLd4AVunKm5/9wfi2wW03yMa21EiaKDvUUr7mGxV/6b3Ty0JQ2xhKUsuZpb0gQU
yvEO4WJUtENK6mYEkiA0XBqpgziThX4Us/zFtMnJG0R72eYNEnSmstkBkreW34au
yFLbTq+Lrzt7XyR+b2dXae2f42yfD5YeVgeg0tc3dnr+9sml/MjnOCdZUCvaab1J
WjtIxfW3a/0kihVwXTUIHalXlU9t07TXrI2w8wcNYNn4FZJrDVfZgsvHsD8MGPiJ
SnDy/qXzWAmNtCdRFIfFBeZgkWSBJMe57RIqGqGLVC4xe15+ZEgc4uk0ZsKmGfht
W9jtI75fA/NURSUYgmSjNR7fLMuuUEeZSDBNviz1WayLrUTQ624zhdsSOEqfEZuM
4Y2Vg7XsyjhZRJO9MUKLhyK18EymzyEedK3MiA0eCvZCZmSpgk+T951N7xUW6Ncg
Kgvs4UlTiaP3ns/k1QPiEp3bI4a39XfOeEKCqfxOFVbIxtradvULFqmNc6n5LpjC
G6U3sIr1xxuHsZyvkwGh96pYsog+j25YkHhMZR4xy6/KtWBQ9G6V9NO1yY6MRuYj
GGWL8YMrdv7fyROk1vIfbYNFn/w2j1UhXkbYhiiToSfYBdBdZYnKclSghH8SIEtd
liXsOA5c/jDJoZFsLZlTY4EMY27XNPDdq20zBvQbigmwNQ1kR+AA6eMxZzFeI8Yu
vMWUKBipE60gMbovDj5X7yuMj//Z5SY02XsNifJGhSn9sMyBeVnl9kokkFFq6scC
KBTaIVJUR9qOeGfMrLOZwKNL67KAm4tkDwqn47eGks1mGuuwZXphnoZwGOk7gpHk
khfG7svifya9iUYP7A2AzWsVHYuIQGMgvz9olQaTjp4XX6IiQ7o2jatgebFu3Of1
uYLiwlIdQuaNsdguk0UNwHZtZBefzDYKoL+fDDD1ZULo+mk2p6laf68hpB0/bQw0
LwwUl+I+Ggntqm3ZAQ67xNHVpx1S0Vgn5kpYHTQAGQgsTrBFc37LVHBwPAoxVaGP
RJjR2qVlbJQbsVb/jjMVckii4J1ZRJlH7Orjp+N2SGiVGm1+XrtkprPIgsaurUtI
1fBXmuax2tPrE5aasglKE667BB1BbKBU63bcaeB5gUTPTFsudJHiS2vaLKcL0yj3
FXuURPJj2hXbPaBoUTLzQmSfbk9sQPvYOPxom7mKvsViF8jp1TXiiU/AcIffx30C
Go11VsmUAVl2mR/Q+TrqNTGXWzH9MPr5H6cQv2qcQfDBZWn10FZ5XjU1q6yiMBna
SNV63HU/yBLJO8JiM9Kpcv7THPs/sykM49BJ84MotQM++1S4PplU0lSIr9pon/x0
qHBye2QltQJI2JxR0Cz0dQdY9FJLIK6eU0nzl6ThkELMrn1ST/wcPxMM1cHaRoLV
SUwT+Hd2e4/mZ8ioaWfaYe9ooPtQCsIuZaMH8Mi5zCAHzW6vMTwTz17Z9VBGOkZJ
1hplVH1j0mDfX7SmjU66LlZQU4ZV5BirF8D9hBWL7NzGRneTL48/V8wJ3FL5uytw
mK+f0ANC/ZKyzik0i8Vy9g2nGqMYH5sOa5aUbGSwyFpQfOvvAzhPKcQ56g5vvcw4
Znx/dS9r92qK3s9x1bDLOdSzRYLNiBLn2PggijZ6o6BlKc7m6I1DTCWkCSZGr1cQ
EGJC/gIK5q4yhCmpWSIc9EwnAfJFNCcaEYBGuMTUkNsDGVwXwRGd71GrIKJrMnSV
WGBowAzIuPkaUg88jJAPB9WjWDO5DZvibzGfktdutX/Yir0FsVCYpfEr44J6E6WB
OI+BpmhZvX7WXB2n56Wwm+fvSpuUG4hDm18Dh+tlRlfWJQNj18MEGVYuritA1ac8
OR9RgQK/R6Xk26j23+t5GmG0NkYecOwW0C6x+nizODOTWxoSlfYBoIia5YmUldgT
hcP+k9J9d83GVjtc13PcJcFdmqiZYfDPi/WccGcNpaby8Ei3m+UkvRm04Dn55a22
upqyfj5RqzB5PfQtDOIEVgSyJ0RuOJqHlJzbzBjvICTkh07h5eMShAHYGkmSaffL
pasosMC9934f6wJXOSyFGOG5awQKGOVglupCyNO1UaYmw+XuST/eUiiDRXZKhIql
s7Q8bcRpJ98s2XZgUOSBVIKAB+gtqBhYRb9sPQ1tJEl3EOPkmGPPGGh03fFxDQMv
AivB09fcE4mhbY8cM/4W6khunACUmDIeR9xWCb3g6MVRmZUweh4cjdMpefhWJk31
b7YKQhRSWx6hZRXCdw8iDIBOlcOnRyaktwlfPc4VpRP3U8iCHlorQZpnhqJBCOb3
iSe4gujeC9GGAn4mOIStUfzse1kg9ruLqEVrK8fsFWa3RgWNsRsSIcKAcG0nBxI0
PZkWUH1ayu+geITzMqXdA8wSk96+OKW3XlcR4KObrzKrlPIEQqnxUItL1Zo6BU9i
9iZsiJRXXbtBW2EU3JJ678BGO3+m0YPAmbUP8lkfXdmTuHyHEPhRXblriBbRFRAr
EFLOF/fy0qIYavKPBS6Ci2In2tFL+no+UZT50LoeazxHPLSKZxORxMqFv3s/n9G2
4MNvlm7GhskfBB1pqrkYLnE+vk1dMbfiJvfveOSQCc/jdpJrI9bsRSkGpMNl3R3Y
WFo05RYv97TD+lMpqKOaQnf/Oj+XrPhc9AS4qJOkUphQ5QWu5Aeom2b5/wSREG/b
qew4ZwCHzGrtrH4s165dbMVd9wivRPphWsHYPFMc1lRoraLX/V9g8ZSrZ1egmo89
7gollJj4J4oWjYXkP8ug+22kcCuDwDeLTkiJW0MJla0rUzFSTZIT55pvgqMZcY+c
CKCek9Jq9ZpDNO1Y+6BgoLs2eIYdBi0MfXYHGNt3uovrTApHI9n2e7LKHGZKd2fN
X062R304/lyDfZZkj1ZTbfhTizaSV+shydSR3j/rytBbE/dAyAWhvLhJTW7Hb0Mp
h03xBy2UEFKFTmH5sh1Rsd7ISfIBfsfdPPcdmxLPNdk3RLKlxQDeDRn+YNinHcCL
O21isIowVhKIE+/VymXLhH+1G9mK6QepRzCJCJF4+gT0P7sDuHnXv3nFmX+v0C59
LB0Zg4ylkGuTYcuirzyumABUUc7z0qXA23sg46rJWs0TQ46TqfxJF3lDeXqmuJax
HGZ037/YVX3uzhr0MNY6/7TwGaPThxI8LYLsT6JDZKFyuzS8PpsIxMLpyWP5fX1n
kYunrAVE9wfJ3Qf75SVvUAw+NYc2g9TuYlqK2LJsm1MRWNzZJDJurqGn4/8lhrw4
HtXzU1HuCnbzKvNmrzHpieQrjOgyGgQO/MoniYxK/zi+U72zPpbwH9VEZJo/2t0g
N/Uwh/gSHXtq761I3g6RCVv+MIZwudTA58IznBE2Akx0oZk9xQLLbSkx+IC8Kccz
Zay2FzjSECn+icvl2RpITGslPA6K6sRawD/B4docjZoqHpl4GvUnEqbPhR3nhPrZ
YbQ0pYCREijjpg2GkUFv+HCeR59iA8H2JoyC2HMZFmGMITKkOAAMz6MPjQy8I6Nl
Q63c77NWkiXtymoEut4tmUTEKJj9sAG8MEPof/SlFL8necP0HbGHaoW27/WVTwuD
KFTiZ/dzMxvdeLJSNHDya0qrI74g0nmhomAAE+vBUacYS74zlm4PhJWm1YcCqd52
XYD0gNAI5MHIuKkysPXhIlyNgecUDBEQ5dijPQevuJraFO0KK6cCt7Z8kfYRR69X
FYgIXH1uHMWU/6GlNfFTSxSFPuAiu6u7+QBgeFSsfKdl2OVTui4MQlqMnD1LvHy9
c6T9+gf73Otm7ZFlIQtwE/iewQkBt7NROoOrhz+uVDlPjH/MLdRclt4eUOtJzT6z
Z5Stb7LLNQDVBo0WvbUar5lqHBZ+3iPXHOBeT9tksE+nlbDu5q0jWifIOzZVcB92
2JP31ba/wMRcTt5E6l3DIqpU8x+U4XfOWJRSWxGnHERf8lEKSxZX8OylkMov887m
0UUAQn6lmPwpO5gbSnyxCH/mGgaKQ2jqaVl2eftYpKzgn/qvqM8bY4bxsBb5ylD4
L4kFE7XvyS1Y9M7cA1k6HfAhpzzbzzSl1/mLUEaTCKV0tiRYe/xUOha2GvsrMnNU
R1/GnfVGvx/QcusWr43XhjAp7HtntX+5qkopd8Zm7x3ViILZsRnfInNHwBOzB/ay
D0XC15aBI0Tilr2cGmSqvkC/imF8FUqzm0sYnXdinWvbz7SIRZXAP71P09hkU08B
hHUGv9kxi3aLzPv+9kfFWKwq9FScjtdBdHlRQxHU5k4gw6ud9Zcd+TctYv+jg6kn
KTMWwax4gr9qEB2hSzDKw0cXkdmUlzNIuVsh/YvYHnXmvA5Xw7jwrGjvwwrfg9z9
LwVZNsn0LhXZHGWZl+qQy+wt17If0ScWFQOh8YjkhbzQ79poS06TU6Y0FvlcANCd
iTdHj4WAOk6oSmxGBBWbxZ8brrH8rBS5pk3/Q5AYkh5P8h41tDSjAaOODkiuIKFw
amIoEjkGIw0QNLoHldJy52S8ixxizkOejeQyb5yLoYvW48oVXc/sscMjctTmVZml
QZwN86+NNM0G49VtlfGYNw/31XHKLqbIPjzFuYhAMPhbZ+ro4z9y60JOr1bJJ0Rw
XQSaCEBRBgieQQxIrZztPMVxDjAHRkS2gi/+ul6atPMWne+T22pJLprgn9fhI8ty
5APWQYoNHu7OIAdpXbJastntaiEyb5dVg2ForzSJu7oR537T4mOJZUX3OPngkHWB
tpPUIXxvRauOiOqShDxQBPilVRkxQOwY5P4doRkFVdPh/HKQGpaYjFvQ0TUA0/MP
y+6Pp7FSF9J7lGaIqbXTLSFd6v34MsgsLo+Q0OIhgwhOLaHiAgRv9bu+Fpbw+9QQ
uTU7t7uMFOzQXZm4PqoPFkUV7OzlrCDOLnR/HSk1wa+uDkWfOr4Vxmbf5GShE8rg
ubfQ3Z7pSxeF692EvZU8H6KDn6kLf6v25+tYHjwLF20L2QN8Yvs+8HQhucBCDYes
TX7Z4C8Y7/zT8zPFZyQole6wu9QEqoO85wsCZf3+zlUulP7hvJKgUdNQRa2GAZBx
IBgocN0dohYj/kurgVrO7L3WWlcTUanrp1ZvoBYqndLMsp6jNTU0GhG9HgqaSikw
Hvu4e2D1UEirIc42gsOI9mKf2mr1zGULPqzGaZcZ0WHNuN7/JkaU78ygBAmYoW/D
QpgTtTKg4KClnQPnPRI9hqL6Fw/rJVX1aUNslXOU/7mJYZx8SI0HOWcIxcvYu3oo
IVc9ELnG53gdMxgyuzgSZoErYSLuQlnqVqHhIjRWzbJOiTiLFQP9EVGoqmsBcILj
sS0eCBb6eusVRm5cGTC/YCtuvJ373lK0dieIRSoUITdoBeoCPM3iRcav7RKkoJ2o
xzufVWDKr0qLV+QxL2fto+0tdU8ZKb2/0T6u10Vie8/pHEt8IZfsdtVlrlnVoVQ+
GTHLM8EbJ/OW7+a/4v3J5Smf1MrXU2lBlo5aej3vpA7tT234EG/YfNJKYDbgKUy2
m0DkNNA4lVuHi+ttGB2P09L28Z41VRzAfdWINd6P2XH2+s2+TR3ugHLWWBX6uBG5
dLq+K5dzi9ph+XeAAhbEkHqAHPYm515ICujOfR1m4lLT7Z1IAoQujHHRw4cDSbjk
twSQ3fQU6TGf7hjoLWIl3iCb7hv/FV2/fTz91DA/8lMlDS/bSevdHMFafx0qI45u
hxb4OgPlDDHqE4791PEH3WO8tuYnIAg99gKIovYxOftsdJ9Sw6yk9TSBGqvhCLgQ
KfvDDyQ+J3jjjHM09YjZJ0zvDRlB0RwUaw5mPJINxW0tGmeqnNBTfO2XhWEmxrNk
J7Ak6+gV4oafatJQ3/LalDBdQiZnTlNL0tkEUuv8Qu1rY8votIo92AhePUPT/nfM
6D+WZGLiY9TYoO8sc/kONDZBwm93fynaAHSvzj+GvvyvkKmD0Rjur1F69KNEgPf8
bIQjnmHuW2WOzpWr057L9UXf86E9t/PpZBJL3le8Rbcbi8QTaRM/psf+UPTmDUDl
rwhwDzlUJSS4wpwzmD6CwG61YtdcrKXQrs2e1kojklz8E3sAqxUVvo44u/MXxeLO
gVNnLZF+IATwSYffxaDqcjKgHtIvuBgxYnTjyRJRVixo9dJtwQuIy+4EelmxSRuj
uAtVnx2He3nyKB1uZOoaP8YSzJkB+XEudmJPARnvASbMxQaKvL6Myc1SXi+hoJha
OAaY1e6SyOvwMXhWqsY8pm8S42li3ZegV9WYhLzUIf1DOhJ/KsjtWzHQiQS6k2Ma
Z+IEUaoZ67Bx1hGdnltOskodElXSW4Wd/nMweeMWANN9098RJqxhXg3D4A4BAvy+
rpPWo7pEENX0zGNe0BbyVxfDw7dG7Pb52BHt+DNKaKDjnmod/26plIg0hHODoa3Q
xNUvHvOvFBIlb01+baydLCQDhsOXbfQTwevVyBlA9T4SmAr842moQQo/iMUwV3sF
UAUgJZtp6Xqxfk57bXQk5KX1e6oDvltCa0wNDeSGe48JkJSGPOxS0GlbExSfN776
kFPGhFI5Swgy7v8Ez7DQhAhM+URKhUfPgb4v0CEvdyrjpmU9e0uwTG8MiOuG13ed
Gwdkd4R9SFU9vIrfvEH18ASqJgk0DWpwouapJzAdYwlrEIooDuMZ7ovuTECTwAYA
WpcXjGLF/dCy/iImleZo4SofexUc8fCobQQpqv34x44ZkC6Nd6dlj0obe4YrE680
+pUTg/4wSvgj7l5/xEjDGnzG38DgGSEoNKs5zcSeYfMPbjD5U+ROQ0ubxYCQKu8H
LtU8F1X56tJbZOZ7HqmC2lM5gGhIOd2IqC8Amc1Oml/5eFNpHAQyqprAOp5RcuqB
D6Bepgi/q14bj4v2SxBmmz9P0BeQB2Y8mZ+BEnQWKbAmRwOnjT4+b7JQ96sHyIFW
E+2VqWXzz5r4Vdw5VP+ErE5a9Ikh/vjWXXwjGP0roi2zmbljdOT3n1Ef+BVdFgmR
3k8WMTyy5tfzF0GW8ANkmKusUJQms8NvIT/3zvUWiiX1hXma0evKJMv2msIX8E/Q
nU1Wn6ecTwUT6GaTrs4dCvGyWljnzdUu/Qe3JoY7twvGBD6lkLvJMW+EKkWvwapV
9TTWFqzntx/4jxzY7xVQZM+8/EoMZjGAl+2Yx3TjeSKa/oDKKQryoFSp8nFtW0jb
lbYMHoKzilXm6rSE7MVdDnahLSPEsPzYeUnh9nRcgIjlz4URfcNzq/wt/eE3i+nT
cvutBNg5YMhIQdmh3etc63E6MvfdJMLNh41yrtzIZN2yJoYJOxobhASBAMGgaKRo
asmP1fHakK1lhHwlRr6Uu9kltFykpoawzeyeV/thTuJlaYP84adstL0/7B3Cy3kX
c8HGElMxBq7sPa0thV59/9Po7/AALR6WnQY1FqVhai77QZRcEpLyjY5IS4oQZQ/n
dIC5CKmRZEs4zENiWy+GJrcml9hCmqvq+aTdEGXZkM03601ALI3C4Wd4z8H84+bl
JFNUELB9T4fCfc9AnYGD59shvlhIEfv2/hX5TSy6MS3Iqk3TByyL0c3q1KdYky/B
WJf/OH3PjpduhgoA/4XuuUYKuv0OCQnjcJcG76nc+i3Ze8lpXMLwkW8jdzEUtZr0
8TlN1JQETxLdKOFf8OAdKbTiYDDlTYAO1cnA6ZtWFkcKe1/5jGl6nWfd0ziI/I6f
NzInBzHFea3K0RgCjdMpo4DARjFONgmXwde73aD1S9tqJLQHc3s4z22rbq92pYmg
IkMzGQI2jks2pUl1gDwl8b+Lipepvwozga+x7sDwm9onC0Mung/7dbcOZQH6VJ8k
hfTITVEV32CK1JB+CwPpitJMlu2Vf5oD5ONzLONHEJGsTa8VNugFL8HagBr6XqPV
gT3SllCNs9BV332xQ7KWZ/Czoyo9yY4opIpbkoqgFD9MSKRR0rZfowab4CxblrtK
5dkh6/FHWKbz68fSP2Av+gXdbmZslD0EXONVkzWnUPdcK7kqI5vg+7v4QdK8BAvA
jN51UEfddtWXGnBjuKZ3mahPlhEmhUI/QMWWIfQV0/Y71hr+JADZrWZfIgt4lVRB
1n9egqwrQ3DgcYg3rbOt/F88hY0xC0XOfRtwCD1zFKWwjj3dm5tUkUcdzLpPBFGC
vQr+1QwZC7IitzyicJqEa1wajo4ZSn6tnsRFlyh6o5jjLRiV5LOP6A/HpcKc2bJL
1Vwp6osoaZElf8jlJD/wSpTqZb9Hh86rojiDKf4ERikIBrKkKQ6oEiGqhDTiqW+I
qECxIIdLdriRvxKl6cLFV5iWIb3Nf87jljPlbP0Gs07BfEw8oiJGQu0Iq+S07uni
DgyqIL4aSHHgYDK1L/QmSSrwr5f3/7lzmV3SWWJi+VNRWwoszwexOutxUbpCy2nI
oma7EUgBDYtpj3ov8rUtYyGeEs68nZTOKIX9eqTTno02qdC2EWp9XXFxv4RKXRmT
TnqUkhvA0pYWQ5Zf95xHzr33DSZj6WucavphxEJKlDcNkEg7o0ZV/EhOft58NPsI
5Eb/XqNo7q6oqEtX3ZlCRC5etOaRjz6QvnBE2wX9CH+4a9kB5kuNJUy/S0kXTFSM
3O1hCE0Q6yunoV7v6/w1ezBiI472ShSHDd8Hn66tiGHotz1QgqNeOW+eEkwDDyMC
0Hny1Eod8M7UlD8iGr/Txc5czW84+y++p2IPl8J2GhnUn0upbBFAy2uIPuEO+/Tq
4OQ0F0b1RV1wKxXX6DkmmeXzaq25ofCjnlIHpR5uI6q8ll3BzGRmefiXDVn4pY95
vmK87/dBBdMi0O0XmlI+5TMAqT5DhWwYyxVkYOoh3hMOAPvkmY0JvT+vQAjIeGTi
Xs0DZt4GfdoRExvQOVGgGd/3l/f2PrZYQ4betRo+dzMZiXEiA9kQvW/SS479LoqG
6joQHfu1wWFUchxHT9Lu8GZZBaY3VaxaaPi94cj80ea1ABO9yTWzSClLX5Hs6NES
hyAQvqbRo2Eqvud1yIiz5UW5MiTtUrL4r+Ha4uF0CZEDwjEPoANfditGZxxDHuDn
v9lBfqc7838TJT8+X2TRPEzSFNckpw9vpCTChJk/T3026On3OREFxlgZt7Fr6CKr
1uaqMFhKwXEFiG0UJPQhh9X4IIGv2IuZdFZuPUJSHuYM0e912x5Sysi6KlHQa/tH
VoiadEDoNNJ9b9Co5jTZFGBVHs4gPUQ9NC0xNAEia/2I3tQr6x4gt4HXzZeApAKK
v/84EuJfabYDIKb2cVEMRYsNuJwXTYzwuKvVzXEIvAi5vVf2yVze5bE/7RK7h1RA
eyXXcYpI/wyp43DXL4e39D9Ki053pI/B6SyzxGe/P6BZMJZeYXl85hwTRcSU5bhx
it7u20+qLZtCsLm0KNjsj0NrmhPUIbKsE5XLA1qi5k3CAYcKGvUsIs6wQODpb7mo
UtHQ1mimKBqeWa9rgc9OuggqkeZKDobPj6O9iAA3fyWEG9dpD76NNMOoTM5vsgbJ
RG2tKu/AgzAtdt4F7AeQYVNEio4EwP4L5LnjfBk51fTGmkM31WTHgBR2Wuc4o+Iy
9dM3u9obYUrQ2lQsnYiKuojS1yi6nwo9jciPmtcC6JNdxPFHLQRnYQR/g+tNCoa/
L1qKWQkbd6LoD3eDi8zWCZzzN7v+ED+tIhmSg5W9ZB1pg7n7eRFYdAVx6UhkaHkz
OPKqLnJ9gJGqQHumwivvqglJwQThkna328SIg69CzGcOs8iiESXHlrxG1eDrvBxd
xuEQ4fjfyW4ZKzSWmmcjuuLGpbFQxKMz69BjEnuuPHtoob/Ln1IL/gXCYAl5MjmO
lPs+/DVpTHd8lA2PIro76GAQAbk/n/pwpnecF8GGLAB4SORSx9SgvmO7BRAC/HHm
v5yCZrHX8+jbeJBYbm3g69eZFYRESZbypo7hh0SqIwNzvYQoPXswXNQE/nmYW1Hw
p7SWWtRuwUj+hGUxQjXPTY1I6Fd5f0DflOdfsHFeIMgJXaP0fPDA2AqSgnqKLFXY
LtnwghIE1Ntsin5Onmszv04Y2hkh4wYwGih3NVUXLnZ936mTj1ibRrAajlCddMcD
0ysCuwsJ6TEKAXej/LlwkaUSk5MwSET0XH59E4kA+YAW+8vfHYhDv0Je5mVtE+G8
o+ZuYr47b2ipIfL9ZX/ECSBrJIiNk+ghfYezGkdErptIz8mMW/3DRVGkv6lxjl3s
Bxsr7ub7tHTBEk0gNVX5+DyLvBe36cROFalBhuFohZwpqTKoptfIXlmGhuDUaT0m
bIc5uzpemFIWEZl9eR86F3YAnd83EBEQTfpzrEnOehG8s8RQT+azbB0VEPmqSaxB
GsknQFnOio/j4YJCg30XvcYIL7U74rwQ7rfQcNLLpemMZivkD2bo5YxujzeG6dsw
7H4fRBJ1ju4f5YnLmEq1NDDpBRAo/+zrE0Y23WU6XVk0VTkGY+HfACHrv9p3I5RO
kuBYkbRr45WJOTWopoPLqkZSiWr4uqULoVMWmHBe8UB5q8YDalspawo49Ide8UkA
5QHnci4EkUIwFlJe7mCsRL1Bevoi/+1qVXnWEDSIXiu3rok0m3KSiI+XmjcE9kq2
UKuomj8iuTAf54C7OMVhLjm69lghi4gzDio8pp6mJ/uRw8HLuTjzqGUIa/vqdT4t
CJUF6hOAQahQuLf3hVheNS96sIKXNo+CfaM+zZ85L9M2gzHxNJp/II8kGInhKCyq
avcwfvofQFRw0SYyGjagcnFxwLvqwdnGxNE8Ah10SyXxaJGL3Ly8OJYp7RjfNwW8
QWq8AamSyOlpcdhW7JPJaG/+ZpW9BJ8hA1J4IGnbndfMajKQKU1baHmEpt4iBres
q9ajFJvbl8PtIQ/QIp+KuWZuJLB+WIjokL+N2lTUz7Mo3La/LgU9hQzkzzLgE1+6
mVcKjPQHwrpg7na2jR4Dck0fTOUke71UqOApnHV5uGQfqrMyXBTC80tVKMy3GGGe
9kID1gNiQOmPGL8uWHrcui81C5luoxgLa/cc+8zGSD18TnKiuNZV0E19ueLm+/vF
/F34dG5QhfvzCZb9iQ2r6z0Ap2B8CIkHhmddsvLcHJWn/u2nyJqitp7L8F6SalEB
sEEoZY5yXtMrqIZxkht8yig3AjkbGLs2OJ/kobT5ikJf73jrIimaj4LKmrDrKR/h
cdsU8EfZ9ZhOI55p2w2zjtYMiukGH2Zip1i8gvPpfzPq9LnaFwYX9+3TJY2KdpVX
lc/9BmAb2le6y2Yk9lJp9yA3GjdFD4Qe0ElbO08LX+sTr9wJVT0tLUkTme5Xrf78
3J7qjRzHWmVD/cMYt6vtKzuWB4QhLeaiiZ4PvB82AEO34gBry8JgGroSLb60TOqk
r5sOo92jix6Bq70rn9Pg+k7a4faEHNH6jo/OkzvKOJtj8WnTE42dHVD463VHz34s
3Iak5cpZhg7ZgvhF8IVDw8CoAm3Z7AdAhi9SkzoK3OAIiMHKVY/6Kcdrq1sFIGKK
oTI8EV6lk60okcm3hoARUZxzp4ifcqFXfnjOBZkfd5gBKxTZV2J2n/LDURN+eK0E
5Kjqk4VHoQYqwJI/acMpa12KUssaDzPk1W4DNvIRLm0aB9phNOw+jnXUOjnWMkUi
2J4N4HzFDKyAx48UL9Wmmhfr+0BhCySU/wfoEthCQpimV2yJPexH3axeKg8voKS5
q8s3NUZ6p2IOd8Ncv7o+b+lhdRd0fU/nSvy1H8AqYkZvOlx4JQMoA1Hynt5nnamH
VRZC9GWiDSWPFkEiOjRMHQFcvhg3W5+dIcZV5D1ej7o821q9e+RIbUVOCr97zifk
cEskWzBUPqJiHBywxuVdw0p9KMHccV3ALoMfF0UtcRDnrxu/SGb5+/KgPeagkUcD
UOSfSBeXeeWlVazEW+gAtvL661p3Yv6X1nMc34JRGA8ngYeE/c8F5EjIdkwK8Uo5
8duwS3BUGi93wYVx3amEOVaw3X0xXRfhtNCDibjP9eSOHiawQ+biYsXUWVbQE/1q
sAPtzhCqQ0+1UwebI//GhfwXT7VwsHil2Sqb8P/5Z/hi/IvycyTyW7IQwgJ9K03v
qaDUsMJeUzFvpawvNaRkBezbf5PD5LQJ4xTfDHo8I0gGLVf25WIXfAUqYYIq0UXS
lrPCJmKKSRFlhgh0VwBuC9Wpa2FhZ1NduWBK3XDdUbVeEQvLwZ5TSUGFv+B0gmLc
qdeNQJOQIApWLeAXX09KpWCgF6I+hBYrV2qD6KWNcs2cDzTJHaTSmUHPJNJKmTFK
zC+P/7GIoyXY2zwbNnTyRdqpBtVYljNFAE9COBESTHXsSzBGRnc68S7RphJ0KEqh
2T8gvV+SoL62E/Rn14b+4jifcwFz95eaOE2uddEoFwrFfnRaW2nxOIRdTizqukbz
iWpWOg0hvY/mIc5IDfK+3K1hOgtDK5Epe2vkogGOO88xhaUxcHo1aOT7LTvMf6tW
pyMy1DCSBwCif/joYye8Ao2BdTT/+LCFEoBQctU94Q9b0GqA/ah0QLYO3EIggKdd
CVZgwu3ORA+e4yWGEg6F8nyfQUZSsH5Kri06gEC7/NJv5wwtaPIhO5iAZRI9ObAN
tPx6kC6x08i5if/F2IYhcr+9zT7ESdmSZOPbBAciXYw+WhuvAcbaUJwWpZ+OfCab
eTm4ezQ5QnvU9bouKkKC7xPxLD5y3UW7BinWXZa9ngtZBkC/aUeNYMueJ/54dySR
r0yo/uRNRyDqYnHtVha2wa1FyKOlO8aSlwfrnR1pVOk1maaGDrLMGerWxS/xyWg2
mCfRbyq8lCjjUOMk1cyagCMw8yVkEYLxj1vDcYq0jf2wN801EIm88Oh64vpMbUUF
OxyQvxTLthiR3WWT5rXCneYA2venQy67JIFKBOslG/PGVPKiGw6uzk+J0KDPS89d
ElXdCGzuy0aypvlx5yTfemQe8cPB3SEo1tzYKj31ORazNJHBFq1fW8FAtd5qtECD
fX6dEa6JWG+Wn1XmMq02BI/V4cSYb+8/i5JeSiuOxiw3wcaO5HOmjICsd1816wc6
qioSxAqhdUf+mPUh+LXGnf6G3zI5om4y3L2JcId9Zp5T8j41yGUTOhA/6OUHXSqC
3Sa4GLBNTJfJHpBwBGNqnusZ9fjP5l7xP8Gv2eFYjJZNqw71vhOYij0uObm9FdyE
a++aeiTpUa5divNbGTeDg4ztY7hr9s6mRH5It0E54m0tFJsEm4xFX5AkYjoYb7n/
vhWplgWJseHg58VdGku2WjzJKz6YcH6dqLcevbDoaLfo09jgsWV7pvDeiZnOX11E
iyu8JmxLlUpx5gJAE+AugL/6QBuAZFwRdINPmWqbkZ8pfprCiIYA473IR3e+tFRE
fLbKvSFtf9+ZOsCmI+h5oP7Gp/bB1VjmrZe/+ImQO3nrSRkChvlf94G0HoUpiVll
Pmw2lxcgd0ysXrpLD1tLGZki3H85KwS+s5TGbk9Qd0ybBvRB541OI2Fk5XzogDZR
a1dyN3yhzs1rCljrrwRE5flDQZ0YhMCjvFTEbHSRbmidT3hwiNNXoxOkImJA64ma
omO1LL6wk9uNSJutjQ2MgHP9d0AyED2yTDeIjaA/dKpoOiZ8p529JTxx36rwQ5AH
klerkQTM3FRiEI/gJn0JnXddX8QA91uu6remPH/cPld+xaf0FcsFMXRqjQcsPSRV
E62pF7yArXFfmVSGOxHXycrmFcU2NKB1pmY200ycUfkTPvOvoQjtOoSPywQU5ehF
WHZRbe93EZ6FILIPDMlF8BTjQzAXSlzaKPsgFWBnp6rkAlvvhm0fnO79RFy2t+Q6
+Q5dF9LeoZ2GQNCT2scXAvz19Wmz6Y3LQPqZP+OpniSm5ezGaYJzRUlCZ1P3DTqk
7LKODfw6ZRqKzM2LTu1q0DGC48XKTTVvxdjPJOpw+xs5pRZdH8xTBbteTUNWTfHh
AxOwLcrvLQTmCAz9gGa7SgVQ5V90mPcTgePQV2yoy2wTlyTVC5dXtknFIWu0ZS3t
np3NveFLbchTTFm1icCT+daYMxXxJIU8ypoVSv1a/c/KUNM+3H/aEx6w/EoCxHle
fY43/qjbbkPskpc3UTWWMQKbNUl3Wb6NiILTqliqZFTqGNYcTF3wd2Hxapp484iL
DHJ3AD92AdxE0bjdJ4gm2uXd5SIFvbQV5i0DNe14CCtW7wBI4PAREp2Uo+Tan/8H
Nf5SlS3cnshctKocaYkTqh9GzdnMcxMnh2XUhZEN+m4/mo6ogYqSpibFWavId8B4
UDjNWqLYo1aijCPe9i7VDeGOIJiU/Y1hDhd0oPk3e59pw4qHPYKYAFxoVVMlNGGd
l3S5SLE03Xsg/FxZ+6Eg18lAX5CglMRZpajBhdVfYOFugctzmH9ibItnuRiFYvX0
6vuwNij8HHgETVDAFAdCAYRBbrSXl4r9RWvtMEgePSqwRBtzq8TPYvlxhpTze7+l
/OaYuI7PEHwGa7S4+4TB1vpe3KqIZbOPCukK9h2yhTE2DVf4BUWgEuQLOamiZCMo
ZVnZoZbd9YgWBKZe9CrlsKD3iSDb+8SSN+oOvF9xVqvGC5rzcn/KIBlPYubecayK
/xYutjHaWw1AYc2czEOcuv73RJQGP7uVBH/UAfUDUZZVjEEiyOHcSDzhTztKDpPX
l4SO+COhQCLXX5bmiWpY3UA3JGwYqmmKdEmDHbFhvlu3OKiOTtMQNewOPD2DJIoz
tqCRdxBpwuATt55rqT27VXflP64GdGCo/DsEB7gNg20J8j574GNfkcL+lnyMHiGl
sNPiIV235omOxVwZvuxAGFH+6O4IkgjMGoGDX+Ob8Sv6zMHZCzjFkyl1VzAEbddf
NnVwpn86NFkhpFR9+T0gbVcfpMJ1vsitug46uGCg/l1QLtEgx54PVe2mJu7bUhVa
R5iXzlkb7YRkbib4zPifwe/tl2hCz502EcDEoaekZ0vNFQ/TCc5FwmwTRjGO1toO
aLqrQBb3aW7JRj16y4MKpaEOlSVzlfQ/DWvnqoDrToGXAv1KdQfVqJJbdbCcs3h0
BbK+FXzq5jJLsPIxxNSDZs9mw2vZKsoiZSY9cgLgdcxEBhRYSG3ziAQUDLwhWElk
vksBf8gH3Uwqo+msfCBq2BxPvpmVx3v5VYaYr9EsHDOMTAiTB0MkNIKvH47ECLwM
zcxStUwsiRDIskDEifH4f062LkCaS30SACjpnrIvtxsYGX13FjcDx9VzfbxX4H41
MT63XOdQL6l7M6kOwvnq/GkqB+6cbRMXnHON60lkcS0ZVyBqq4RFKnK4FaZugBQl
fa8C+viCa6K4iwHxoUpK8wvFTkwPFLJI2M8MmQnXhHw6RZDRNXRpi/iE64nmCx8I
RoCAGjV7cPAZriYTzsEg5XU0pggsm6u/gndQxQJa87fRVZhPYiHQkI4OqCrLUV3h
j5m4QhIzsEhlhayEbkAQeA==
`pragma protect end_protected
