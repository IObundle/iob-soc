VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_32_128_sky130A
   CLASS BLOCK ;
   SIZE 558.85 BY 435.09 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.52 0.0 129.26 1.93 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  140.42 0.0 141.16 1.93 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  153.51 0.0 154.25 1.93 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.79 0.0 168.53 1.93 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.69 0.0 180.43 1.93 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  193.97 0.0 194.71 1.93 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.06 0.0 207.8 1.93 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  220.15 0.0 220.89 1.93 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  233.24 0.0 233.98 1.93 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  246.33 0.0 247.07 1.93 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.42 0.0 260.16 1.93 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.51 0.0 273.25 1.93 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  285.6 0.0 286.34 1.93 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  298.69 0.0 299.43 1.93 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  311.78 0.0 312.52 1.93 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  324.87 0.0 325.61 1.93 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  337.96 0.0 338.7 1.93 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  352.24 0.0 352.98 1.93 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  364.14 0.0 364.88 1.93 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  377.23 0.0 377.97 1.93 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  390.32 0.0 391.06 1.93 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  404.6 0.0 405.34 1.93 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  416.5 0.0 417.24 1.93 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  429.59 0.0 430.33 1.93 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  443.87 0.0 444.61 1.93 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  455.77 0.0 456.51 1.93 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  470.05 0.0 470.79 1.93 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  481.95 0.0 482.69 1.93 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  495.04 0.0 495.78 1.93 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  509.32 0.0 510.06 1.93 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  521.22 0.0 521.96 1.93 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  535.5 0.0 536.24 1.93 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.43 0.0 116.17 1.93 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 165.41 1.93 166.15 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 167.79 1.93 168.53 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 172.55 1.93 173.29 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 174.93 1.93 175.67 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 180.88 1.93 181.62 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 184.45 1.93 185.19 ;
      END
   END addr0[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 33.32 1.93 34.06 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 36.89 1.93 37.63 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  47.6 0.0 48.34 1.93 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  164.22 0.0 164.96 1.93 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.55 0.0 173.29 1.93 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.88 0.0 181.62 1.93 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  188.02 0.0 188.76 1.93 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  196.35 0.0 197.09 1.93 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.68 0.0 205.42 1.93 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  213.01 0.0 213.75 1.93 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  221.34 0.0 222.08 1.93 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.91 0.0 225.65 1.93 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  236.81 0.0 237.55 1.93 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  245.14 0.0 245.88 1.93 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.28 0.0 253.02 1.93 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  260.61 0.0 261.35 1.93 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.37 0.0 266.11 1.93 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.82 1.93 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.41 0.0 285.15 1.93 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.74 0.0 293.48 1.93 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.5 0.0 298.24 1.93 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 0.0 310.14 1.93 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.54 0.0 317.28 1.93 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  326.06 0.0 326.8 1.93 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  329.63 0.0 330.37 1.93 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  340.34 0.0 341.08 1.93 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  348.67 0.0 349.41 1.93 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  353.43 0.0 354.17 1.93 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  361.76 0.0 362.5 1.93 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  368.9 0.0 369.64 1.93 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  380.8 0.0 381.54 1.93 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  389.13 0.0 389.87 1.93 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  396.27 0.0 397.01 1.93 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  405.79 0.0 406.53 1.93 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  409.36 0.0 410.1 1.93 ;
      END
   END dout0[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  8.33 426.02 552.9 429.14 ;
         LAYER met4 ;
         RECT  8.33 8.33 11.45 429.14 ;
         LAYER met3 ;
         RECT  8.33 8.33 552.9 11.45 ;
         LAYER met4 ;
         RECT  549.78 8.33 552.9 429.14 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  2.38 2.38 558.85 5.5 ;
         LAYER met3 ;
         RECT  2.38 431.97 558.85 435.09 ;
         LAYER met4 ;
         RECT  2.38 2.38 5.5 435.09 ;
         LAYER met4 ;
         RECT  555.73 2.38 558.85 435.09 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  0.91 0.91 557.94 434.18 ;
   LAYER  m2 ;
      RECT  0.91 0.91 557.94 434.18 ;
   LAYER  met3 ;
      RECT  2.83 164.51 557.94 167.05 ;
      RECT  0.91 169.43 2.83 171.65 ;
      RECT  0.91 176.57 2.83 179.98 ;
      RECT  0.91 182.52 2.83 183.55 ;
      RECT  0.91 34.96 2.83 35.99 ;
      RECT  0.91 38.53 2.83 164.51 ;
      RECT  2.83 167.05 7.43 425.12 ;
      RECT  2.83 425.12 7.43 430.04 ;
      RECT  7.43 167.05 553.8 425.12 ;
      RECT  553.8 167.05 557.94 425.12 ;
      RECT  553.8 425.12 557.94 430.04 ;
      RECT  2.83 7.43 7.43 12.35 ;
      RECT  2.83 12.35 7.43 164.51 ;
      RECT  7.43 12.35 553.8 164.51 ;
      RECT  553.8 7.43 557.94 12.35 ;
      RECT  553.8 12.35 557.94 164.51 ;
      RECT  0.91 0.91 1.48 1.48 ;
      RECT  0.91 1.48 1.48 6.4 ;
      RECT  0.91 6.4 1.48 32.42 ;
      RECT  1.48 0.91 2.83 1.48 ;
      RECT  1.48 6.4 2.83 32.42 ;
      RECT  2.83 0.91 7.43 1.48 ;
      RECT  2.83 6.4 7.43 7.43 ;
      RECT  7.43 0.91 553.8 1.48 ;
      RECT  7.43 6.4 553.8 7.43 ;
      RECT  553.8 0.91 557.94 1.48 ;
      RECT  553.8 6.4 557.94 7.43 ;
      RECT  0.91 186.09 1.48 431.07 ;
      RECT  0.91 431.07 1.48 434.18 ;
      RECT  1.48 186.09 2.83 431.07 ;
      RECT  2.83 430.04 7.43 431.07 ;
      RECT  7.43 430.04 553.8 431.07 ;
      RECT  553.8 430.04 557.94 431.07 ;
   LAYER  met4 ;
      RECT  127.92 2.53 129.86 434.18 ;
      RECT  129.86 0.91 139.82 2.53 ;
      RECT  141.76 0.91 152.91 2.53 ;
      RECT  417.84 0.91 428.99 2.53 ;
      RECT  430.93 0.91 443.27 2.53 ;
      RECT  445.21 0.91 455.17 2.53 ;
      RECT  457.11 0.91 469.45 2.53 ;
      RECT  471.39 0.91 481.35 2.53 ;
      RECT  483.29 0.91 494.44 2.53 ;
      RECT  496.38 0.91 508.72 2.53 ;
      RECT  510.66 0.91 520.62 2.53 ;
      RECT  522.56 0.91 534.9 2.53 ;
      RECT  116.77 0.91 127.92 2.53 ;
      RECT  48.94 0.91 114.83 2.53 ;
      RECT  154.85 0.91 163.62 2.53 ;
      RECT  165.56 0.91 167.19 2.53 ;
      RECT  169.13 0.91 171.95 2.53 ;
      RECT  173.89 0.91 179.09 2.53 ;
      RECT  182.22 0.91 187.42 2.53 ;
      RECT  189.36 0.91 193.37 2.53 ;
      RECT  195.31 0.91 195.75 2.53 ;
      RECT  197.69 0.91 204.08 2.53 ;
      RECT  206.02 0.91 206.46 2.53 ;
      RECT  208.4 0.91 212.41 2.53 ;
      RECT  214.35 0.91 219.55 2.53 ;
      RECT  222.68 0.91 224.31 2.53 ;
      RECT  226.25 0.91 232.64 2.53 ;
      RECT  234.58 0.91 236.21 2.53 ;
      RECT  238.15 0.91 244.54 2.53 ;
      RECT  247.67 0.91 251.68 2.53 ;
      RECT  253.62 0.91 258.82 2.53 ;
      RECT  261.95 0.91 264.77 2.53 ;
      RECT  266.71 0.91 271.91 2.53 ;
      RECT  273.85 0.91 275.48 2.53 ;
      RECT  277.42 0.91 283.81 2.53 ;
      RECT  286.94 0.91 292.14 2.53 ;
      RECT  294.08 0.91 296.9 2.53 ;
      RECT  300.03 0.91 308.8 2.53 ;
      RECT  310.74 0.91 311.18 2.53 ;
      RECT  313.12 0.91 315.94 2.53 ;
      RECT  317.88 0.91 324.27 2.53 ;
      RECT  327.4 0.91 329.03 2.53 ;
      RECT  330.97 0.91 337.36 2.53 ;
      RECT  339.3 0.91 339.74 2.53 ;
      RECT  341.68 0.91 348.07 2.53 ;
      RECT  350.01 0.91 351.64 2.53 ;
      RECT  354.77 0.91 361.16 2.53 ;
      RECT  363.1 0.91 363.54 2.53 ;
      RECT  365.48 0.91 368.3 2.53 ;
      RECT  370.24 0.91 376.63 2.53 ;
      RECT  378.57 0.91 380.2 2.53 ;
      RECT  382.14 0.91 388.53 2.53 ;
      RECT  391.66 0.91 395.67 2.53 ;
      RECT  397.61 0.91 404.0 2.53 ;
      RECT  407.13 0.91 408.76 2.53 ;
      RECT  410.7 0.91 415.9 2.53 ;
      RECT  7.73 2.53 12.05 7.73 ;
      RECT  7.73 429.74 12.05 434.18 ;
      RECT  12.05 2.53 127.92 7.73 ;
      RECT  12.05 7.73 127.92 429.74 ;
      RECT  12.05 429.74 127.92 434.18 ;
      RECT  129.86 2.53 549.18 7.73 ;
      RECT  129.86 7.73 549.18 429.74 ;
      RECT  129.86 429.74 549.18 434.18 ;
      RECT  549.18 2.53 553.5 7.73 ;
      RECT  549.18 429.74 553.5 434.18 ;
      RECT  0.91 0.91 1.78 1.78 ;
      RECT  0.91 1.78 1.78 2.53 ;
      RECT  1.78 0.91 6.1 1.78 ;
      RECT  6.1 0.91 47.0 1.78 ;
      RECT  6.1 1.78 47.0 2.53 ;
      RECT  0.91 2.53 1.78 7.73 ;
      RECT  6.1 2.53 7.73 7.73 ;
      RECT  0.91 7.73 1.78 429.74 ;
      RECT  6.1 7.73 7.73 429.74 ;
      RECT  0.91 429.74 1.78 434.18 ;
      RECT  6.1 429.74 7.73 434.18 ;
      RECT  536.84 0.91 555.13 1.78 ;
      RECT  536.84 1.78 555.13 2.53 ;
      RECT  555.13 0.91 557.94 1.78 ;
      RECT  553.5 2.53 555.13 7.73 ;
      RECT  553.5 7.73 555.13 429.74 ;
      RECT  553.5 429.74 555.13 434.18 ;
   END
END    sram_32_128_sky130A
END    LIBRARY
