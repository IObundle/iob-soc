// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rADx5toB5LlGjfW2VNQL+Rj1IKDnafSbZBLiah3GMQZml+Y4NUQkrApZGQI+WJxs
OdwzHe+2Bf/7mPLW+BixarR4mZo0vs9WiQ/ReUISrgfrIPVGvNigjkmzCIqNxU6i
tTORbAgDJhSXfwsEmVq3oYOB7R/toO6/qenH1B9CcqM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 195920)
bp6yR3YfLLPlIl2YM+SS2/MK61w4gFfm6bZ3jrXzztIu+7B+BAajwpV7cYDvC55Q
KoXc6zpjF3x0Ve6Bn7d4qT9LGfhMJxVEjZCvoWn5l5Bv6/zNAxYrioi4GzHvwORl
GMUORbN+aKh+dcjBNHKPYVyL1skdkRet6a6BedAGAyrZXZS5H2uv+QA3lLzLu/w6
MmC5X+XXgv9888x4iDlafZP/qIL1j+jQbDPj5B5m/6kohZUvfrgExTrViuVek+et
+WIPbJQuywgQh8DgVbzC4j0lnGpp8CNa763wpKd5h0aUrum9/Dcp5D7viQ9OgX4h
+cRxVRYBOonXzxpWIXw7ThUbEuYlN8w+BGzxWsV0kmWqqYZrtDWAV0t4ir3nDfnd
RTj6tD/b02E6FWrHC3wX8T1qg+n5fcmXys6yqff8ExVRfpNyAssj7butm9/cs7TQ
laC64PBeywUiueSX61w6q1q+9nF9BMCDTwOyJTsHgGnEiE4eaS1//CgfDrEqqoDI
rB0/tjHKjFvDjlSXuY/uXsbxfgk9PhugOAZXx1OR5UMHygUbNSh5RTC+VmxFqZJu
YXSNIeMqpIljtU2sIuac3kwF94N8BWgvJaboIccQY7Xj2/9PwF4PstdckQRO0Olh
DiUK34fBD2sqYullGAJYQz9pXghue73uNmn0VNZntFBHylxrAJ1j5G/VQ/iT+qcQ
GgDYERbT+A0sw0p8SY3jXD2uYJ6/Gd+en6ReMR9nM+cKQRXDRKLWsKoF+OmtAgSV
FOEqRHvTh7njNuR91Xyw10OA6pGvX9Y2U9Iwug+ZEnGT5fvBbNF6D/QXjF5A/XQ5
n6eI2Mo0dUEf+MrkcE94kI9GCbUTzcIbwJXb65ZlOYTcs+sFUB3eqLxzckTl1AAr
itFf3SBvOWJr+tdl7AuGBIqZjJadADSDtAdxeOVZx+4mU87BE79g/qd+E6+e29ax
c98giEqd4f+PMeGgpsUOTDdo6mq3poKRcWxnBKSZQ4ccZOal2bSReXMaBZ7p4pAD
KAw1rrW6CH+c0IicqGZCrNTYHbXCSZR/dcyzDFDDtwRH1X8tWmZF0cs4Do/j6PNE
gMJWxaW3xiWJbd94Rzrv67MJ/NZ/Q/Omub08QnosmtAXozPJefp7TOaSgnPISpwU
MmRYQn21ZmIzt948/vnrGQ9roon6gDuk42TksNwXUcY/N4G+cy6abh6e+YgYb3Fp
yZ1H8I/jTc0a+B2dik9LWdVMsnIO/fImkaIO3JeKnxvJTdlnDSKU53OwHz9sizwt
KjG9a9ezX2yusN+NurH+Kd58COQtxF6Fxsm5vNVmbTOJJA9yRJmNfYSMkBjCU0k+
EMfqMCMrELYe71B9vDDajrQetPgOX+A6KD0jLj9zAovKffzFpBZm8xh0kbGZ7AJk
eNhQ/yy63nfrJOpMc7Ba/Xy8xONbkGc0xaScuj6juW9ZwQLhfxZztcQzGfXLWQqO
0eFDLT+dC6CcwRwNB8XOQcMcEjpppHoh/Vmh9xiIYdOV5T9zISp6v22WBEoPOSzo
OrfW49U8nZ0ZWFg7kFY+w9hirVL2/wFRaLcx/W7hsB+bMKLhJSSaIwgOTO0RCj4q
dIZ/3d7sjUbk22wrcNeg22pBg7gABTsE4WpAdJeGk8ICCtyjn5ip0sdIGIq8/H/U
rarMbzXj8q4+lHfa/ubY+dKl1VqM/O3UrlmBJ/bNgG9juPHobAbp0OE7WhhpR+GN
abkH3PfYyNrxDQ0szyGXE/JcpfAf7NVm8xHp5YRzMTEmxojck7vnXqjOmFnjgi2n
OYiSuvvhXFMjMMgqn5t/kNl8U3v28vUBNiJN+lKwduxXbRAZW0NpY5MmFtu/3SBo
c4cnhFcM7Xv6amHHPYgQGahbt71fWidPtZylPMFwQKbAh98IByjP3M2ds8hh4KF9
BVswATJ2WbGxRp0FcvR9seTgbDMoB+Wy99fz0AOtLqDrCMoCdyDPv/Ww/6p/9wBz
1oxdkQIuEcGRW89UIJrAcayDObEs23c3QVotDYZmJEnL0S+aqaH64/Y6Pyeonw0B
KVgllyp0tRIhZjga/y2xTfBaGCQuJf4kEWsEUlyY0DN8jbOmgIK+QdNAA4suyDnl
wtqhBAlLVEEyo29IADRyGzS6vRx9iIw0Ns3ZJUszA46tdAi+4OgalGGS0NAHpxPh
6l95eZm2ftlf2rWNwpkEcgKI/E8C2kt5C9wSeaybAGyj8tichn0razHd3kXIvo3J
8RMPmRZQxhwbF9bdTjXEjhRVHLh3+SWRch8KUD7B1UpfDG0PBBQffNQETeKWIe7D
1YZFT6w0sqIj4w5BPVcsHhbuj9Xw5Tqgb+YeKo3M1ir7q4AAG8vh9ZgeoE16b5fY
rrZ9XRbK2MSrPLO/+MS9nFkX6mYH+4iDpf0BAqHvFJYqNaEqrobUFdNQEl1O4mYC
uqMLgXT9rvjkzoUiDAyczY+WvrQ5/n4PLgiBVUyzIhSzS0rHZ99eCISzarE3wOqr
Nl2aQtR0uGKdZjH9+LtAeKjRi17k/KIVkBsLOZTkfiRZBlhuV7aEdV/g1PtobMdi
7tA9IaE+WfFvm+QYvdj4lKnynJacA+LfvkKN3iUJvLTRxs4o/95VkyXfyVv4piwu
CxhwfTNg50zXXoOcB7BPM9pOWxUSA2CPm5mKi3UGTJUNhfIYWFYmxxELezJPfOzw
HDOOycN/zEBWswRCCgDGMC34lB8oGV7l6GAgcnnb7sSoN0/bcqB3W9qsRc7vC9u/
TkUoWkVQ2uyl1fpwqbVz4Xn8FA82mYIej7jzVNlX3QIsSp0Bc+8tOUWgaBCe8S4A
gKNEgXy65K7lGY4rGB0IPuDfZBVrEWbEf6vTiSIkLaWEgdYRslRLrQ+lS4v4rnEI
Ninb7zmNiDZOC92mFkkzyt9ylXJtM47UZr/CTAPPH502mvPvNc3tViMtkTL3eQlC
fqRhNVLGijRQM3ttxvMgqQfZrwUD6okrWTKNnS8wvJbotfCWABOf5qZm7kZUqww5
Oc60wHK+A1nK0U9iq/vv27maNM5dmLAUpXIrk21D2yiPE+M0eK6MOOUZkJDYkHSV
iebTWsnmYu/gZIrwpMR5d2SfYEmrqjGjeyqRMIxalh4YfrYLKUj6SVF0TBkZP26O
ZfnENFisZLreUskcYZ9Pnv9qlW8ons7KFz8hxkvrZNVk900Z3diR34cHFld4/xeX
7W0Rp6qHuCytyQV+V9Mg2XgKKYBttvcD6f8nxnA8ajlmCO3S+06DHE0yn0yahCPN
8bEOQ64hFHYhdi1OkYZdhJFqB45o6bHNDvQGnyKSF/Vg1GiV+kikCPJS3P90POwf
yB32zSZWWYdZrcK5iFR4ZvGotHqWQQEEFtB/sTOW6wwnlhXct+DyPEEqOUNPQwlT
nOKMp/OYL3n2Si8If3xWXHKBr0TcHiZYy2E7uKOxBxssoYYk1J9MP0sct/uUr5/e
NG3oV9syy2P8wqEKgKbPRCRqQEJNiULgvp4I8bVtqEAAmAzoM9ZnVmvoIvywwd1l
Dy2DkP3Oi5dXaJuRTWHzbMV9BzEUk7Ca+LFuXe8zBh2vYkjj+Kk8s0xpYuYnBtsK
MjUiCF5IplTWrxCVixQLgQJr3VgAe4moUfNeaUbWbsH1/LlKuuYjoNqaQKZMdaZZ
05V1MtQr0HMmx5YeSmWC59W3PKWTL6808evytDSqxcTPHq+MWyRt+9+KPfOIi8wJ
XHuSflrtjc3z2wGyizyHS2tedRQJZWdFEr36dP/zGVH3Mtf3YfNPhNN3c65tmaMx
UK/lu+XXN4krtw5JHhj/mEI251pN+prNI+bsxrgyA1LbUEoIblY7qOJVNaA/yn4Z
nZTuvIh3L3/B7O4Q+2J1gW/n0fg6gRStFWaD8PZQRQc+yt+hC0VjS6180V43YQ0W
KROx3TGtDD5vSS6Es+ru352fexv77WWxJLr+ju78QmQMP5ecl9Yhrniu2Qs4mCav
fJU9UfyWKkvTtuxuCWfYCY/9Ia12+akPHZUcWRJKqbiOJ4cB7+g9vcZwC8y7Jnl1
E563hWHaUNVQkOvMTyh5MnIfHtRAbqg5n7+LrqsOkdV0hXXU5Sln6CSeqwZ3tf9U
q+rbWwpYBMlV/KenTIgq75Ls2IuA+zoSOEKSl8sMXVsNFiSxQkmLHmFjPn1K7rD/
Bclra4hIC5/av4Xe2E/U2s8YYzD+CrjuA/oinwaj3dXtf0m0jqSoXnPbld7LhT7r
TEhm5Jf6M8ikkh8751KoXezAOWVpMbDAgw2VKPGFEQeHOrdeab2orUnHR6CheM8X
GHhlXk2/paa4Q7NKCvIPrKlLM7IAt3jWHkiZ68oyUGg48DJtTZq0hibXiDckV0zI
r0MP09j8Nq+MUYYRWUuHe50a7+g0c6H09WxGcmleE1A81c44/+qpT3o21oUTdh6G
xMhG9ITlLXMsqiXBn2sdPXfhTKKQtmO/uORmDo/G0hF+detUIG10IKxeTfiSCD5O
1Ra6PoQCReCHF5bXvypnMN8m8DDQGynKeeTa+qnKP86Dz5q0B/D+tnKgNvfXdFlT
kfjjVmFtOjmw2q+UEem2rp6r36glTzSo+NWymXRgfaArkO9Lwr5nS/int/yr+/KF
KzJApoTXrzU9cicqBC983VKwsVsniGk/Eyt+Q0xjlokeK91hvgeIccbj+qqBKiGK
WU1+PtUkp3bk6DCkIjULA9BnY2c2Tm0pvX51kcaMRnT9/NRSWbBgDYtMEch92RdZ
9Rt2EAwZE/5I6ARQyJq6fTozQC/SHUuasI476daBox6hjOsYrfBJzsLLu/m4DXtr
+Wv8chVjt/OJZJkw4qRj3njFsHWAczRfiKC9lDA+qjAI9GPQKbyFt29un+lsWlb/
snEjHRy5uzR1fwcLq+x3+vEV4pGSQzM3B+NtNR/hk8fN13A9EBeYXz0PzTXfCHAG
KptOm64mPjlB1FyaRhUPog+9cpOAs6y/h4SxARz05NpxDzAcGPXbwvLBhC7pw4RA
mHEuKFKU+LWEt8yES75Z/391jNusmWQSgYmAIxGX3kW+/qZF4sY10+uruFoPNz7a
7PmC6RrQbBtQgwZd2n3SOe8oPvzSw3xliZeju2wTz81oVKB5oW1rfy96QUAWh0EL
RAUstiDAEFKNeR3UbEwwaRJMdfUoVkiWivvTOC8A2NlD18o/mO03vySyqyr7qnjM
JZ5RhwlasgCUkLotrUMCxJNWbwfCXQbju1M1y+zcoxlbYVeheOW9cRFIMB1YvSJw
fVF9zAjQmCcVJW2VsB+TX9DEmxPQEQOHw21ododjCqOICRKvvJhQe9TlBAW+8LIh
0RtbZ2pYacArZ9U5m+PJNSiFEJw3BuqMk8vW2GkCFtIAWK3nVMvSVD092ThMHxDe
op6k6J7c7bwKJSepKJCSDQY7Dym5I6T7D7YHMC3z0wEy1FfwH9zWVLV5rVOGyU2Q
55ccY9mwhV1ywJ0hcLiomso3cJG56qXu9RRoybUuBLzhCAmdc1CFWassZ3pfYKYg
yf2K5op9qYUOQReeCBlNA0ra7PohMCaJDktjbgZYTxVDEp45VRIo/AZExQEbW3Q0
GibGwweHylbtWe1bHQaMyW9xRPAY24ghyuufKg82iVxzgtgZUWbI4etnIyFZNet/
srd0x/GBA7x134mRm0B2bsHlm5+BF/pEpjSxQCQc/VwTGMT3kMpF2H2VzW6iJTrU
0ArIFYn9QcifWoR8AlrlCZJS7Th5Ing11OsjqfNTVqr2cmaxGBmggcL8z9rPWuDV
UrYznPsCkQ0im0jk+tACzrvgSTNHc1MslpS6j817xKckLjNyYMYme2OqxDoyDgf/
N5aSlmO192i5Rg8k7aWdAIeffL/9LLzJO/lrGW61eP+q+vmfSS5hwYLJqJpy87ZU
GC0gewfjFq73FGmhdfc1cp++U3oS4wadTAPvD2BCj+liRR4jBQ5JCkKMGdODGuFM
lXmlKOfjqO9ZQeP3zWxgZBoJ5HVSqEzaxhNe7yZ3Aor7gytApU42AaKwnsvwbu+/
fzPQa1Tv+Yr6803A+N1m7IY1e2dFPbPB5ZF9mE9koTc5PLG+v9BPvTLgJU3Dn2it
lQczyJsKLISYJZBTLqBrnvZ8rhImYcoEVS0324KSMSR/n3Hm9sYy2fBGCW/q8xfR
vrww4SWP1YtB41uHE92Xa6xQZy5AIxNa7Iwj6iq5BZoXy0WecAKDgeyWFtMBH56+
09HBv2oDz0alsuumcvfXe8yfyP8ERAie13NMRQagdvoClbJzIg3fHdHZ1HB5Ui5Q
Zv5wzqssLlqhSdXjanjjomGkfKl8CW9lwTZ6FRWFrwYws5wzpbBjHkRXnDi6CYwp
oAFu1ePISzer2zpHLTGEJBDtUpvLq3+FEVr+Eodzx00WK5ltREFp4QuLa4aoQX2T
g2QATBs9/JwEkoku43NnuIRUlQ3tPV775oybrOb5SCPnB2+sdc2sEBEcLa0r2U/j
G496WB5yKxwT1CPALMTitjOYAi3Nf+zqAWLgZiYusev2zR+yqIzDxooq1EZx1IEp
0+SYIHJdp5exOMQ1Cs2wPPgiqELOI6vppblnTtiS9b5t8E5R5e5M3LP8N2tkf5vV
4sxbqDqBiDUrnt7Tgc7T+OtcVbgyGPrlLiOqM4yXuRKCp//sj7fLfPcFlY29wD4d
Ik1OIb2xpqCdXn1GD1SM2RtcLLzWUQrIMxn32JxurqRYkzpi3s1nrZBHMBw8M8OK
8uf5Ao8+AkAkDTK300rro06L75e1FGMY001vwFFLUOHxKxJR6yLikGtcomCH5P2B
JaASEXnJcpZkKV322tRvw16DIGXT3H2d/gte9FqA9EfzaVm1ubtXO0HjeTceHJAA
3ePUwSZ5zY0nW1UCCuziKfcTSXYsavKmleH8jRn2OOhENfRqr1V4YDHEWUEOOE5V
BiUgutw5BkD5el0yd/ujLj7hiYQlKwT0sWFEpNE2eqlhj0jo2aCU+9olGbZ1jX5W
vxYFZ8a2bu6ncU+IX61Gp+bj9lQNRcCCla8/GfVB3vbefOz3/K/zOfndi5IxzE2A
iAhbDfNzahFW3uReyhs8WUb6eAxyq3cQQC/tiUkfCqJmLsWe0A6Q5TQTIzIOrre+
k2KXNJMQn9l6tXsR+Yb4R+q+WEXJBIh22HNDVsyDewy/laUNEquhfLEv2wunY1hS
dvzXA3sX5NxJl6ejCgk4PoqZ3J7402thttxj14bBO6xjvfd0lSgRTMfLmH1rqypM
pASptS2+TSCUlNasbff9a4PmBJXc33Wjpfl/RZXuQJgj24FnUQTfIaCmEgJKo0pC
koVtvgUUhZIFnmUX7hU+ZMpUvgz95swKNq1UsIRwlnbDwbN1344g0dLpj9U0Tp2N
p8Qtsvgy2AQhL5LxK4RGBShg+Vl97xzbtxGeXMcY1oNb3JsfByQQrSgrzvwjh1u2
twvUp2ciyWKzXgKBN4bBd+LT7T2jVEznY/kl26X8nEGltt6ynEJRJL4bbi5s6FVQ
buTOgD4ThWsfJJmo8LPM8ktZLkEaIiOngw6zFrQb2ew1EtoB55r+/W665i2GmtQj
kZSah0AJ8f/NKMNr7hMomRhrhFOUczcm8UB/Y0xqgPQ/d1K/fI/99+pZb6H8sV2U
o2kLe39vWAKJmtdtmt0mtud/JldilLXCnPewqC8HzcG4aA7FX3RDN1KcA9+RAnb3
vijmuWFILf0ca7wz+HVFVDJA08HTVAbREU7bDdCFHfJhXVNi0mplGJGXg3SmATO3
GMVB4PNlmLRnwT/O3VZZDzs+bxVCXkVEDc9RJ+tEktHXAqXPZHDJkJ5ybwWt4G1m
4eGMxAOanHp/xeSLPmE8g1eueHWvHKPi+IBqH7O919n3qOnphi++B1GfiR/8CYD7
uevB/HClTlwSpa9YhHN/tdNhW4c4QhBm2uEcvS7b9KfngxOU05FyM9jKBdornq2y
avLKWc1uY93gogl0MxAA2OD6HV478Kw9xomt5J3rSpHkOFjYCOwZXe3i6RfjG5UH
tgBuBPTbj28kCwgTJLPSVbk1Pomr/Sl0mY7nE8CHiWpLHkqcIYfdizlIiVfvhnbz
up2XeqCPghH8sDRVexhBvx3xr7VAy+ygZGPMOuni+R4Wi3wCyZoNddaXe67geGbW
Kcp7aJDim3+ydWCjzuPsfWUPN5W1ysRiEoZ6Ss8gYVHDM6g5ZVOn0wMuh1MF2Hzr
4HdyyORH9PgoOgVR+nlrrQ0+E9q5AMuKlhTmkaF69JE2jrTbaiSMbiF5yKsOp0X/
QF2HnbEzA+172uftpJ5xb1tvz1MrmlYw1r4wNpuHmKu4sNMjHJoWZo+zgWq9i/kz
NbunIBvbqusQ9Pzw4HIg4ClFU5gCZE7tIy5JdeobwOUiQdIu0Dlq9UdnivDSO8km
HLOuXvZBMRr1Rq7XMe5DX+Bpq7WV+igUyvoaOkzRWGMJk+tcadGLEGUyKrI6ZDbx
ZH2kOQEHZJVhjH7t7UbuITIHjZE1kCrtYNIKjTM1mSWs8Cgs3lRp1qg/hVGOq5s1
Epxoead/BrFvXChM5SumT/1nLYpTvdv3o0F9oNGJMVYDiUCfJ3m+rm8NPVv50m26
mebz5V+t4ZNzj7JuaYeVVyWdGKrk5uZQi3oKp8L1jHyN3iZPzDGz80MiwJ1LbDCB
IzNcTAG7VpBTGNhj5PwAO1rervt6j5VC6rF7OaDUx6LxQJpHMD2s4H0RhmxqiPcf
gKaAxA6O9BWBWQDSu12qXNEi2ymPRQSr9gHQk3XiPBY4UKg9yud5mEEeCfLDpBbu
hDqQ39lgytutUIqLs5Qi6m1DiPHS1Y7kCpg9S7FeYO5p+kTZu3x4GjlR6lvcHFkr
Z/2mkIQi+gxOoGnqpZ7PsnaCILEEYi20GBpl27WVWOfPkJiycXqi4wjsMSWwhA7V
gcps69NT22jPErJgbsQtpAgcnI6+uAPT/S4w5EfKeht9/z9Fc4bybF7j4xmZMZ1P
uLfg8jR9yM5S6xDTS9yL2LTrUItO2O8UV/3l+2xzrOV8QbTcDez4V7RKbhCv2Azs
VkYqnt5VSjohEhnJZg1Ns/7xVVs/yx3HeCIKRCjO2lWaNrxg+ABCq5ixlEo9I+f4
W618l7yMZS0+bdTTWhLa8DCxoJ/T2fNgxooGnMD1NSMUdsfWdHDZqBxtqwt1x6Ul
fGqIMbSoK0jWSniu+7yuZewvx4EYPujZUHIv857yJGN+LIIQVjN5Off3ApKqiNOf
PHA8fM9Kg8T9GntEqgJ0nGYxX9IbXYQXkYium5eRvnkiu63O5r0zMkQr/RntbSuG
1KQjf4ptc5z0nbP46CL/LT7mIxQ8ku+BeW1tkVdpZOgn7A+bm6sPCwmMdVePuIf0
YG5MADE9pBec587n/aJtupszGtR/y3AM9mGPzN9suuYLxID+8mk9yvl27E30wpVy
Y1yHdklBlEtLFuJK2FiCtSCHMAOkzs9c8MZL7c1JuP64ETiHZawSzkV0moQy9y24
NUAOF6xMCMqhmdBHFr0KCiCK7WONpRDFsNC37M8IZAX1lZmAkHAnL26VxDE9FbSZ
GAvdLOmzg4kqr1U6tg312sFe+EmECBN6W3bdBgp6xP22Pp0XVhkSfeeqIwq3g4zN
CPPowmFH+QwLO41+4WZd1qE4yNYgU7eP3AAYPI0YnxkMu6X5XkYei/FZ1S0kyWmD
cCtvJhm9siNCWsZhT0MGTxfRcx5XB/hHw0dggu36SH7tneDCI1zJStxYjEWr6t4P
M7ft5yZRi/BXLAWlFs0b6rEb7y6k4PjEyCNcaOBEQNOd3/TAsldhzxmugHnBm0Kb
Bgud6dQZi3HDD0ltde9I6ySTWmV16mWWlqbdsLbz/yXs6N5AdSvPV3vUNBgiTP/c
6VUsXLPpru7/KvcD6wo5MmLd8RRpNjoiH8k2oUD1CrAdSI8Gr2vSKwiIbb58J9vT
S1kNs6VnctkZp0Ld7iOjPFaizM99NEBt1LHXA+CuaiHdMGEX/CmDzDIUI3vfh50q
1FtdMcimY6zeYH1W0i91SpLWcZDRpsKhnvi8LFUwWFjZpgJtLlp/OSlLmasMjjEk
rBMfANhd7GGHVLy4ya/YAcQ8CoE4G1PhCAxkh9RGPgtUquY/nixMbIu328IQWJzw
DbiZbcyTL+9Y++oU+BqQYbDkreSH6kzj7yed/yo9il+BRuS/5geZuQQAyXHPLY8I
ME0T3IK15SIqt7y5WT+qB88fbhEszyYPDP3Kl2SuNitxqLT9Tiu2+qhhied6Ebu3
A8S23aU0au6pULv5omTGAu68/T+1CXL5zvwbItd1oFzC24yeH3aGV2Nqjj1UTorV
ZA7yxSUeu6c7oiU4eWeVdNnQygK7rRXuksWBsON0mlmK2YVzXEgGBl3Ivin+UXeT
YdZudjYz/EcX1dlMMve5ggojDEXVBprd1TGiwCIYCAOyMW/uSDZVai+TD+tZqLAO
KG9jOm2+6pq1Pcmq2n7+GziOGsZtfB4iQdWq9XJKZ4S/JpJwCzYRDg5t6SO8D/KU
2YK0qQgPlqRXlWHOtr1jqjv3D+CVvn/rUXRbRX/fJMDVFO8PzRYIldSr4qZcmMaA
W21Wsy+sDer5rwXFOE/1lTk7P1BEnPsxbMrTOp5Nq7AEBwlh67ZmfrwN5fjJq6lu
HgA8VtYWFlfjxf4Xf7i9fVrMOzGeEjT9QHm7PY5Szfv1QPt3l1UtIjmC5sd3SIo9
sAbZqBMzPT5RJPJNjgU0OBp8Razzg6UL6GzG6C3i7/5OZ8ZpofuYKc9/duFKHNiU
5npgALa6RBx4Y2l0BeTbDR9xWA7yJt9Vy3GmKzg0Yodsvrw0IsgQNVVCVIt1hzsK
QSxB4N9CsONf5xI4w8ByIEYjBFaVPn0Aj+41ntJ3wXMjglraRry9OT38QmsOsk7P
j/NW1nqeYS2GJdG72n1KjTZ6GlwQKXS4kAd/vRndPCqH09AK9wrWTFvyTMDcWGWP
f9M1xG8KJJbjwF5xX1MDhesAlZWRlIjzVVOU5CLJAIJ5dZsHNxCJVPExoEru5Cb9
lqKbKdt/LI7oxZGzMG2Nh5gXsePHQcc5A3bvx7wY3r8JcTwAYNwvw6YFJ7pOBsSq
j0VV2B4pzcVy7vmJeiLiT7ed9G6W4eCMdLHcnwUBzAYMBNuPMQ5Vn/swvRrPzusV
uUunjd8T0JK4U8z5dg+yGybIB7ypNrraTqrObDApsZlETmguHZwLa3yNkVct6WRw
wmk6VAM4w03aPxdhZRbMBaMChaDmpjePiRjklT9iUBE4jasZtIogNQEEyeV+LIsD
UCIOnutbnzlHImYmJgGJsv+YYHwIb4qkkrK609Nf5Q9ASosN7MKl60jEBpgSF7vs
/TkSa5qRtt2m4IWyWcRLWIhVJNSZzppgxng91OQ92YgLKAPcNS3GZDggtBJ1ypBR
TKn84Vnkw458iLur7IyiICfiovlKd5rxe3WH7Q1zd4OH6j08JX109kN/Kr96Dmh1
EKqIjf3fkLbhaWMNgACvhsifY4aEEArUdnawcSkXGdCofcVl+4ZvYw/K/F3hbqcX
q5IrKxMnn5eyXI0lGDlFgPrRZhHYixuG69USymjaZ8B3qaFLJmVaK+T+DA9REUZv
vhQjxkTz+jb+oDi/BX7L953ev5RQBo8yFeXPfGw6hZfsfIdD9YHMwCVFUZhxr9Qf
vTCrFk2+IK4yqbioCNYoU1CUrqme3Nw2IlmFLUDmY5c6ZsHQVfYuT6oCFh5XcwZs
sBw5nMvrzJXUfk1v1XQbuFb4zkVYYusQbVQtUFioxVP1kDqTCtK0OoeUCKyGxoNA
dYy3oNIv9iaxFstlWF00kKbuXfVVmbq8gBGc2JeqONCdDJb693/E1VLyq4UKHSBf
/DMJTNqvWuz1Jplu+/6Lo6qlasqirX5clxsV17t45Fz+0tLtknm2/wpei6wtwmEH
hFxRIlo5qmicOBZnRXZSGs7qFcresRXZLzCyA8sqYTJxsvnEopKpekMMgpm6zpYm
5n+7oS8QhIlUndug28ZqHeCDpF4pcKmXyasmAaVTduqiJv8jtEZoU3AWJWmbW9gC
cDo/iesKuCFT7DBFc3sxwgZukrbuZVLuzYQQOOGmfolZsjXcxGH8jKIc3DvYEuV3
MBzI5WKZBsiPI0lKMcbOE/XJ1deWtOM3mAKSwd2dXuH/8AL3lgcO1df4abxExWAV
Evgb8MHcqKFJG9fisB5X+f463OXa3kB/nEzx4cs7cFzSUHxpeh/CTzUS9Hwz5PxW
KPs+l6Q23LnbHec7wE375WQrJqS8vv5Z3UIgNqpnKLAwFoTKgpOU/2wI0d+hFZ0p
+kb19RbhtFbezqF6ogUlzTdVzhcJ+KeZXlN6lxOOyN1J10kxgZqWpP7sSuT/47Je
wPMCX6ktKTczEDDD+0PXH6DyocQepKZqgaLkpQwiOlHaFmcIy0RPDugeccc9qVkm
yXOtOi4TxWZv9y12CkiZo58HqSOPK8WH2EAsE0sGkO7rIGP7nV/xgGhnRn4l9+4S
EKJrriRGyGtcoaAQMKJSvim8Mrr/jGJ+2zucNd+1DCBeVaOwIQqyJNGblF2YYlP1
wUYNfJXFsNqDonIO+tJFmGvODMRcf3a6mYOT3KZPONTHOzlF2xONhn5QtomAA75+
aIGVFwHEsHd7ol33EkUIL7JIf+S3EEjp7ULUq5Q8nZV+gAspzusBZ9An7rPkfcZG
xHJweD0TSs8rX2gWcvKSTpq0Q/SLbwa9IzNxV7yZjCOlHnKGyyc2i2daSML9ZRho
wEhEZfmWcqkzj1b3dILfva+kGpS+U1rI3QDJH6SvCNZl58+auqYQhfDtfJj73EOR
70dKVNYJ3PvhNPIqs2yhgblqje+59x5+fN7TSA+9NF47pdFGGd4wQKEdi14lmbVa
2HFwoXspOrTkMM1f8+eQpYvZB1r8makvhRALEKGIrxvxkTi7FSVtUbqRkGilLr3U
K+gFPti7iUxu5fc2URhIyBPWu+IcLCU0hGqXdacuyFNgaekfbhG1HvrDLfCz6uNb
f0aLwcvxwkKl0rVJdQMTmNU9bgoSYOqqP22fLs7BFVsdpM0VVkPW9PDXSnTfOSS+
qAlSdwRc95Y1XMVqosdN3HUkqCW5wAHIabTikDl6OZx0Hu2Ql0T8LWlVXa7OxZr4
tlvjgQ+W92nPaLAiBgWuqdBE170NHvmnWMxgv+2KGReWQ9L+2Qvv+TUKFeDzjwgp
ZQvWc6JBaUm1CVhPYXAbeKIOuP40FSy+FJR/3ggg+URGGDgPEIpN15ANeeclNeAU
Co2FwdsaGfv4vX+kZ751EwK0jr4CHIYyxeVAh6ZjYeCj00j2pAYeEdFKQVeBlFSB
eZVSg1/6xMjKg6O7gRdWD2hE2jiUffvoSCt8aflh3FQ6Ui4cdUgfj2cb+YSS0oOX
JLd3LAUcljgyq3JlPn0IrDJgQEGB/w3ZCQJkE/L/Dkyaj3cnUaL/IGyITn4dLcK8
9zv6GET2n8XFv4hKdrgdAZ3qXqpZyeEBM2XwR+HHx6vzzGTNVXKf1lz/GJcaVJz8
11myMS5lXe3pX3YLWHCAWZ71uvu4SBb3P9/ONbgUR+keAyoF9PsYllLdqDBAHmDD
s+2x6rp/FgO8zsdkUNo69MzYYNFmLFccOZgw7jnaNyeYHNj8s2YXU7uJspZJ56XM
9cOgm+y/ei+hdSkSUsZD/xPvlxjx0IbL+9DN7tWdYWl2h5Gv5r/8q3ECycWRumbk
HOXgp13uXh+90n57yqVqu+t0eW58boOWFwxzJCNojrHaWTCmQejPFPSDrcMPEH/x
K/mNA+aliOeF7kGrXILJ8rB/rSxWeGN2bhp+iUYXEnQpNPtEmYlqWoBOEEMc96p5
sVSHPN0b6la0BfIm8OnxcVJ0JWGXE5ctT2owNbpz0uDJzKiOiPkwWUBVvyeQ61xC
iSONq+186k7r+vle0b25dI6XNV4Hc/PErqlPuPGv4WNK8H9KEfIlSiOxnOMxwfqp
L63AuPeLe3h0pdNwhU3qZ7KpPFo4sMNE9vfwQsW6aSVR2huF/RqwDqD3pkGvyF7E
D4+IvLlnLQXPwKEB8cqw45X5w9n2qkyvRYgu++jhF5AxjS5BipkFZb35kzhOLwo8
+Wadurc9N87TILVRUVBSY1OwkuGKbC1TZn04EJ3IJZ5dsrL1pVXDNTyX4NpxCS1i
Gr04roLD3PdMG7xay/afTwNmz5QmiaYLgZ0hPRzfwrwka82iUq1TJuQqKAvoS1k6
Bf2HwWwlpnt9G6D2f5hvwvig5GKJY7IPPOw2lNm6/qvJkfnLrsB2vG4Yo3HlN7Nc
kN0WK8EO7ozRLB9QKsRu18FXjlhIVnLYgbxOqW892ktOUqslp44rileWhpey8Ei9
mIcdlK/dr14GWZ29fTIIEKCRhtOW8+4JFZi7ycWj+dhqFN0eGyWRC2gGHR54w5sS
S/A/2ERaJh0L2fUwdxcL1dE+4pxaXc55BLyymfnBxRVSRx3cFry21jv2+6Q8+a7W
XbGdyaKvINVwP9d7xysin7hH/fR9/KDFJSJLlnX6zL8fQXCD7IAoTQA7itLSdbPB
lFccwv2crGGcr28MC5LrgFRLH3jGh6kf3WPL5K7QNml8q44N2sAHL/QrjZBM+lbk
WvvkyKG9xul8wK7MkwjTtf/eAZbHg9AJNlMaQisnXG4mpLCB9bKVAp+kbNycW8Lx
FqwLQx8XdsPheDwruNtOtVbdMH92GR2XKWKfH5+wd0mcLzbbZbxyOXlrZo4KPwCo
fpdnmYiVClmApI2jJO/RxMRh/8A4cjpDZJTJU7EvP1oiIPphW9PGgK8DHYEKQTWt
8qmNogHQGIqw6NCyMYmLtgO2rzA18eoMgN2x1lbsThFGbQW78+WMvVSTF+8qHuKv
+XeksV5NcnrD5DI9ioDgcldmGy1R3fe95riRr1/UucEYrLxCf0TYbsjap4mdCX8H
/N+R+5l/fX2d3i1beHMKgGYktpIK1IaMoq5oGmaVcMIv2AUJrzZFKkqefj9xdmmH
Alvd3S8MYN0nGAezSW3sIsk8ami6go4o2Vb8wFOECFKsRlRzklP4/MBrjPbQjXVR
itZXJiOU3CD6/Dzi6vt6fpZMlO5OJ6xJjYOT1YhQCOlVHGSbJDkNouH/Yq34QUwh
yswkjOtha+rTfx+lQbGj4ljGqrg6BAycFqtyx0slJWltdEWvN87FIXYr+ZqKSl3a
fe0knDjNXWsluRSaWNn8sW86XMdjk8qNYm3bNGe05NnLZ8h1IeZfoaCHXqE4X2cn
5fqhaAmPw1/vXDeJTO8we2E/zuiBvJXH8GFjdUKDm9KffI6SC4VADiGBqvl1Pk2g
rfjuSrxKFRRLuslhl2re+sCI4l2J81gTSUbM0bp55qE+y6bNQHnIXMBjL6W8EcMH
K5o7FhHXDrLAZel/3oIfQSEzd5Dp8Afs0XwYTxxGjVGwJML+lWBuZgTtGcwTu1OB
zNns4LzP514YjM+5wfrIKEF5hc/njWZbTMXMr0vL4MGlhOg7FmI6AlEuiZkGP1H2
Cr6DEBinbLJwFIbUKgw1s2cYmHf/ICVKpP8Xx+1u0SAVeIrsTZ2dA1fQFj1JYKht
t9bf59L1hSpXXueMWTVVYt0Nll8iR9uIC3cvyh3ik7FFHeyywVRZYwiksQ1kFJNJ
RxDgcF5UUypVza99GxUKpGGJLKsrJOviY0roALTuBoIMhfmVZw9C6XVzGvs5su23
c+leIyycF6Q5NbZaqFAscRm5qABpsskMU9T+I+aJ8PoufjqLzzVtuwQokY4im1iv
m9PCsoxNLhzEMH8aFM5qJCXvSZoSI3ixZqJg4t9er+SyHhoPIB2Vnq6D0ztZMDgE
jTdTRM0t4Qhxr8y59qVPsofBVjLj0ncsuiPtf1Q8W5eiaOVaW53I90bFd/VT6TWT
SnLYUY0tbOQ/tWxTBo4bgRlCpGgawXovBYT0eUSw/OIWHsAoKmXUg7k1hHa7gpC0
5nqmy+QU/BmbYkiqY3vFsPEXyWh+4qusROlOwf1qpm/ah8b0OjXDR6jORg2eFFgY
cA8och6ZIHEEcbayl9rZx6Ad10e75oWRNNDuCZJar0Fab1M0sjd7tkGbrcJJrkPU
TaGfiAKXwzRSt7m+i8UKvVQm6khd6KLIZTtgbCA5yDlSVLlVYLAoim6W98Izfss6
3YeK8ngGX0PM/i6Qm+LVK1tdPVt6bs335vFwHLynvlz/99FrTo/3daFANpKC+w12
hpdGuLYJWtQZksjbmKQHnlsq0oW+y6H11nghFkchExpQgJ9N/SZsI8PO6CjRcb7T
oXnpxb00NeZwzmt5jG1XOna9JjygDwKTWvmHg1piHYcKSFnS6YW+h08AdMzihgn4
bfKdNCipEmAAxCLEmYFFPeQTHe1dFiWMYmL0cQ92p8m1douHZBL+VwacfsvNWmm4
iohYdXm3S4H0bmfHh2TAJqWEFWtYoSEIgR9JUrCbZVUYO4pcfbAZWFA7obazDpfk
qr7JidpM4XuYy9+nHwMZ/Gdu5thDSZsr1L51k6dR6WtPM5kCd4VU0TRpfrxY8NFv
nAn3UCN9n2EzF2aq6hBpPnbxo+4p2BmxyCifTBYQtx7587VZ+35aOJD4A+iW5BmP
7MwhZNe5KoevzwXQ5y0ApCogXEb/1KqjUaifb7CdAsDm5N9/SxrIA5ek0prl9RR3
gIGfFh0KqjmvoXnmEIE3lzgcllIBMnHgRsmJzSZs9mtOS0v/KcRAkZfqS1DGi6qe
saOiiyThqbNoowXiU3IyK3LlxMexOQ3v9jopPJJaVU7W0oo8ys/+4FQsHB2m1JUt
/aV8yAtL8XzpmD70/hwfsudfcNL5yqU0qxdON6e6C9QgnuGK+ge5LQHKbztZF46J
RR98X3NVhyxHYOjYQXjeJ+bOYFaFl0ROdeydY7XQYrlrfHYqRYkOnwO6rH+SaYOT
en3NemMa/gHi3QSBXJhziWoUkMu/d3A9pzGYjjjm6SR2hI2otCZrZwSRn8u2b3KQ
eaRvQzHrOJJRBdKU1OEIedAkbltqRLHLqEgBqQ+QQAGWOK0ssUHM6jVMcdTU/WdK
YmTP3HggjXL81Su06N1ucScu643e+hdyySedr7ZpHXPscmFM1L22tgJfjrDIl4qV
/m5x0WSm5kmEA4IvEFOVivhCKbGMyLozP+htuObg6lrh1qYwlyo8FT2RobSGwOeq
QUXJqEpYdV8+H1BE3cLDN3bhHHX7+x3Qx1thsCF1lj1SGg+ngL4JtJdXuiTORLMF
az5mRWifsV3GuopnKyDAXonuacfA6MmrVyo5lpOcK2YPF28T6DArfPcb8gpB95ay
4VeRUQwtIwpnw5KQ0ZUWo2cjEaSP/JImRxSYfbP1XuZLLkvWI3zgLDksS4KhkzYL
N703t0iVDwmYaPzg8Zatq1xb4UL6dEeMtOB6W89sbB9enc0S1xzQ2eMQjc4HsYeE
tFJtZXYqPLAZNhxtkT+1CV8gcNivhAMi0veu2HIm5ILaf5nSgSNxLGpuU4reEaVp
JbteQQoA92e+3SJuREnYGnIa+d6swTBF3HyJ3ghWKuReT3BmINpmZPEYHaNs70au
Jwo2lrkp1N8s8vJxKegNj6/7jzr+hL5EP/OzMGa/fU5GwsYPRIe7F8p00Onw3STR
agya0qJSwlRnuD4I8A3MCtkZmInGLYh8ymWZKa982RbF5JEp2LbyFgvglgItlfap
vbQxDs639kI6TRic6vgqVKNDLzbUP8f9HYsXK+1QSw2XOm2DDPOt6h5Fmt3n56ol
23SpCVS8Lxtaub9jAZUJ15nRGWtiUDvtyMuAwAXSQ/UtGB8isjZ8gs6NCLwkrVj8
/MZ/oqT/cQXpDhu6xwKM7+okHPQHTPr5nrBedoalQQ73ZYgpOECPKRix5FZdEiUL
WGtbn79uVogc/lkF688M0joQ0mLD9+YCCwWHxkctysnrRYJtbnK7cthIpb9vjcQj
QJSHBYMFHKtYfVK5z1ibTl1cYih0kZnPATvRKS5pjK8oXWrErEbuqoDRdQYzjV0k
Ib3/v8Qz+RKTEMUnquVUq83CNrYfWOeuvAcygLmgs8IPzlNMcQ880Txl/OONaTs5
+2Z/X5c/+Njia5dwYdR9oLe2egmVjFb/i991NFcOSVfxQyXJuR/9ZOBhn0WNcTOZ
38AfDN8ijwZTa3nijN94hVK0SvVC1SH9uOsZADRh24SkV7h8jKlTDD2H0IVoL9ae
5qcbuXAXY0677C3SqhcLeapTYqieKCpP66Lq6gpPSy7aaRKGo14BtrO0y1KO2N2/
BloSxsrH3ardXIhhJKSWMnkO8/WsQ6I456WSllihFL5b5isL0ZqFZoONrwyhoyuT
fKPBDKWjDowGCPpe+C+cUPaKh9/dGQ4UXS4CBlrR1HoSaLJk/m9auGalcqmvwbL2
xhoyFako3dcy4oqgeIEo3lxyMkB/muVzD8gSheUSYiD/+jQO1lmnm6WdLnYGDfzP
GOFeagZnPzsh7KgX2DP/YezS6EhsjZK5WPJvGAwr8rw+L8z7+5cl8sOU+jNTrxal
hR/c6mBDJCrw7z7EPv9yKuuavfg7IxKKAAs1q62unaacRKi1stXW+QwcXr9EKgyi
OxMh7fL1a915R9KWTsHHqMHOAQ1zYOsvlHk2DQ+Gd837g6OoQNYCiY8Z2vSabntO
Gpgp+fjV5wTG4pPeQrom2mFYiYsqYnXrBbxW5Fua8o8UcJHkOBzTYldEjyN04ouA
EYnhQ5jeJR8+o4YTzSOZklYnSGUGLyFESf+KgohZ2oxEKH03yZYXVUuS+Dp7utwB
oPB74f2YKx89exZnzvp8bSFOCSbjUHI/Umf5DprgM13aFHrHJKTncoLddUZ10l85
K4d7ngCJjo3h2pNA4wGOQztgeuLKSJeah7jhyThTAv8hyZ303cOKOGaq/9PKg6m9
r5EkXcVbRHC/mA+BOf2tL4/r7V5vLOa6ZifyW0an1JvazzMhYbiCGBeiAVvICzS5
yNgAkOWK25kNjIav/xHXUwXGHQOxfNtyxx7c2dqggiqMW02BkD251mutqmBT4uv1
VaHFD6ygaJ8fA5aNEegoxb8ZdyT78pL/68oC5LfSwKLXrV808lgqwdyqiZGL68bK
hFMj22ephYWNHap8tyjeCkpQ2PjR7T53BU5XUgapjG2tjM2/jwS7e/5cDWGFGzUm
q9wGwBYR8S4gE5kL9cGlOTn/SJ6mKhaT6zj/RYpIVjA1TCa+wmK13D8TP0cFTdJ9
6Y+LykCeR5wYUcIbPvNX2sqXQsXEZX33w8Qa0kHRP1cCXdnrcTWfnlxK0tJg5Rhd
+dwzWAODOdf6jVr5bIBDXU+tiJdIJdYKlKFXhRwZkBWCAjDeozCsBiQxIAxjqZ09
a5vb6QmRd6T2lg21ROoFsFrrkXuwzYMBZf4wxmdM9sALrC2L0oTBCwjKOi1EjWDl
TRVzIDKCO5FxFUAONWAhZrsg7JcSFN0BRrL79pCIN0ur9hBwCI/si+68iab81YtS
+TGH4o7GDkxWWPVDhB+5Zx6b5TB42aeg240O2c+2fxvEZaHSQ95XJYbvHLxicz3L
/87haZUDzP4gUGpLbyBex2RMOTxQ6L2lunYcaPWxXrWEXYslDJiqKo1h46RshPq0
P1mQlkCorm2VBGqfLONnO9Q0bbnmRc7C5Iw/qjErWd32qDs+zPcqsIA7RveeaPoH
qvpVzggjzryTQTyl9F8JbiKji5lU2DwDf607xLeprVk41t4DNBA/WMzCMCh7z68l
GsdvV0Wgt59NmTxCwMHYtiWObFELtdpcoVQ0zulKZ63J7Bg59Q7C+trrA2wgu6Yd
BrdGTWog2+pX86804UZbO+cEMh8d46rsXKruJAYVH6p6Ga6KXV0B5UJNRq2BGhFT
9Vs5jqtHZwl0+s3oU3kOGXzlfbB10+9NaC+4r1I2inW0rwRRY+G7XqgxdJb7nxTU
n2OZd4eRV8GimXsJ2KFS3gJ4FLjIyh5Kh28s8niK3EVca+p55/+5hFjnAPeUK1LG
bw9FpC8DQCkQhTQAd74JTj55EMFC8nnbHAYUjlJ/S1UAV0Vy2hGe2AcEC9DLKUjh
SOdWo7P8C5lZZ1C+OFdIedGiY8nVAFEAm17cSXwK0cXIosdmMOm2ajPMcerGRTPH
khmHT/43mb68qbUSztMoX+be8/7uKECG6AV7PwLX5NRzmX06P6wamMTASR9VHv2u
peD31s2MbPTKqH58DJwzixHcn8OlwnIcGorgrFlIaUpA5Gah5kgvNOPAc/Px6uuu
qOB383KepF462dF10ObxLvJk3+IVTGyMyrPiytGd9DAqvwlDB3uechM9SyzRE5Wr
elmPm8hURIOg96DpCPibyFzQeOXOXKvn54+U6chVHZDEqdMG2dnAnie65SFJVkCy
6vBJkO/K5OQtbOGUOgiLzn3jvEZjDPMGACtnt1UDfU5cXYbQ9ykuowaxKttqCkQC
6bg81aGkB9ld5pwieXyhX1P3Qi0zixKhV6txu3Gf9sobdzJgkRRy9cpHAzDTPwBE
xbusIO8ffW8cOPnIxQN6Kp/CepEMvSWEJsBwuu3FOEdFqlUzO/6OWB4PTkennkVn
YvKGdflOIsOPEpDJacIQwDlT0riWuPsaZ68RLB2DMzGq1V8+/REuynkrn0k8FCT6
ohCxPRVx3VeYEZvDrfB1dhhdzZEZjOrBt63fJgSiT2lEbmQMEvzDzA6yXHnBBFOo
LZunkMxExc+5leO08z8d1CsNCZ+u8mJhacp0LTgHFX3gxfg2F75sf+wkHa7RntbS
8RuLcf6GPGp7USS3YBkaP7RShX/M9DJBL4bCU4pbTW+yHKOIPLys6WJZ/Id58tUB
uKTQHHVDTDkSjQoxBdlODL+8TymCHOPmPwNI8fexBn+Rr8hckPb5AI/LKazN1odj
SX7pPAx14OQtVmGVxN6hjymsJbBMaMFzw8bWMRLBpzH6JR5ePq9nNinVgBmFxUwr
JJ3xfa45eKDjofA+EwN2NNO2Y2toI+TkLYSgItGuWp1tGhqubjSvcp1BEp/5JEZt
5Y8ps80/d1S9J32DdWSem0/zZKM49CV5GzYcwONLbuSAYjwZakd/95SOLGCGrQRP
yzLg/w45Kb36W/3Ff1LLUOt1AFPMzDFAxNE29/k184SRrsqTPeTgpU/dT2MwUbkb
8Xf4pjbvWfF0RKgNITiTsyV44IpaVzyvUU2UR77BD09G/S56/H9F3h2sz1Ys2Rrs
IuKAdezma4HD/Ne4JpSJWOuYYOtSUUCbtYPP+gOP3OXQ5sFQwyqJ80MY88vYkgPm
SxC5yFXTu83iDWZxvk5Z4k/8u1e4XVv8xlUErtcR7YOPmW70PwN49QvhbQ+X8891
Qb6CAD8CeTUltnEVZDTjKR32bXxlllx1BwBzekQEWoT1LJC6PqJT9nuXBrlykrCR
LR1nM0PVDOamJ7jfCfkj1rYbf07LLKRJkLyU4eLRUOSEeEIVQbhrmUr+TkYCobTR
hYFhcMMHS+4zsT8CO1IaimTTW0BS9M3RPs/tv84oxuP1yFwRssrrn3LFKLqwz7Wn
WWw5HO5HAeMelyuPYIvZYr292OapNwMZ2eN8M8RGx4GPXFx+bCGA5X0SFjEbqE0o
h9MLEJz8dQ/gchtdmqvomsahy4KS+lvJThGdwJwadI9jr28fxL+nSGXH7kROzvTF
3D5dhax3GxfTPrVFyTRYevsLjCPKvTNds4I4IWuGM4GBrbRFV4zQdGDI7ABwcZEO
86HGz9oFgoX7b8PobYxukaqnPJSd9cmOtRu7UWBsWqt3NmHB6fZlxmU1os9T7AMr
Q+H6RyTcLn4Lqyr180/jE6aYuLmfJZOyfOybGiK/pm9uhm3PTT5mdKSiLvj8tkgM
lSanIg141CJf9Q5yc6bvKYXec8Z7tZeLR8znJ67OKAdVuiS7Hf/UO19P1tiIbuBH
47MQfo/yiVaCXdoaigD6c5llOaEHJJpr2xQsU4asiOlaJM/19/ccITEbpacZoccZ
kd+nETLz9gCX87CyXbgDIRlOKPkUtHUR9KYMg4PXikSjh//FaUcdU8Tv/E6GFF8Z
UCaqtnXzTCLHacgh+FUxYrBpui7U8UwMnRLR4xFdCSV2/4aGwKRA8l3pk/WKGmqA
8RBI5l2Co0WlHW/Rw3b0KTk0qLGy0OkQSZjdjlCI9RjDHtdj3vUajcv5EiNcwDcl
j4lbwAgAFKxSgmlPjErLv8k+9XA9aed6YXQ3EovxWIYxalBWdA57EnUmIc3RPQBb
1IeyR9m+anZo6aVh4194bMc2J8MkPWNKNy4J0HJ+wl0ySKmQT/LNS90SOCTiZvda
/zPemcEBK85va2yWZY+Ll+s5gRTGah3XsxHNjlEuJSAkwE/18I98cV8AqmyryPjy
Cb66k/xevEv9BpEk+YjW7O0fw8x6/VcLu7NjyBGDBhppDlwzgCpx2eJof/rfOdVL
CYRG7gqJPfg1BKWfsr6d8NC/VF7b2cPSglIGdKEGzQvH424wJ0TkEDg1MZPykTPD
QDsNgXymPegldTN87+c2BsNsFf4W78BFxZJISG1eGTGYURsJQZy4Ib/CGtFlgD6S
UsR07z3JGsuZYWrblrNmC9+Nt0LFMWkei1vzMbGmbZC6r3WN8o6RMSfwmwZEp2dT
aJzfGFFBCDuyOW+XBtChWwJRqIWejhOfgNVboIqq/RTpRofxRcDS5Hv0LUx0+wp/
PHpPJ0mmMgUerqG8bIVCo6FzfmxQSZZqrT5biYMGcxbk0Iho3r1UtOFs9fAHOixA
T0VYXsm+UpRvOl5RSvqpUY5IG/rdVT555+6lRgTEIezxF7vARfGhoTQDVbdYEzIz
uJM9Le1xVPHje290x6UGbZgLkpQMMRLF71z33oSQQ1ZJnvpelFQhSsXhl0fICXEX
tGahZ/1ozuB8fWmttOOHeN3B3Zl/sHPZYC4Iq6V++bNnLEss5KF1Z9Crpitsj5Py
B3k1iVPh5x23k/dQ9nZm5VtbasUQlnti98DGKld5XDScruOgBw2+SvRaz8rfRzSY
kOo2LwWFYiSIr9zLEGXUynbG3iyboAkIH7GihdMIB+HfUkx+nCuXj6rNCp6kvSfV
EITwJaOEs1ZzZvZWEtlxzMmNrdAbeMWFDGWVzQyVp+ILBM+RqcdYlT0hgTnVxU0g
W8Lj2SZWSJ1PApjbZ9ZeE78IC8eeXN3h18zr0hS7406RMKmx+yTff0G2dc+4rdYp
egopttkcxFP+GxJDPSQPBaQDWbuTZj7yWbXWEYHfALmOX+h6R7aSHOl9XrLYF2tV
twTG+bnwaxvTruhvNT6ySaQ5lBIZpSjmBQ5lmRMJVXKG64s5oVqyfDN3sbVYO+Gd
Krn4McDuqJ2zhzs6dmvRIBfAmSGQ/Oc2nGmGLDUG5A+lv6jPMTfjgRu4DgkqYI5C
J0c8DN0Iq9LY1eigCymehkytNcTDq60Lp1J6R95zSP3omWSx1mk3rNLVRng4hxxS
jnJB1et7OgMsjZrlUMcYthYyotVkzAV/hoBjiOy+AYijLpPDnzByrVE/435RzfYq
zemYwYl7UQ0GolToVJ2X6SR/n5BPY7WZJX70qW0O9Gceatmt92+BsEl1lGTbNFR3
Cupj3zcTYcgj13J6pn6kWxOTJUoFBsmS4f5tJpQ01gY2hgq0ICB9yCYeRRQYaAho
N3Q5Y2akV2P9F0zvfNJ0RP5Q/5q8NRzER+ovGlCIZI21Qh7xzZcDJ1QZi/+INGPa
lhkwCFog+NzEbB5bUePRGrHirjfdWLSucSD5BtsfAeD0clQp7fe9e6voAL/13udx
J82jsAWEL/HQI+aexglvKaF1s5pBcZBgiXscYOKPlzW7bDIH954a8pSixnTjq2/z
wnJaP5bQndsHPQTNSUvAdqOH5nveN1UOsElX+PG6Ll8rEU2K9WxPa/EbsCXpBz9N
Rc4gr/86TLRSRoKTlM/ZuyJGipDd7K1mS77oQTNVh+U5Q8TgN8+JSGPTULQp5CQt
Ynw59AZSvLdSOlOp4sXKtz7TTMVwXA/5lGUFdGmfAu1p5b9K/T9uaxnGihBnEMKY
/YQS3UOwwIM7mw91uJUssvlEQkxsjx1THxunVm3Nk2ikGnFgcbWVGCtlLQcn00Uv
6nQ4s/5FK/gNNXma8Z2CyIOddmp7LpQfpeef2AGWr3dUSp3MW7nLJTQC4ZDl67UA
HttUDn/vrrDWd+3K5WgJgr5+60aZCUO4s66i5zaR0lxYEqNEEutMrZPlw4nGkqoA
svmC5G9f/PcqrF1GEOC6OHnu/S0hUtSGQw2gtk20CXoOK7AVI9lpyHxP0Kz9EHfC
Dw53VlqT2rGDFuNVXelZN7NZwwMizuLMq8D9hyUnM5PniGTSiAXImgp87x88vqb8
PgngPeUYGNEif7jTUOT93gOQcE4S8boYdsb1sBTNS/Wk3GsiFFESm/pRaVtbv+19
DvXWwrck77+rlIa3EXTWkrdcGqdTr56jOyMt3OVKYkqpCYsj/1wFbzG/fZ3DRhxn
yzbrXIQ4xpOQcB4uYoQ+ioSI9GkgshCQBwe2XUUA0HfjxjR7yQvlN+lxdUVMXav8
CekYVpMzyGBLRxXiQoUAdcu1jW/SUNtm1KZ6643aUKl1zrbS1P/tHLu3cpa9fcoT
C6iMGUBsf2BZF+VO8xVGgtztvWypVzbDMYcmu8WiijJIOt0E7TYSz1ran/yThGBc
TD6b9oM6zOSlELsGz6/VeM/cnPy9bgIh0eGneimXk0ncX721R6Ey7dMHaBgR9Vlh
5Nn/4ffbM+nFJj0c08JweN+kl0IF5mORKz1EHDSUO3L3dSE1W4Hr589Cmwto9H59
OFZwiW2z7cQ3fjN9FAFDHyAxhUEZIAb3IFDQkPrJlEo6HdurWp89Z5ZrwRimkQSD
jRGLyWZ85ONxfb/ms+jtQb92SPIspPe4sBbU9EBW5wdYY+BkZZYnkjDeQRWItSJ3
rAgHDOpZSAC8wruQfCtmRyjef8fiVpRkvWU3ysoIrH7rCFfTF8ISgnX5Pb1D9XqW
aZBlHxGg6otKWsy+39ftxs0fDch5SdNEZcrzVM4+1w2gqzIWvC//t+8mX+Slruht
O/lhfX/Cf4S9lk+Th1mMAW42SqE0Oi44lT1z9x7JEZMaWbDHwrrnUFDhZ3HTD1lY
4W/uOBN8u4k9BWAXNcfD62YrniPCBzQ38Af+dolE1mWXQxbHlVcQhJagQBHNkMAK
LFvCpjrwR/fis9YHYLQRHvUycseKpD0r09UsZQJbMbpKTYo43ftxQ1Nl8Gx+Dszy
OWYAuNW5O5OGPwYxZE++mV0RvMaRTmOfJagAOqrlVNOUPl/6iiH2NYwecMOOiZsz
1/KIe04AEMFUhQRkNzsZD1w/nPBDNtSueW77lswmkQEgsIX56TUTr/K7DkbuvlX1
VF9FGT7BuEYAET9n6xEjFHiac1qnHUIv2uQZr9HqmPQB8H1Hd4E65s9A+7XJUsCs
PJXwc1ayskmEh6UEYokYxUNrzUCHxXMaq/kZohtBwMTYGlBNgXr40TGHoh96tfkN
V/OOD7KruydLes020mdAVuCGJCHqwCDqBPXnXCRNWa2VOfm2AHwNBcT64lty8vrD
G21QpAHB/S9g2AVF++lxgB6c7K3S7XM5+j+45cibALRbtt0SCiMeAQ9I07gsbg9W
uP/64MKOtnDvzcLW62W//CsiJsOaYw9Tdd6DQHHE1yRPcgSFqRHeK+KPrTmNOMXG
ckUIpPRr22Ctv/9jXbqpA41ixVT0CMhJWOioiIpD83OU5S8ilZuaAtBRwP6Ef2je
avkjJTF07ZgF/Iq6DtjvWNV6/2UY5CQb8NiRWmV0woXQ9gnOlQl7thqfKVDr1WKD
9V/80CRzDNoVT8Jps3QrHf26YevHqQd4SpHSctv2LCGrYLx1EFsyZy89nc7jPusx
UvRTXRYswpCGWCY/72wMXzkq3blXvBR0QOoLKGcmdwdV3gfqnThJO3J/pldxzIWt
qMrjpdz5+CqU+JBWMzf5aj7ndlYoJkcLG4m6L/NtedpDt7n/c2iE+D9SmNN6zZqe
xzifT+tmonKwtJ331qQBcdoIt1K3mn4XFXjCohIMz7ItjwTlO5Uh149+Q2JYJ0I2
oAZao5gMahuziD6dZy3DWj2Tze4cTjK6T0k03vqxMaPTslkd/Nf18K1dPgwcnC2R
Bo7ToiZZ4FEfIvrmxCIL/J40T0LAVRNKWWThEpMzNmdU84FsgYqCdux3sNrmOHo7
j7P0ADMvlJtNclMBJ6pS9yPlVo1r5LMLZZIs/DQCa14OETEXxgOxOnY0uRmnTl1H
FYtANHeATC0S+YgvM96BQdsUkrd6JfoWzXlgqVSyaXR2CTpEqM0f8Rbz2waG3LXg
uFUQyf4iGMQTI5tA4X+QdN78ZQQ48057ffIF3WJEwwNPdyqOyoYLIrY9HMRJHMkN
zG25gcvAZP09DlrK41KaxG06Jt1INm8HPRkNZ8iwN31tVSngBDpNGJDRswck+TSY
WIA512misLh0tOYdPB/SCedBo/3744EXGgXxSIkK33tgDTo5WgKuS/H5ESZqKc7o
HyghurkHSuUHWTVy+ecBBg/wxZiXxPBLM7nfPp2eROHFBIB/B47J8VfwYQeaQ3T/
SsZvHxkvP44dC3Wmx7EvbCSi7boHrrvpjOzQtZpt/3CJVFxvmmbMZNculhGQglcN
WGvLCmA7Vq/K3d9U/o/4TCNfqoZX1E72bQ+UxAZA54eiybxBKkl8HKPoBRxw4uFM
qwrFOstOzd60QaVu1Fg2J5TOk+YLNTcLc0oNSAPJpA+NCW0HO754qSQgQduzNhdk
Wmd6a3KW2ZYvSEbwDbkvMXkk/DDcK6V/9wx8tIf/egLtwrrzCoeJ9rjTt7QgNEkt
BbxBOst6eialaMwNi0PeENdqqBHg3W4BQcMir2iiTVYMU+fT50CFyp68zgCxBofl
movk78m8HcrDuZVbBvHpsVNr6j2iJCthnU4NY5615sc2KjgKQlqm7ymiFH/rILlO
7KVBJnxBjVR7uzzeikp36z6VMXRwIYcQE8SMD7/34AOn1sTQ4OZtmFe5ENoJ7e+s
STaX4m01+sKNn2K5KkX3sQxnoQo4F9Ii/3aE1F9o4YulB1hUarRAOQVkKrOEgnwu
8hRfJzN7yW2YPWgJwMDTV5nv0X4zFLz0ed7cIJDBs7ArkH3KZWYg8wGXZOfFHWGO
ww1iC7D9RiPOc13Sz1yvhoMMERk5UTL0qIaHmwTNAE4MfW1/eJ8K93HHJl3onFeA
qqRerb+oohoKTGQ109cmsT5fQSiR9P4h11jWhrRQmh4Woq1zADpJr72XQzkYV4AP
HErmbgfUjs2IKFg09tYFmWekaMUGDvLyJfNm1Cq0L21E5rDcIqVCaCKULXwbR7rC
o0I+tE0qcC3tUPML3O8PFassLnLZZvl5vJzf5giuYrao3Y4/ZYIfFQ+VvKOdlawt
9Zo+hL3RvvtkYlIZxg+pfbBBUVhMvUvHTJEK6NPXIMjprGw5GXiyXIaeaFrIeGQK
6s8opA6OWZkRPW8yIVNoOtOiLqnyG0ypIn+gcf0cgxBv0cYnc+Q5J5932DKDOfYN
RGBSfLoaoKA4jo+F6EgA8gTXwR0pnMLL4pEHPu5R9FvzVjFtZxWTOxL7/WUJit/v
qLFVC4waOeJX5Tmzf+MZKTWFegI1i02ANqZapDWwqva644P8+gKO2pACSWNG7jeK
P7BgnRuUOHw+eGWdyBUY7tMAhVXUj2SrWkMtFYr+GyF1sVJRYGuHudbeT/e5W1vy
n3l/VZbLzCfDlqP7NUqS9rN+/hcjXdlD4cmEspBeGbjZR75EkFD5a03Fh/l3c5zD
OkuB4CnaosGnjnCkEWv4TthRy0TdvT60L7Hf+d6gGYQRruvAuKqPSKnvpi7Kmh9j
p0z3g87yTh4FefTUqZVA68SGyyluUeQzAQjWFfR7ze93B6Uv7I7TQkacRGTHMHYk
PTgQxKFGp49fnKgWFoBNYzIpQRVD7EzGl7Ne8cC6vnbcJeEU4NbH944kaZ1vAVMh
bagXvGkTBgGHCuV9ZV/TzSXfGvcu8IwjjhyLaUEU0r/tyHS1VjQNRKQ9ud+Wwviq
Vii8ZuTG5yH04Dd2TbQTEb8ma3ALOvxL/KNYWtaJwv16L0Uxbu/YI97Hq1fKdlCa
G+A3YVwpjfb0skDzFM/r7WFCoTvUorkNdzlQwYnL0xxZkn7hY/GJOJ+AU4EOqCBP
rPA8oi2+KVjS4pOzW5KKjTKP2qvCiSsvkMjA3Dvs3LRo0ZXvA9X/Z8vy8OAJoYow
K+h135Y+seuIJaGir+EGHxaCrnXTWhE/0l6Qtqc8nhsIB3d+STBCG4iQ9AhuVYHF
8W96TcP7IgorAAPIykO/SMtVD+PuuB8H8Qv5pwU4l2Lq2GwMvUiYypMugX32R+lQ
EyJ06rYffcOSF/hQMIj0QkeMbkCl3qpsUf8InptJ7L1K1T5di7ts9gzvoD3n07Fi
LCqk4LTjePRlbBktM5GQMARI64fpSpP2B9TXWhOG6XmqSmW10GaAkbUpcGNpR0MJ
JR1HaDq8aVdj3jNo0TOVRj6ZISmJ3siXHB9+Xs1MlO1F2VIJbSTgJkq12USz0huY
v+j1Eh4Bz33BTAu+FOTPT96NZfwmqOqg1Xv3tIPs/n2zSlMFtxlGcPup0/gi22xI
UnUoc8oLhFr3fCQHzYWo3WuaTFkp4v4Ebui31QBoSnYHupifC1nyVliXb5ll9t4R
PEW5InMCCifEhrcm5sW0/dlh++ZcrYgtmSW9CL3OcSSHRJsmUl+6Fr3iYcCsHIw8
VG1lwvWvJrK5kOO1MR8I/0vw7DxSIjXwSIh6Mquolf9IXuMzPmXP8rZVkAa1OdcB
1Uny8ilhcKEm8udlu6jdj9e7KU24nED6Nnt3J6Lj9zA8EK1nMdGVyi0qF3qvETDN
YeEISqVZyOokUE6eRojQRV5F268xBxZprm0dS1d791qhEMuRqRgt7lf8SJTTDqs2
kJZQjXIXxTphomL8E9zbpuhOQ9uvF++x0hR0IvkQnrzRALvE+XyPrAObKHP/tbpA
j6hD0DUlL+gknLmnjsspoP98wPecQCf/iMbD6hhaSaXiBZUBYgOcC9ZAADehWQzD
33Ny2mZaNiARV7nB2rAs+p32ozdpJyXlBRykYlK+B4PV1kXL8vjARPEMIhxj6eFk
klMiRKwd07RpIJpZmpkbT8KvWZ+RJeOuRkWgKMwTEx10e2Wg/26o6l8aTqaI1aaY
XhEzC/cZ/mFS1M6JmVRkNmaO16/55bxiRBBh2+gASz9IMwuvPmR1gdIbpN71OlPd
PyMM/pYiYY8wtpWyCGpn8lNKDjaeMJm+P4NxwQdaqJ4a997vj3c/vYrgZa8mDGb9
Zfz4zZvx9qLqgix49V9dBAgZ+wUgRKTnvC0bqWZHVegghjDGm802hwniHFYw3vGT
TPk6Biez+6Xsqc98x3RomfMD05BMeM9wwamzUzAlTzAxFYNIByd4qVj5kWYqOhMQ
QbI2KHUrB2kL4bZ3MZ+RUOZ7W/JqTOjnEG4fY+Ft/MZFp8yyU3cUHwp15vFIDaTu
C9jbIbTZvASaFl73ranQCloJRY5bMy2vR0GrgCQW7JnvVuuIFENJEQnB4Hj7Qqz7
maD1oXUA4fadblio2uqXeaUJgrKSdPDAQcq6OIfqdfQc67cJNIdl4M8AH3MzV4zs
sUs+ZiUv2pe9HvMh0gt1ak7g5BVb0q2ArdlTDHZsZ9cdmsCPEsJdVqHFzAAtwVvY
HoE/p10hxkBAeocOhHwbhcBqR3BuSJ+MO3TbQv3iwbkzLCJx2U0FtDdDqrTOAGOh
gerNKDYZhpfg4r8ApkRqiAkM4wYUOkIThQt2ueljVx3FPc71/F6u7TL2wk1evo+d
wb3DMct/khz45OWNxbxIwQmHmxpapfPzAf+q2Sfr1eyzk/an2scFut9ZXNcfS8zZ
fHpq0EgONPJ6JeCN1Y+VeeMgZa5MJR17C4w3Eu5qm1obkDxhqOcavszdXjm/7tHS
o7f3G1IrQX61Ga/ms7wKISY8OMuYUE993JF5+75jwEpmABFE5cbYTDABewBHBBLN
ypzt8EJq0fjBAcHFDwTvwJAW+xaUK3ikJAN7sqoKtggrI50MgHAyMQG/OgKiOeHJ
7nDUFrKvAuU3VfjVvtSEw8Ye2NZPIBt9ky+F9koWJBwTSJAEO4wOsbgm4vgp7bO0
E6tHISst84hEbPXFgqQkingCKRvYE0LxGQzszldcysH3/k5ZmeQC357JpsOWBfvX
pyJX9dfchdCd9sAH1p/FfiDVC9rkysdducfWnRt2BdaI/cMPu1lipnHnAyywJtEE
TN9aPNWn+lJ+NLRyD1gkHJU5soPyoXJONI1aul1wcnDuQm+5ZTl0RAjx5YTyJz+X
uidq5DGeU66zsnB5leizXoRw8yu5yK8LuJh9eonTaRoIlZMFCPSsP5REBCUeqjZ7
4GlAWZnoB7V/fSFd82BVWjgrOUk+Rb032ZZL6r7/WrYe4d6HmuQPO0YYsWlZ8Qgh
xRgn3N0GAyS5hzYOthHSijb/eeKPqJDG9d33MdO/oBrQg60ta+fSBCBV3mRAmAZ+
F9byYn/lphCkkZKr6huPB1DXCIhZMaOQY0z4F6h61lRZGwXfxBBg0QkQqM2VPxvw
wZ3mCc/TrHL/JmB6Gk96+g0QZ3zYBCyafFUubMNOKkKKg/gHEhduBp06lOMAZmnS
xpgwzcZBaEHI0PsRTct/tDyyV2jfcU2rrn8oqd+Qh8a61hJzJBtvEuRnyfYhs5aU
ep6Q4/NCHrEIQN1ACjb7LTVT+1pkrlbig0Xh3gu8h6odb92AOEFWAXtUq8pW6iRz
/IvucW0232chg7UEK0sGF5qv/LYb9jSS70Y0UrEvkFqTdNgtQBxx4V9EkIozXRxl
EXH+SQugU1T6r0q3XL2m78HeTOcGqcHeGNCIyVH9FkAYPgXv+gF+o77OIgdS/dXK
zWtU7+EUX1HWkoAEYDBa9e1Or49ucwsgEQ58RQL/zmouvyK6GKSXhJTnRIIRpxEa
VR/RCRb9nbO8BxX8WGZXdzwhZ46OCBgP2DAKXsMid2fu6iVqKsuGyBQfagueVxT8
h6fHhjT82C04pEQ7YaVhGWnTHEowfts17A9Vw3IujkDyD78IHT6Gnaj3NFwk71Q1
EBOvFKuZ6uy6uZXFNjQNSYfry+KhTsQjyTu9hSZ23/RjdkMGF6HpMxr7nyZEXmgI
LidgkGlxjWq0QfB7yBq83rGzuGGtXM4fnVx41EDSJA7j+OgbGGJ+yR5RBRdOStQn
faLGJU8FQ451miXnpORtJJO0dt3ST+XO4kMugh3Yib7HuWLa+cUogpwjHX//JxD8
7LHt9KAyBicE/2e7D43TA6KMgENO92aauyQO90Xh7DndxLfI0XulXenp+QKiBNzV
yg7qg2rwLv8Eb5YhXz/w4yRk/W8bkNbZLK6u8dZOHm3JZnSTiDmx0YgooSf/fRuh
ADd+7jowNhWOU8XA3u/acowgMVzUHMVDUGmTElxKZYrQcPuOBiD2ghm3oSkP4vXb
2hnybhG2TG4xg9IUtGGcQK5+HLsfBHXN0WvP4roWzz3e4jxFEEdUf3xLpFdJsvTm
GyeN+F0PuBChyXJBoOfZsk3D46bk9+GOKPHyQjS+rGrGJeMUtetJE0kJQzhB9dzj
OtHc3qVAcCGJNAQGhi/syhhKrJ1fMylwLVXgp5zAOiecS/FB59EWo61KIujTtitV
f/FNt339U5TSL+QbsrkfD/AXDtYYPC377UDvKPW4YTRNqpMwDpQhdfbhuuWtDaEr
E+tZ/hHOja85bk0tnsXokJod6MSwanAlGFTbBPMwG/xRctZFwwRNJJ+B9MOcHARZ
swN4KY76q7RtcLqfnMR4SSguxXqqffQwMAX4j5HAO4MpBoBBxWse1gmdeYouzgeZ
U1eHyR8o6rjJoCE9OUjiqylP9a4pXoXtW1+p3AToDsuR6tbPCiUFpMTdvT9CDy+R
vDBU6YKB+zbvkgBehrq28/ttciZdTT+hT2XItUMp1cgiBCyIjeP6/xMzAwrcFAiW
yX+dqcwSpHGOm7JSL2x6bJoFtbnAqc1HZao0XUhy/ML2EDMtaLd4su/GtKW5se5P
3XXn/mM/nflN+zEi1VMfpgl2ZntcA/W/IWNLiCbJ9qS1cKHDUCqBJVGme66UlUPS
F7lGL1MP+3ufNXLz6j1AO33dK+xtTZ4ToRYehVTpksYoLPZtLSFONqEz3y1VPK3t
tqHArrLdwm4mFw7VBYw/AX+pKwnqIJsroLyc917P2i/gMC7O/iKOd06RtQ57/JUy
FKWwKZ4CyWAk+qSdrXZGZeqPJXXoMWnsRJyLojP0LTB2r9ZPTQvJrcJEujIVa8Wx
IWHw4snpPfq6PwV63cpRBDj9AcGy//AhZTwUfhWMcveVfsW1QeSDqesKR06EmR2t
HzlUpbgl7EOnrzhsSNVFYnuNDR22WayfwOUL/cU1p95q0QvlHEVvxQM902us8xSy
brg/IEzSZpiq9i/tR0HEpdKtyVAR4UiRBJC8Jt1nrsSPFYNX/KlGSwll1EhsatnA
nq0oFMTEwCeNE3KxGsR0lHourNWn5FcLLUlxnWY9EDrZWicWBV9qoB5/GXxS2VOM
0e+PYI1q4WlMudMjMxymgvra8vgJjJx4QHPzHED6i1kRXewrnGycl1jW49MKj7iO
3dF4H77SrcfoMFPNBL1dw/se0IEvlh9QhIgCDT9aATM+t2KJH0DeB/WcpuKX9dJd
kCvC14k3DLz4gOROuySYbsvBdJM+WNKoi5ZKO1nPQK+XZd/qpDTEkv+U/E04zP4X
N01T7Zn21L8YzOROoCxFFRiaNSL0J/mDm1mP5F1nJiRLDKDeldElpI6ypXAQJHMv
nK3DfIS0CyJNNaNdTJN/QxzxUnxdW03yOOsjXLbnjKik63A0bgj+1Q2RkAXMbmgD
mJt5wRaKt1Q8QJPDu87U+BwDSlY1Ov8A9lZi53anscauBzA6MB5kOj6+bthplv9M
/8dshLcqVodoUNs0uXC5ng1GRkFc08UeoR37EkfzZYwaxMS+dfm6DP4/eG+OnE7K
Pw6f5AyqJ+6IpcUkr5sSJoMHEuVX0YD5xj5mdxO4Q/W6Putu2frGd5u8PxZDcLSZ
kQ7tQtK0UsACZBEnbpQuKQFAYl24exqTep31U16pmeMPh4ldjaMLRgP91p+CPEnT
9g7C8m7GOURWfTgGwaBvuFGJ7Np/AMALzS8LZ7ELOl2lYhPOAbpquNVbQikyMLBQ
1izN+Nl79X+TzGkEqXChVg3TUxydZtxQQu6Ws6tcQsFEtGkXnN58InU57uEw/PhA
FRcr70IW9So35y9XB0hRbVVwc4UKNWRVCAsiQRN48YXVxSu95qir4TXtMUI5BAeX
yf4DCutlBIRq4ULBJQ1EVkUF/kyFpJWJHUsJXcq9bmwroJ8l9n6wqTSRryiPoZpG
Zq3YhS+WWxfw2wgie7Ykc+AgTcvsnhneLyHLWkMa9YAkNSfMioj/H01VVGwXpFdb
2YPB2i9zXWe86N+FFIE8jchSEPc2iLAIOsZfoDbQXC9wJR/SPEOZwPPVrJ3xE3FH
tu+6aeZ72L7F51ZRiG3rvBlD+2LFNIAbvbzwLn1Sv9bqHyzL0znBlak+s/Ut487t
rEQkxxou5XpsIcjdbkxWJmDCDp+GXT860EW52PJus/RDN5Kho60sjH7+38uYmYCR
QruwY82Rd51Fs247RVn9rf9iczDIjJaaeP3PfAKybEEk91zHRP+mAXL4GieZj5/z
6AzZqZd1q9tNyGFebeaNS29n7x2O/hPJyfz/6vTCI/oft4exdRUwryV9N6h7mAfp
rXCy/ijaEt26bukMNUe4RE41pADkYy3YEm3DXrMpe8k/vdSYl5r7u5X9yBNrxTWZ
Dl4z06SfjYxZqNUHxTKEOBRGOPzN6MGu9oU3JVdZiTSHbnWLDQEuGabwJzBRK/gm
ejEwgKY2BCNNfykRWZ7FeKUEo8McXHwPxBdY+e5CJNaclnlOd8PK2TDju6JhHRIO
LbWjsJijVpNjy0lwE8UthjrfWAtrWrCb+5Seqo+jBywIQdyk6UYoVEd8L688UzhJ
a3OFhBsZ5IfoWjnSia3cnox7YHu+P77iuzXFB6L/ARJVCzlf+FTShHiPN3TmzT7P
i7nGMrLmIY7pLjPHXFY+tD+C8+wIR88MGq9PvjQHQjD/ZvYod5zNyeVLxjX+mfBx
O7ZbNa81H/YK+VhMVD95Oj30ruWT+01Flzk7a6Jt9GxGREQ0WLPwo31Zc9V/id9R
MEymmcvkOxeZHIR7snONUMBdyLfQOS7gavE7gu6CyxIcSbCcmVtHTNSTpd/XWPds
stTfRAJ87JUIhGMr5YEQIeQUy0dxkF033+mrvbodKQXfXPgKVbYnFi8xGgIGm6QI
SEVueDQCVsYNS62FbfBweOJf/hAgQFFfwUcjCAjXOMmNJajYJSIRy1/jne+tXDs2
NxfnIHc9l+QGZYQlnPBIMZo/uNlJyp3A2LFa5IeCw/Yx9ty0bmFvRy6RD5SbXD14
Vegc5J8GZNEeLp9LSgHQ7EwIEGY+vl3pWzwkmRSSpcK4LLjRgs3YA9yHaiBHVfx3
RnfcdufDbEDvHMPzAczRr3VQSoTE6qtGKL0C4FRNKHk47/lKmvPKivbdiime94Vl
1yv4bOkTRJuh2U6aG15OZ0FLuOgo025nFKMTMRll8BwgOThiSOD6Z8XHH7QpA/Bk
vtQmggQ8Ji4k462Iy7hRAeYZDGnJgiujNhH9Y7vEtv9f2APOtQPtqQg3Efwg/Elj
wTX9B/66NHIlWRf+MPiFe77tfAkf7MrkSZCToY/41do9Gaq9isF58ZjMdfjHyyPX
nt+FZhHo5jI2JrNcMVzPifyJiVLQwB4SNuceJ8qnojcaWXkrqhNYCqsBp9J8wqrr
PkkwrFGvuVLDMKd5sgYGvEGGi8i9jG3XQtyuXvnaOlfsDO/8IF/AfdKXEgLOsevL
767ut8OHiL1EYfFmmA1fe7la34jhRUuIV/C5lAGps0vQRh7PpocKcZL+aMaa1Zsm
9u8tUpSRMdMnIcjaVXvtAE9YA2I3odNnkEKC7iPjM8TBhwwL7YqRjIcRdA5kELX2
z4lFMOLUEEVpf4mncLa6xffWqia0g0ZpqiBErjnXrI2RNHQ27Uey269T0MLAUbGn
+VyTN0EYyV6pWyLTNMk94GF8Q4AETwSwDWuAuU6tPE6La7QuCwfiVcuoWGmtnbPN
J5tPmVyRYGtnoBRcB5j0AIGgZ6e2oB8KcQImKm74V3HtzG0VaH9Hux7pG9eqlZO8
3EXMAe9lWr6I/D5Nj89Sk38xqBNgDS3uksgc4R+Ui3MY+07JzLUz8vVCGLhjuGxA
1pLSTwiELeUCIMHacrIxsbT6Dzi5UHlfypYP8++D5V3xhBSqcTF5WtC2DJBeTwk0
a14/1GVwuf67si5NSFC+KdDMBNPMBV1bNpdlKHegDMGn+VTI+0apZcbIHH0ETnba
UE3qCBVxkuFJ4DtxgBhnOsY5IN48atTowXE4CDeiM0OnWs4JWzPUiyEQYHDGJFRR
iRTlycs9Am6ArJfSrrjlpqG9IP8vmSliRXtrmtpXvqPs7YcDuexGpHGF5aYBL5TS
dfdFOBrJ3V0Gw5Ib4TcsnU3CLm1CgJT8gJBoYjDN+hGpKxf/+RrwaHY+Nb+Vmd+v
HZCYQTEBnGqJu3gs6ruhP3Ekz69IZTe1c/RFcjNWLKtcTxQ19lHO4c282nEsWEGk
mIteiMwxa69HitaFN1XEcCDSwKTHLBa7lvTPNOSBglPgdMxE3OA9LMjcBBsvOWbh
0ftGL1YIuq5ImfaXo2F7RI0C1s7RzgjU3a3LFyC4CmJRpg52tNMrpffXwGugSXjF
HImDsVD68rYl0VhvHv9jiPCgvhYsx9QLF9ehaX6A77Om4PlVT+6YMltmb6hYZg+6
3+Tc4OZ248s+7IkIa5vyJEfsgaM685sxrDu9q8hvE3JqVzv0k8mWVCWp7jCSPyWt
wtJV6kTahoIziz7wBs3zz/5B4wIuqpXYLn8qc8jCjyWFjb/0/4vruTeW1pdaSwR9
Q+17IJg7Ngu11lbDQIaz7YX2dAehv1U9XLd6Q8Ywo7WDjH09c6nw9vVsNU91mESZ
WJr1RmznFVehGZONhvD1BHtLnoAFGa/Mnv2Yi49Tv9HpyObG5GDVUeJYl1ffKz1v
tPZVlmecqlSsPX/FrCGlzd/6YbWkiwMeZ1tZo7rLOWUg04vJvHpqYbTl4HQaA8fc
CFyJw2oNB/adjKdHylQhK2CVT+8hE8j24OvhDYfMcuyGUaZb/UNPXIPzTpio1jt0
2et6U0StpjY+d/XPSKuoWJVmb/p+93cZOl+lVqLD1owsIP+YEGXvDSF87l81n4m6
umHJ+xScAtse7BasroKSqKd3GMsWnnbX+EE+8u6kkb/iCOZQNYSCCLfNxxOXujpz
qrTpe1KQSeGN/o9z2Oh7DCGArAQ2H/NW5KRXByE6r/5Y1Zwzy+2zGIXXtwv8Ixql
GsQupoLZanpxXlnIBGZQGI9S/kDIe9n2/wD26xZ/jax2o+bnbnJi4rJF2woS6QHq
+4UK/tEEvEjrOKrfX6YfIbJNNuIztmbVIxqlcCKW0us3IVMMB9Wxe25dwSUxUi0/
ysF3o0y9QL5WxyZ/mYAfR63GLRmMG2j7o1PlWOZiGX44lXfRlN3qG8XZEsj8d8dN
28FV4SuAkhs/6Ie+wY0glcFs0np7BpLmZNzCBx2broAEFPAwsPVJoCZnLKxRnGKz
ZhAkAlFJT9udP+JylNH+4G2dCboyy7lAbVeNAeRE/s6jr1KD5j64cVrHCi8su2Jg
xOcaKaCMErnSqm034V2XNOwQwVuqv7p+C76HSX9Elxqh41Ed7lQpMNNRztVEvVIP
vKfmQL0Ybo7fK/64QhGCnrFIrM7YKuRO5rd6SzZzWlW2Pli+SUPWwwtAXUwjrG0p
PPMhkeOnmQ5kvctJoKmf6c8ktAwqn2/vrFE/ftFOWShGeT+svu4tbUgObmf3JJ16
Z82riBWt+tERWPhzVsqzI3ziuJIJoUxzvl5fvjtwAQM5QGhDkcbx8cDHul8DW1ok
3LhvZCaz4/c2gj31RsprP9pv49e559KlPY32aWVw0XNw80vGaHnypxcXCkIPDPwm
VMifKMzwyD5atBgGWXHyc/5t8FMSUss7kdvd3DtDh6/O84Q6yJ5cwJbKEe24NlW0
Kf8tNEfmBpfkEVD6ua03I52ldQXIgvR2z8DyvfqYjlhS2oj0P9GfW8QMduDZIwhX
EAG+sjw2mLuBB/K3JGCavThxLr4FePpHPHMnL4v9u1vq5SstkKbpQYLRmf2QWZH5
tHScAC9uPpFk/vPGArbCe8jSwxFEFySJXUjlhsdG+U4PKAeA8bX8QLG6EKXaMqrH
tc3FUuupJSwyQqom7c1HbnCYgRXXitYw5nQXIgFlbz+T7IcJwrz4QDjpx7nZUmiO
vRGuE+rYi5AjteJnl5RWWQqUfrlywJRjGBE2XAmlv/LsN4wubB+EngSSwWZlPN9l
w+pcLG2AfK0PkmjJ2UUgnyv3GBNjy9Rr0EO59DfFTTHHnDqBzDGZEICDWY8C5/Dp
CmOKTTYBYfXGw3W9KsJLeZBCHdDTbwzA5eFbHy6ukp6wBXEnVOLl1apjgfPVawgM
D/8dlwILMVk+nHn+c8dXEL2fQwZvDxfnDv7PfZoA1behsKPhcuvLX0ioIc3Pn7GI
dsLZ4uRi9t+JfVBP/1l1inVWguuJ0HojEm9kvtFb2J3Gc4Jpl530ZUjFGsccHcrE
wpW89t9HVVxmBiwR+qz6/2/bfBJNNha/u52CGPf0bzkzPmX8Wc3oAXQPPqXSyBZb
vuOlfxfDsa0uXGFSKBGH6lv/Ur88H8GaYTAffwj/zvR3EjZc+EPw1tle0SvcSC7J
jc6Felj13LkeNuekmiiH5ZM1dDN18R5jvkQWHTh5jtWDXf6+OZe4Rm9OB5WveIXK
9YSgl3UDkMjdOpM173NzrCQ5eErsuwR1cwZlE8ZyIdIeMR7BIptAWg9nkmLmRL9z
euV7GObWC6l5T0kcw9zosRhRW3MYOLq1akjJI+BN7aD7FRLxs0uryR7iVGb69D9w
pZa3trapibXYgEngezyHYtEHIrZm34pwS7y7izdipZi6oL3U2NBKEHv4sUR4LPb3
QWyPSszA/U2uWVns+QGGS08vlrFxNri7jDxyycWpuoVbF6GYctrxduo7VL5RSItT
07hLVDt2WQvIOSK73sEyYhLsP4D2UyedZPpbcq6M2ULoYODMpuOF8+18v3xDvyaE
Df4DseqLxyctw1WalvQfJGA5k2pAJ29G7JhlWx7jj+t9mB4njRgVX03HoE03xF2z
Rw9hh7aSdY6ZrmKFsyf0FAYqkVwcdSEplZVsmTUgo8/tVczZj8ORAr/K5sLOS3EB
6vx3m3sOvqJzGMGuoX+Df3vW4JcB450Xk1zaGjyIPSb1Ham7GIUqAFkA0APhWkZm
gnuaRCOwU458bj//6Z1gaoT0bhEhX2BKLxCPT58R6TNsiFHlwpn2EZp/3H2ei1hh
rpx6TCQ0L4M84a9k069hpmtU1u8xF5USAjWejYGsQeZkaiSdpD3/hYgkEF/zOUHh
YNDyaSU4MPXlxAG09rx5E0r+xA7djQB91+C5G/b7kvCYjWZY82fxwHC3GM3UX1ZL
8n/rYjy6CDl/XkCEqml3tPUxoKXFmEXvmXjW1NTrCQl2cabW+O98Ybnr9wRYlfhn
yJp3eGRM7RX400CtegUa2D16k70V/P8prvFxhErLPv8vvDS+vvBN9G6KApFpeAHn
HdwbXIH+hYTJn0H4USBiqX4yVbODexvhHXn6zUcjsVka7pa9rPrFV6InayTjksJz
ZP6fH5ttyJecHmnFmbhJ7GA1h3b0UPewnIpjpGSspeHpnbg5gu+NR9Ub+rPBtAL2
b3KbDCqz07DAdZ2+kVV1I/6XfEaoB2KT5RJTKCJRwOcMrn7tMTFoVsoF2/Yc/Rla
mxjNQeXh64qJhyYoeA3wJz8+9AcCnkOdyn/pV45J3tRKx6AxvB3RpW5YKVU8ElUM
l1EMkql0wsoRGjZCEjT2YfF+ZwqXaFvMZjN5jkfV03KFIBkwkTm/zYe/GqvLoNXN
4xN7cPpXeUnSiZqn91xbqrx4Rin/Fesa302iM0qzEWwkCGemYACXaBnOkxX4K7kF
Cp5oE+oywfNH//6waayqoE5jIfbuQqFh589XSW65eRXIr7cm9cOz8MqhQXZaXiyi
Ix/QpxqyxfmJxNmxrkcXMfJ/6E8b+6Oa2ZT5UuuByWsgEJDVqsiYeWTsE/t6Ebm5
WgHwFEkBBIRLlGbkup46J74Cxtr68Ih5zJsbFXcplp51NxQosWuFu+DhP/CtgrPW
rCoZLjYolw2fhz7X9SUt5/tY2lxBfHUCG35rCrf63FqjIIjN4PZLK4dViOOVm0oD
5S5IbOm1QA5rqB+8fwVcq0jNQSONiWhze8Yk33/GnYuFE/L1sy6tDvt39xZrsXNa
KxkzaO1u4ozVvfb8j2lgAAReJnHEf21LYCd4lSbY+BJj4dXxMFy5sAakTncTGNWU
sNhAzRtvvdh9ItXkAqoOQNy7FAba/fW8RPLUL6EUrsENfGAeRi0yjcyQyHaW8Wbf
eMkOuKWSY2qik1A0DiNuNe5CqHCes07gBB4kLafnnisvJSc5dLshFGRHegUNyCXK
GTCsFaUIksbp2mynAnNhSzHA73/FUqa1phs+3fmuM1eBwdwFBwDypqIW7dXU8ywH
vl8pJC7j6AA9hlRPpArSAbQYFcKIJm93JqOqnUSqKWjQ2Mqt6HJX7ksoJemks+8l
G8dixYuYmgJ8PzUdYcfNtI+GilMT6U05ymhFV44A5Fu1147n8mC482gIeA1QuYWi
ph/HneVDhCQcSSCvlcT8pB0H5U3/ILWIRslqwFRWPbiphLfOSw+6Tna723fDh9VU
EYGC3zWZwJ/3fze5kQPZuEyNgKkrFkDyci1njwidySanqu79a02JgFek/fT9L8G7
tGywphdpQ/h9vNQbLUbNv11IU6oVbVTn/Z45bW7Rm5+WSmhtxHjG6Hyv/T3dxwmm
VB/FVDQQ2zrh0UA8rG3zY35IQcKr8+myxQKNq5dyVhuK9s+H305+0xZXwG6HKjCR
2yG8gBtTMZp6Tq2v5mh4DhXVo5SCJYW2lOwNfYebTOgvC6TZJnrZhDtqdt5BCh4K
yV8O1E1Qk3VDmRB8Li4gV+/kjHAX1G0Jk839l+mbbOFwFbF3rW+Qeg0ZM2BbJQ9C
8VCxTarr8MpZ4SKIrtBpNczsnjD4hZM1/8b3j0IME5h511wPYHedEw1Ky7UUWwcr
WsqPi2lIG0+329BwGzG8vNdOHyE5xMM3r/81gCA1BcuE129Lw6IpuFyqsHxy+8SJ
6u/JrJ3Kp8shNDeuARuSaKb53mgZJX2K+tkTaJhqX2c3oV+T7ZYQAOSPlbHmr5XJ
Jfcj2NyAFTc7z7lhkfpiQY70uAbLq6iudC5gXDxyifDAOUHTBiMC57bhJC9OLYz5
fd81mORd7HE5xiePsQGN8RpiGZbNZcUrzIQP7TOKelybUq7F80t6lypvk8wmxBLU
oGLptP+ezb/aBZz+FAo6fZJ0j9UwamZRy5x2BgWNKVAqOUKa0vIXkfc1SOIryHQP
EReE8QGqIexaNCNkr8ohxDTYNNIPrU1EpQm6D91nrG+cwDDcEWOwFxn6bVCk2JPb
SWAaZw4DVy1TctGO4vmsyMb6E/OxnbjbNW0jDCAu1l9Tx5yYTjvPnKGqeqpJS4uz
pckWQlzMw7uaVmCOdbdrj0izSLfDMPmTT5VH4aFDUGi8IecM6OV3uFF61+HGHKTq
VJc/Z6y+OVZ8tDkyqfTGQ3X+ru8W1USUF/8OYPpBLh26gvTXsYlCUXMGSP0aLmOv
hhZ4lvkftMk2yHASJhSt3/vlDHaUkaZ9lmjoF2HjeaSbana+nrNBEmpt5OrxryRu
yVMj5DIzeBFR4S5pQHaKhksaf3hsK8SGKVxSqhg6evaYpn/lsSFCvcK9BTqytkJH
B4QFqNsEv21MecV8mvCamd/wteUs2oTDuxCD34lJfMEVD9HliaN3CO7Y1c4pei0C
/6dbQCo8UDyqrydZ445CvaeE2SIIsFfrYRGZ3TY5BW1Tp6KzBULgTKvmy5eUl9U7
ieHmVvWWe/AY37EcXWBQs9xmd3H+nTk+gDM+HvqpT3izzERua6c//JVXKYUx9LLO
HSWiJKcy8nzUlG8x3+H61f5XQKh87qIucDs08vLIJlWaND5ZLNcu0LWfc3hFcXGH
YtA3vEJt7u2Yp3rryuKO4vKwinhNxovPmzxLhEczwtQDJBoZ5SdHltOY6Xr5lCtk
qCH105JFlipQkSWpTFbYkc4SBxGNOMD406ycoC0gWH6EIx9LtHum6gCJ4TbJY4wZ
iNu+ZjnsrjJ3EEQQMyLrRu9SMnh3nszHT7uLYKFRuOaK12zEzklUgfSPnkUnHc8i
3bOmgWz3AVCtlYkJHluL2ADswglcsEelJjPuKiDwTTyFaMrdYT8mw/fJxZazRsWg
07ba3n897jzFMbFgtDfhq6nN2oaFnat24+QWqLXVVk75bGU47w6jFpnaLg6k8Fts
zcgUtaJ5akZy43mnU1wwlGnShjCMH4vwgVs0bdVW82iVr1vVumvQe2482FRbbRaC
9678rFOscNy6/HI3PMIR5LY2lLHyaqL5zhmC9AknJy5yOM9YT33Rl5yAcGkXlDkL
HKBrBFCVgZ5w5RlrEvPHQ2IY09D2jNKOQrFFhQBm8GZAIKi229EHef0Yt1SEygsP
2KK1yQuwLqScAp+4Q/XdvOocstMxJNYoqOilhJCb1ZRo02n5/5Hm2t3iUPual6QS
Su3cTd/os7JVUNuZNCfLrkkRlJ8uRCZtherfC0lH9gHyDWbtUvFK/ti7RtYzUQwp
a/dtVOLUO8niUuirhsapsbMAT/Ikt9fbLmILAvMpOmdKSDgNmLyp70JtiUyqMaNT
imb4UM80cs4Psz/Oeiaf63Pq09WSgYb1ZMXZ/nXh4XWr+C8TLi4b0xswHh/c/laM
f8Jif8tfStup6OfHsrpxM0tFwG/6CTNlSjx0J5KYZb2bY8/bhyHAu/IVUY0AFKpw
yEUoCVL4zprkOg2h3NBlwKzaZ6BYS3LqDEhlxL6TA1vZR8GMPB1AO1Knt8iU+exx
F2yRkgXTL0TeMVfNVxbMuQTWE3yCUwPu4kE4zhIOPZo551cYhudCi/TrP1uTMdLv
bHIxWaH2LX4oymrpvgdAfHtX6x1SYASy8iZaRLZcU+Sdc1hSovF9+J52+ZAUP81L
cIt1/ThMTjudZHLOQhPV3ZqamJLXYjerMl8N2ZUoh7+W/btgGF/Zex+NEQJ/3bne
1Fl40R80XUgnhJuQl0tq9QDvh2BvGepXOQGw4Wb0+YzAGVceqzeTKrym5ADvpEhI
7Bm5eZyupLln+MWAdkZSyotb2ttZxzUE3rgRmJGYhkGZMfIY6ORZlrC8iP/sajEz
e/7kU0s/H3yLYY+Oufj1hflZzbPqa7v4RoTnKl3hUeNw/Xjy+XjY5dSmWY03IBMX
S8CNWkznjA/tkzhnPbF18KE50OEu9KZ0oc73igsCzDCdPCr7AQCce6hzYqE498Vl
5to5/fcKSc+Fr0rHR9TCcMVydA9xyfj6v9Xsc1cruF8DkSjDtLkFmOv2RvwjLSEb
EQIdgxtzmBQ44QT65h4MFdR64vbo/cOc00vmii/1Iqslsv0/evt+HKkaxZXIDLuv
LadS0qgG4ETpQJS2CHLgkrgCm8SjBiH0z0FYDWXy9dkp83N76aLgAab+dism2mOH
ViBIkTUm6E21CPo/B8rtBU+sG/MArPWYmXpMDUmGFChtVdkUbn700AtJ6JdInHir
ZS72uI7ojQnX6iZPNju+4a3mQO10tz98En2iO6iQviovaEgezIz5mSZFss1aqKPU
bfXF20szmF06CHPQS4vziqiYISlYvhoHDx9lEd5oD9XyhyHtS4UcrFulQJN67TxR
bUO13UrP0pD7OUh49K5GK3UAEDJXjGv03EJWZ3w5SY1qHgy07y3pJOgOe+SZ49Gg
Y/oGyhDlMRymZR+AuQu2fvZYFQiFn7WMzcfuOyP/ialm9L26UQQTF4fP/ig4IcO3
fKPaANg/3by43VIVQqxWsLM46qXR7AoXALHGZ5MjycvvReMWj5QXh2FY/zxiAKFs
reC3fORBQn1uVhVOhCA0l8fsoMrOyJye/IPHD62DyUy73NaSF+6bDm+9hnbLWDh3
k4K4Vyh8eVWgmMMKOeFr6VwpsBUEJ8vtHc/PfyH+lr0FJvicdV0WdUp7Ch72XJw+
QXKGTLlF93YBBAz/mhYZxHxrt4SthCqBwVm4yrm1vJRLFabIlXN8wjsUqwIAZKOf
3wIhjW1xAlvjP+1ptYNPC2yxWdesfCIhTAgQFinn6JacaAVy8B3U0I5aMfBVvH/Q
3jsGc4Q5GeyNqisbh78RddkMuhaUWdpemYKnRqT5wAMLn8DDbCmqwNVnLDmClmEY
cAMaEz85trgwokHee1189M998AKf2ZOrUrkCV/3LjnGCHEDDcrDogZEck6Cx1D2Y
c4HtH4DGPZWGVSzQXzdDqaz4gsaxy8tF/WTC02XjYpYcgftOSBr5coGndgRporlJ
JEgkH+TqiXM7WbRpy9fXtrKs0UflNA8Kde1kcQAae7/rnc6RSMM8g2omMDSlgw6n
uQYJOADIT6psox3y/AQTzcQjSqIFEGMKtIuurcSGg8AsaVKAXL24LyinV9HY9imO
6OGjqvFlFpVGyh8zBsPGQNJUSkgJ+ICsm6CzidMSi5AVmkedg8KqezYr8ZvOTz5z
gY+i/ADG6LLWfCy00EK0ZyGIpFIHqjQnQX781sO5CFjFPKjrtyeVlZqsmhwPt5uq
nHQSXG6mYEHGWzXnf5H9LUfWHSAu3Pbt25HCk6KIGKsme5zEEv76BH36N4WFu6r2
46ejMNmlbYiwKcJpc7q6AGq7pEf9qTTD1R3aVHeWLkeH2PDDtEVqwDbh+iJSrS48
WeQhfpQ1tQ/R+qeXwiEnK0uvTo5nK6dW4TCh+GnOWSYS8MEHcVvpMcPRBYuzzRtj
9fd7GtGZlmKqxddiWY46zxO3/uYgVj9hXsT3NKigd9x0EFChhD+yyOXPsf7ir49u
II9aMAU9eHxlYMg3J08cxjRRmqvpqbFWB0k2smUEh2u/HKtkLOJ2dOKx89l7p92p
tDCC59kDbL0+crEzBtJ+GqDH7Cj9+BNB22Af30rt5VGMnHsct9xZXNNyUb2rIxRN
7MB+fT3aLA3/IQ8GoeYvAFuE/nXk2HMWy3Kbve+Py3PBXDBxjkOP3PM7kYI3iHNL
uGXBKmqHJjHl4BYejk5dydYnydmj5LaatXpvgodOeLQOwbAa2Ht2pNIkB9fYPc7l
TDCc5ON+TFuiEmJX4sFv43UcTYuADjmSlaOJ1Bi1JEix1bTAPwG+ujwBjyX/NPTW
x3N7qSWTlTNOvwPXLvUH0j77TLdaClE9yuHNXAEpqbxJ0uH9aWZ4mHOWDuKsTb2c
L6jSrfhOL0qV4KBD8l09YBIxpF9g6o6xACxKotvHgHPqI+UMXcgOxLUFhglw201S
nYI8hOJ5wUL4+jyyeNc7J5J2IrfKtl8qfe/QmbcMBEV+huc+LnuNeUD7nMIghiet
AUl70g7ddqlssPlamVFCiIR86+myiC6pr6ChoLBjraXscNsYLzTNO9+3AuHTNYUW
ceVZwI1z6CYbl6CpibFSJI8QmiU3A1BxV9iw6+io9nu0baa79F1LXnj6ZyCECA21
ZvavhMV3qJ09gL/jbZtdOZYh5gQRD7V0OFhL779e6fOZzUVh0LYNkEmDytMwPKdm
gIusjtLpBzrDONceN2HaCaH4eElaYy4oFpp5R2GUwWDlU8PJKkvFlEbsYyApsD0Y
wcyBsO0rSTvFsWbiLESLuXuJtkUiVaN96ifLwS967Ct1sx/ZfqEEYBuU1LRFkOVV
beVJ0WsO38reNi2UrQmVqd7k96Zoi0wkYvBAE8anH3rbXEBvIMmlTVqpGqo9V62J
6EICro2BkqLbpHT/TihaA5VyZoqohE4osQXpx1wL7aoxeiLGU47eESS25AyZSiV+
TNOQb/QPCitL5MyvbmjkovgzkEbwjeQ6a+2ZaQcV05MzZgHoZuPsU73gmAP8c+fk
3ZsCR2pbAFbLPdMidtHztqQY/UAyex4yHRUwdMbvAykLnqG0JW2qiMkjvpaqvW7O
Majxsa/dOPw6HsRXpai7Woqzc5RD4NdnUflAN+zdhGBOcarQGXeD844j8nwMSEu4
YM1Lq0Wf3P6FGnr40A6ygjEl6NcQ8rTiuTZF5n/1sAiLdd0uG9XnfkDWbY7bNtVn
VYokil3AIU2hYZ5A6JrDyxfKjeEWpGFk18we1w5Ml6Ic6gzYfwcCUt+aLMtC3MvP
GuMzMiDo90j4mrmotIQF/4edY0n+ArwemaqnWkGnziWfvVmbnMKQHna/kttimhxb
s/3N+8EG/c2I5mggkHQeQpYrvPKJJPZljIRlhzXTxXe/Zq/DgPawuwHZlVBn9N1w
u8Kq8TOl4+G3y9zFP3ZiYRWEghaacg9seAA+AsA6SHHwZATYQwfy7HtO7/XGOpgy
YwbmwUjAQTy0xRnMMeSzb75YawoiI66gs5XktYBMFZac+ARs+XdqTx7aDzNJ5ibu
jtqjec1YZcu245/yYt5BpcRqH7bcNRnjYpgBhLBIftcgLOhjRnwVXtoipUZ2h9Pz
V1ThggkRSI1FIWbZKkdCP/pXU1ZqEfxz/uIUsL7nmvhGVGcOGEmflUOOylbEaiia
hvnK9Izmotsev+N7EX2Yh4KjfBzeH+aahcV9hW85az7meB9218nT3DKpeOg8e4fG
o/8bxvD4cE6vb5qSEsVXjjCrRgKYoSFHZYp5zxxcj68Er8VYWJhI0N4SCM1Oa4Xi
nHqxfuVBIgplVj57clRTHZMu4ZvNRBWofarpf57m5xfYPoeK4qIRWMIxttlfvxFr
YY0hULS6ugd2b4YKUQAoipHnJ6rCy9vckr97r7XPYScmnODYRenozZNq2Lxh/K3J
CBYFThcPtlXZ/QpI5KaXOMJ2nHZgEMWj9I5Ocr7iIvZhY/fXOO4wGsH7UHFs5ZZ8
r1TgzIClcyoCN6Fukz4tn9VQCKxuU41m72X83+mYu/A1X48Wfk5xzzXPoiM/TiOE
O0X/CzvEaclGBlKNe6cSQR4+hpX8ig2hRV7xkgZAfQztfS82eQs4GkGNwQQ+cxNI
VUH04LcpGDfN6Vvh9QcEUWRWUfmNQS4joYRojZSR/UtPoEIxNYe+Q0yhQCYEkz9m
CqPuIxkSWZrNnOwQPqpdQZHVCwnHevM3wvX11oWo0jpLhJaeiidBO0T2stWeDEIO
3gVs8uK4ZCYLoTnvbcCnhseWP+65fjhzF3G77rjXXHSBd/ODKXKHSB5Kgho5rAoe
WLWHJV1U8cXEXbt+OssqSQMXkOl0NYRRTJ1xOikbf3WpsCUxTtveAdigExjmP0Sb
ST93Y/f1wdoKKBakfvET45IhniIMhBFL4NyVJazCH7pxaEcZR8EPKKWCOB/Sp3u3
iD+aMrVVy/NjhjUVVoE9OR68MovsAFn9wPnmVgSqyM1b1p/n6Pg0nBZ8R97qQNcI
KfEhToaU/1mB54tkO9R+o+apskQP3qfN/mK8vlZb+ZynB/IFcVGZhdr/MKs4SKu6
fm+Sij/6ta2u7TpYf8EF6XoVmX1twfo9xnjmIEaJw5e5d12uW4tb6h72CNnBdvl2
paMR/1qHa4uMrnTs4vn8HhAFdyhacuCSc8onL/qzbOUi2WC1+2rM+mWz0IkkIBXO
OsFxXwMY7mGnBj6XSOMkbGYkFKxkWlS1+QhjHVkPYo1yA98VBDfHFSyu1mEUewiD
6H0KHJ4ipN4ZTxwJdql1evRp4NoK/Jny9U7/hUvvb00jTKWOQL4uYryX/A6cYibj
WV0jFl3PoU/7NLx6B/+ywPmnTqAG1yyY2tCPQhQFXf2F9/AhJ85Y93vlqSkdB8Oe
4d5t9SHNB778q7uI5qXmXKO+wl8Xtijafi1NruptBgRV7/IPRuzalLY4dKJXRWzi
r3FbO3MrPF2PRgm39Wx3h5RO6Qaazkl46RYsJulijQ1i0adcQPhNsS+Ioxtn8FWU
r+E1FiGdZgh23+gzlbYYcMruVuzES7pC/9FbODLuSkSH79lQchtY+363I/sRyH2q
NLCIeVesBS7YTIppFhQ91s39r/EY+hmeXlAbLBQbfaQTNDFRNgziSqFK6i+rNuHP
c1PNndPBjf4GuX0lQowau857K09yPhs50F5y/F5RhxUwj1EqgRCK1dCB59gCYYua
ghFobE7lHcP5KLT+BYgGZ9+Xt2nQEl6mBikmj0uFjvnfWwWTb0biNG8I6k5i+5u7
6A6XN59+aR1jajVe+G3MIoeoILqOBqRYTSWGfOA+05iyqIAKHXdgfnnJo0AprNFb
iM6cfsz2dK+rV8u70EcYMMun0cC3ZgZXh5us9H81rane+asuDtYOexuQFmR7yeUS
q5Zu/TL9Hs1m6soPAcVqEkJSNKc7yY1472L5h+KL1XHF3ehrgEbKHu4GKNky4HfX
NrS67eTM0mxNESLBdEHadBXSL+WWNBg5z2T9rYaWVi/AdAeZy2tk+SsN1soguKUS
4wUXnig45A85kNb6W4Os+XBVicSvFz4S8l3JzHbt7pG2+y1XVcwjJvWBztyGFyzI
xE4EkA8HQM08AYBSmf1CEC0Qv/cxMm7sHZph4oBtwImcW8/3kPXSEyKSCXcnFYJ6
LH7DKd6DqQKwTZXWQRNPCipVHnAyj17a/YARdSjqUKVO8QhGSM9+oX0xKNroPKvi
7I0Fb4OD8FJ1m0iBC/uwPTBAfUFPjiS1ylqufDi6L1cLqMRsX2Z/4v557392yxmC
HdKeNUPYS9usz/nm1qikL2MK0kZZ2thD7iI0Jz1bHZr0U0IQ+03qUUcK9lLQOABl
uOhoJ2BNi9QvDSIjHbA6wh46ZuGzFQzbU0UYAwbbRCf7NNuJOMpntKyGhvyhXViT
dvTYDYLsxeY49lRZl3XikcqB+C8BtWDchf2b0ohKlYs4f1bn92r24GgahKg7APJc
b/gMVhOW2H5WZu3HYs9H3dIjXs84U/o2xs7MCWQrsCfRtS8ex8D5BijcO6fKNjAV
7WSbS0xFQQl0DXVxX+3NAWolQj3gXN58qGWp3h3LXlue0fPTFAMnr9xVCIHrvDwE
1D5vy9vmf8M7iH5zB1SZYkjpIlfQqYegxQWyO5le4fYgZ8DNFaBB5rmY6DHdzNp3
RmDlmSkwHEeP5yByGY3l/jLpIwAKucLceDfW4KIOCPzFdveht1OslWVP5Kna2RJc
3y09M50qAg7TgcC/ww3s7BkuLHASXBn1ucFJAvBoYEoB4XcOmO/cogTPjsN7Nudl
/c2r5U6G6/E5WWEWRBcPyneWWp74zNv85IbDJ+MAwpChKui0zWRGhj9D0qPuYgL5
jN8nEe2b7ILThFrPJcIuf5REt7SLPwkZmu1KBo/b1AQjiKtMraLiKXJHpFuD5wpr
qyNh2meTfHp7O6Jj9cK41kUQZPaCWFsXKB2N3r14Y2aRGW0QL5sWUH2g7jNV/y+i
XOHroXwGvL7FauNIdNS2Zuk4rQtmNI8/paqPd5XVyGk9Qxht9GZBaaKmK6jRLfqs
Qfip62SeYGx+Aem2TkXbo7XEfhr0bFbirUpA8Ucxf+BST3YYLCv2QlkjTaQpdSRS
vCMgbmY64Po9ofLJJ0puCw8UyL64aIoZNwAzFeOrshAyotg82OCBYXPZwAO2E4xL
399shJAD5K71CoJF0Gf1hrMeZzhJ3WL3OUNRVc81daYTJNGgal71W+LSrkgw9qnx
UlIAXcrTR1lnN1NiOGIZ4DFgztKKiAGCThngFr4VYCNt+A6OtBsVA2Br44UIWbnO
dr7M2E9jYY3v7uAa4QjYLMOutGwcthSe2XaumlUZFQJGcoU805GUFs2dEtZ4Dg1v
nJYkKv6BVxA3U55ruIbJwx2MWyl4XBRjZMFRyjY51aQIa/9CiYSnVR09eDwH9kV3
EnzzJ0fVVLaTTzcF6dNlmtqRuU7/8mA0Z4PvcRVPbt/wRZdxtugW1qUtN0Yo3Tbt
0iL1tRHH922rUiZg0rXNUTCFLXoM9jBMvdlfpCDRZpIDbYyw6l+bpkFoH69dBdbN
loKrb0RxdVqrmiEkxszCN1AAAJthss+LWbE3sh9992k5FdZbhQtNGT1nclBv++WH
dVtDI2cA0mjyAd8CasDEkTma/VaoMAuY4OVSiEo2xeHZhoF25uBgsObioqHcCyOC
mfN4blpY/dRe54iPyeiDLWZdaGzi7T+p8T8kryO2wwfHpmMKoojYKKUscSs9AcLV
gqjpvx+O1QVJpUG9dRLuPgZEhTZI+les7Kr2xAOO751BnmmxFYp9QlzA9qYtnbcC
md/EFvREV65Onqyd0dOCqXxhoFUoOgY2Ux9ptmGMxYJYLini/h5QYNGm4mM6Dwii
lwrkRY7eCN+IGqQ/4RjgR0uuj2xnGtnI9bxh3w+0j10JqtZVbaGVd4R6fWBfrkvd
eQvNqT8fX8mL/WyBmJx/ljhZa9p1Xt7z85KfdA2yNofCFSU3lr8lBFrwa5Ke+Fr2
f6Bs0gxljXfvXa0Tc72dO/UNOuVlD5DQOFJ7un7HN6PTux/7brv590x5rSz4PNOu
lGqNtxrb8XYzXne074UkUChuOEFw4tf+0Q4GH46eVX3DDndWQwW1mYgE1nCwfsFi
EAUZvKN2VrUrn42CwQPLpx2SBbiLZcfAF+7t/jwH/QDlLIKdELuZp8qk3fbsN8pc
+pZV9VbpEwqMz8Llv8lXJxUApp8KOJb70qVPj/+xTMJOdcHYzVJSsyegfBu/sHiZ
1Ki3mMvcUfvNyjY1ZZN1cI1t7lqkw8SxGhRypKEF2OBPuXya2oUob/nviI/aq8Kf
E/R2chRKdUqQ4nmRjnWOBf1j4oEpkA8cSAuabCddg9lXGWsUISCz4KzoYjJy2nPB
R/6X0o3NE7b6M+vGmimxI37EMQUUJRNMe29mC4HLuM6bNF6WUy0v8V3E4ao5FQa6
sRtT+WdudDtrM3rrXC4yh7AA3Z+opRcBU0CWAkEnNwSHMj9reed+k7+EAjf6dQoB
4r1ml3Gkje1CE/UXwIhuI2BQVfJfAe6oFkv0yGm1cvRBRQMqX2Qj+D9NY/uaBBvV
07tLD5cCedE01euiIBxqQviS33Z1p3BUMxdbrxf2sCgK8oWvFzDoJZGUa59jxApK
1oE46Szp1dQVOLjvX1SUetb/qFpMOW/Y5+wuNP53T2s8cSCITiUzA6ovqBOvJwBM
BBtjUnCgbjedyzZYonGURCnnctN+94X9Eov2+muPGTuUTb/BBJ2Ar5e/xPBHSGEy
H61pbsXt5VOO4GWASkw/63d3ULi3+eK6zcVh/yo9cqnqbM62BdrLKDBZ2i99k7cf
PD4jq2gPWUhLjrj3lZW2cIdzT1SPcvaNAZTx3nHe+Qlv7tqp706FCB4vCpF6D1z4
UrtAUlAi3mgyu80pTx9M5HoKS3Q04Z1NzFatdIaUjx9PVbELQdOAjqQ8Ay/d4VRd
RJ3Bs/yJqrEg6eLpeRQTIeTRo49qoHn793xEXerAkMs81G8DQijLbqHzWBd50gCP
lwMP2P7QRA7kes6sIW4y7Nth4GgYdEDa/xlfpKZVj8cScHLmGitepCi+B81PUNPG
OCJpuYhqvLyT3t+7aM0kl9AszSJTVHDeJPCLgAWH0slkvqqFNZWi+Kl6gysGGZVe
WFUJxan8s6+6NfGsRVbE8q5z8+6iAOvM5YEJPoSAmM7vMrLQ0bmpeF2ov0Jke1kr
Dnp+BIDVPIymFlW3cFBXMHASdE61WG6bURJnrRSwNIiU/F8N4qrvCfraxej9wcBp
bTAaOzq2wPN4dJUwbOkYgS4LXURReYnIB/AC4d1jxdAvzsay3DfSD6oYOC5pxnVA
Kte1E2wPr+L6BWi3n3KaCA/ZGabpGyApMk1NEMzj/DqLXNY4n2d/VDSQWCILoOaI
twgp8GEjsBkoHbo4/zm30V7ier2REyrBVjBGIlz74yvD1bpnkNKLnYaWSLWFFa//
mjeCafGBfZjbUsNcGGXlddJWtPZE79D0vuH+awWLWvegZaN9qIQ5TIydozLCbPL1
tyQN86BxnTbf1ZKnwkp/gcrqPDxB4iUJeYrP9rkdVIGVOLehFGHmsJeWBL/PUFk6
ySraIs2VXmNaJKH6KQq1jxrka61e/kAoK7F84CMWP/CyzBPBTvmFF7UGjT0FVW+v
T1u54dXXrAJw4DytuYjtImXa/lcHFl9moPxN/TlmJEgaCPtiawJUYbnoRvHlTAIC
Djnd9zdTD1dpfhp10e9WhEgv8JiIvJ29t/Sd5GJCkDZYTxw7SyrzHMwZIuUciQ63
WKlH/Fh5MZZ4q60gefIN+TyZyhay269kkQeiG1uQNqlFgaZ0XsAOx9oXy+55yOpX
iXV1X7/0tHiRy7vxuMBtFn+81UNg7lCP0QPyS1BpgkwwwffeiiN20nfA0kRt5Col
DfhXxj2dOlDC3sq1lQM86e69Nb4sd9cNAyTbqZTJ+W2csqd9DNqGXQPs6Xivv1El
W+H91BBbeeUioXomIJlHdHfP9L1rtsQ7wAG2Nw4HGPc5NDQVx1sQlUv5hPIEvgCb
da1nhratwqtdBUQrLLd20gm+cEYiox7nSEdYlRUgT6j4RiQ8Hk7YNx0X15Nux9z3
fTydycYTZks+//Pc7cm8646dSlooLPUOR8qyMsDU2OmMUWBTLgJhHSR+VGG2yTqf
EB5sMvIn6LPXpsYAI/Ukg8GqpPCa0KSs0vx8juztFXhOMgM+m3apWEg+ciM9u0F7
BmthkU7xBMLFo7g4ETvb0TbKp7AS2iCHvFFQR+BfMi1O6n7IO/UoC34lcVwaXLu4
rYNZJyn5mPFaZknWJEGEbXQTk1AX3gw6HIv3rIBcEYTuNKEWcYWa4jAa1cMiJ7RZ
7tMfSM8jYiCYS6z5t2C7VuwPd+1Y3/xQJWu8H5Ns8ijYSPiIofumUjuALAsSgbZ0
3oall1KXd9+pReKxM79uxnihxY6tGKiPFHETYcYITmyPv4hqfVGDOljcDUfGFYBO
yzVUYFLRE7+yaUCaTxutW3qGxYYAOfq32STr/zlpCQuba48zq8OBqPm1p0KSpj+e
Z590LxVszaFUxANdver8OdrIDvsTLs6krVwJHFd2Kf152IfxTFaqukPybk+/n+qR
XgySEL9CaqMradWT0sopVzFpG4CIpZI4U3YjQaq5zeb2iMnc1zjJgrOabgWWjc4e
dEmW0Y8UFRffr2aHBXU9qnwzh599PUrGjwxNcp3atjSwFwxLfpzt/krC0lxRowfT
Ha56lBxnbzcFgkzOUULEJl+HgcesMwp6zW/efJXWetAnkG0sgsUx5OLHjKgjXPZh
Ml216qrLjFJueaKV5ziNhea0MYZly8iLcyEv+MEnotD9a1NKYcRmX7WxOTZzjBWJ
3F0LzpLM4Z3OhMNT0xTwOl4Wg5J1DrqP2ohBcaZ6c5aDEXcjRedZN2oojY6xSddb
FUMqoJz/hA/JbQl1IiDj13b2QHLgcrvQtmdsxa4r3j9b/hMFlSGh6lgOSt8TfenT
dxoJzD4qIl1v7LNDUDwfL25/D6OFhxwtQhVSTMbeJ27hIsNvJF7nEmuDWHjRbGEQ
B2MH50Q0L7z7O9azVv+/CkN2F9OAOxKy+o0Gn3ndXtd1lfT0oSExVpp8inW7fk1Q
rRbIxnr3cHEkG6Nt8lAw5WFb/J7Zl+AzdfoMwWQkKNzt3UAD2XrMHJ37n3R3nHlc
4aDrF0532bb/xlXnJ+W1aMGAwmba46nMyGhfNFgspP+GRSQZhhqYwSYOBu/p/q8w
V+IKaJ6G14qohq9pYpbrhGrIndugEloUs/0GZPjQvFxskSNbZ35zxZ1VHtWnoXDD
JF90uxI0rcMFmBHyq7Kfq/B09vHWmiFLsSiUYqzV5FU6h0Jahgvw8GaUSdj5hMHr
Fby5qRXOMzr9iTLUm0WA5JstnxpADY0D5ZpusuzmyprVA3v/5QjW3k0WJu1dfjo0
RkhtOmLIcNnXzxNzDMjwqvIWa6pQJGkIib4Vvcq2DQTaWSHpJpHwZknk4M7vN8h4
zQRHcasMZPiW//7FW/9Vu4xFvMHy4gnkIJqujZgTG8JooMLleXfJZjC85rUdksJp
LElw6+l6NvDSq+AxNDtVTQBg+k8lBMQCISpXSzkIzQ1eaKaTEWaB9DkW5aJEIPl0
f7UlaUdpUttFldTsDPQU1cJh2YuBVVWDVo93JUGJbiM8k87+yHWoBARjnHv8wr7z
1/14p55jKeTwkVMe0on9uCL/I1sGV+xTQz2PZ85YrlYWDvK06iRnSvINZ7Ozjn2+
slJNlxXE8FFYyg9LOCyxchA7dttrzbwzHc1IQaWj3JAMlqffjHo44B+blEX04t3k
C55LRDg5A0f2yMOUdu0M6p83Fp2cG35iTpjO+vTDAMx/mIIqVhSM8xXsdYFaGXHv
Ehgp56Fy+np5zngHDTkOjEmmmfw+6dhqQyuAEFKl0WZOpLlp/acYb4g+/CnSKGDK
/B3Y9NNYXIxdWX7X834w0v1FhxmXW9Hp8GpoCkCuUZmkp0TlKI02jnUEw+IW2Skn
niOQvMnxXEK0jrZOgfnKUlGFV20YvUjrzhloWQKsvuSaGaSbPPwn4w8HyTQyZ/zN
/g+4W7iraVJkYkPAH53mmPn9Cb+Iu7+FmYXAbKtIiBhlkniavwQyd5uddiZY/apq
xCy/F2wLj648MH9ckViM8BL5e9EuUO7Aceaz304PPVWzqZ9Z4AAriwXQUIY4HPtF
GB8l9ZWvGGnZlxJCsp+W98PxTRAod0/jm4TWHv/pNv3XrGqgrzWc92G6DrhyYQMV
5j3jm7uj1rmWl3kmvJrhkR8jH4lM+ubtTNtzCp2uSs/tM6IdDVSDIvBUf2rhPx1p
WTMEqv8oNKrIOY2ICYAvQekkvEWUsOY+MO6maULadY9x34tNaECKyaqzgF0dSUL+
GkEloNNlfcqFwtuaVmjGHq9neOXcp7wT8Ex94PDAnkML1XdlESNqec+SZrgGWU0n
i+SwO/R00X4eOBpQ/OA3By+pkYAr8UJ1QSLy3E8dztqOchZ438WwmeElj2SEalG7
qtm+hpUOIvaKMzIT8EtpfIWYUdIUS7JN5h2L78RqAY56qGm0Bvnbyi0XS8H0ptah
ChIjko89W3QTZza2ywE/AXbawtiPyHNGa3Yr94NJmME0dVKE5gQnlw3r8Wz2PxUu
VHUvHwKmKeo8ts1fd8jCfInLg5x+572AHZqWhZwhk7Vehc5KxHHpmw4xdQKmzf+m
Dq7K72cxMf6r15lndEfpapsVzjh+p3r6uPSVCuO41eFt9wDnbK154WwPxoAQbu+C
vPDw+jodY8nVST2eSNsBE30JDMZhfH5HWPSa/YEe39WoGndXit9sz7iIDquB1/2y
c5CObL7qCuba+KF3LWQcjsLxw2Q/zUZJmBhnWzpItB34jNTh/s3/PIUYoeEZCVrT
07UURifUZuaAw2gvQwvzOv3BgVmkbBw++lfAW9LmqzzB0qiK3jjqu0djeiUlh2KK
uIKJkr//JTJSAdz1+DXaIgJOSsLDXzS7utaVkhKh453LeAvOSakO/q6n2OkclB96
YL6IpfIfYlM+45MR0DqFhN6h1ophlJaeMjYjIfc9FW68VyIOC0BOiW7/XJdwju3V
etLw3wxCO37jYKF1DFgm30ZLKo0vt4dbrBq9JJA7OuoHF+Wbe93duViNZh1f8WbY
oHedqTJvXz7mAztL8jXhHetHgVSge3eHNcqxmPrPFJDrmjJ8RK0GI4CI0Uf0z7ox
32mmNIk3bJagn5RUgt4uNuSRhK860RBbQJZsgTNeSPQa7UlNvbpqkyVyO+0HOgNZ
iKCC4Zd6VNturIqyZgKIAd+oOsJATqXrCqAhXE4sSUjb/rLrUMjn/5pcMJb3qvDQ
FENJFReXpFrTP4mc42V83p7U5GZBqrpasW/M1vk4wN9H4BIdlRdVNPfXO6SF5bQK
1SoXCO2nCVp3r8DN0nnzmptnWt4D050W2kN3FWVPwtN8KStUODH7iFGJG45drhz7
9I9S6iRxNs9LoXqlJUonBn6RcrpE2+fmJVWiseSRxl/gDIxq7OpyrQ9Dwy24C5tX
B7cN250IIW0HvRQ4PwijWpdunIkCG5HjIWCL3JYrYQbUh4UhpuajKlZuq82rMWze
Sgrh6452cNZuGjoKfXCXKIdWPVdb0EfY3kVtRqArCQ6pN+YYv6mjhyxZ+LZhM8sE
iCrirAQ6Ygo4xWHx+uhMbDIkKSKiC4vvUc3/4elrDXB1Q0vE4VVy9y9AMe1Bx1zU
ZXRHL6d4OuDaospxRGrUn1u6lapcdH3cwGUSLMxwAB+ajNgJjXoBTDoDykP0RVoN
qzCSVHCqGViDwIeqs6UOV67ptlh87GFb3vrLg+7plHAeE63P7501yma68y1gCYlW
53zcWSbb116gYl3ucNqkMAIMshRFyh/A5MlzQIkwSckguPQ+pMr1qEuoOFMPH7Zz
bx5Cl3XjiR42gKyXCC/8U1+EEblIo606N2Qt6zw4G7HnxXym3JpX2dRu8GDE0zdU
QxyOoJ0At+DBmUVtfFzK34bzZyo/w/BZkSXtuCxRrwAScR0Segl57vhk+YBzq8sX
RurLpuo/3HbZ2g+5cITb3PvE7ADpFHIaORD6ZJzvX+i7qLj9cz63QMw3RxkWlmoN
CffQqmEV3aBSalw0EbZxhMsyVhJIVo4i1UF5chlLqYAQBldW75zwvH/zWc6IfIdB
koJwGIsAZGaNRzl7f+LMrOG+M/xmVQ9CXriwxD7DozNPrSeSLTvdrZ0IjMLZApy+
3i2Zn0ULLjiPAfVoYYTLgjKjaQ5kDXs6aRxsRagxPWbP8FtG0nt0aHDleRuEuR21
W8YN+b8owixDorXnPMEolfCNaC6FeuorNY2djgr4RZX1tQvtShOZ28zgGw0B4Jud
ULZS1fJxQxmMjBil0AScQbJuJ/+mrZ6ibRFL6o2iCG3oWBXqaHG1kvvlAF+zmpyp
945Kanf/Wj3ysOCIpgx0aSNA2cSvdlTqwRmH0zjrrrspT8vuLNcuLILOQiTg7hJj
3RUhLdrLZhvRvQHNB+PTPq3bgyKuLGZy9AtVtpDRTgjHjbmKFPyIvC4tzLYWnaTF
9yH1bUw2o/rdg7PjZwGKxJw8qj0YCbcafvl324eZjai3Rb+fL8YmXK0KdtICPAF5
lEmzjD5rloTjfZroK3TQs7NrPz+IpYOMjjoCm6n/BXh9AeS4u8A4tRtPwkVW62MR
sd3ZtAx9f/t9wBmMC1nDk69TXEiCoHH5KliQ0NdF5WvTD7P48SNN7zqykkr70WlI
pAbWLs+TOweEQtvw2bzim2bPtcKXDTHl5h+cmRFmvvCAdduB08zpinvDve644gD/
9CTxiDkbHRGNpghGSo7bcOCGfm/KG80A5KKy9RZj8g4IrX6OfJhWl4rGuEvY1Tk+
x8gtZ5rrU4GsWQWZr4wqu6QgWhoCggZbiyM3O9YXS8XmZEnLqLvDA+JTgOh0kp1S
wCLaJKbZeP0WwN52VTUJTVzFWiOUEJ6mM3cGSKmKQOXjp/Vlsm9YUEOSHpWPxKOG
/IfmZCK2NVIIKNSoUBX/0rw88VY2DH5m8RFIUoDYv1dmGzzk6Li0G54FGyoyxTv3
pYLIlufdQ8YYFmB351DbjZah4Kkkaf8C+ilBMZbGqEuq/uR2DnST6Unmq1KHrGrl
LrJU2MR5vghzEuTTyqcrjlPLrrpducNbSD5tiazAKTLn7GdiqAK0U4Bqv9yOnTT7
Ah9m6gs9oiP/A7TvIpar6X5Yzn0hQu+06gjwVKmm/Fj2PE2HVHCNJVFhNv3aV3CP
zbhbva95rTxAXl4xb2b4fAyICUP80bFeUI5uP8C3GpsiUBpMJuRgwU6zHV7bm8kS
bBvPAbEU9lXud65v2dbtELawp+krF/fF2NGNEyEUMOtKI4zqOY2YYEPiYUnsZWSm
56DZ5vOAoTjiyTOSy75/4OaNcIB0EbQ2LYefVd9NChFT8o0H+RlV8WNb9ymGNPA6
vEkwmWXLOcKsfC2OyPmBSDdAEBjWKHl47NnYLfA6+t4/z/yEQqBzTiApFZd0IfFy
DE25p9Uu2Ep9RdnWfCbkV0YK2rb+y5BjcMD2cuY2EkurJbyvP/WIV2vYNNE0yoP7
SbA7rJ0N1dqd1KUIHLC6XLOmLRvgc11Clz+HnEtbe+urBs0SxJtl10lrBpPS8Fdp
nyCfGXkYpGi1gWEpKaUmldJgT8W4eTffOLlTFAG2/xlpZ3khWOLkDX2i1ZgGQClR
2tvR+z2RTRM8b+O2cezuiQmFk5TwC4rKnucCGfEXnTEUCmC2lHs6CRw4RNeitPi0
72kQ+Ir4hPJQKivB3nX+ZPu8s0CCn219pj9laJTAU+f4C135aSvfjE/4a4mmd7xS
utGDyna/zNS9uAajx1iLFE6Dx7NN2rltjcgXynLUI1S/p9o9b5Eqhrn7uetffweY
TrAcsTZP+ao0uJkacr0cfe4+QnafO+R9+5V3atQQIvc4irEOjjEF7UmxJnwtltOh
F41eYntYBQ2qprxjA2sQps5vt7jhuepoujKa06xPJX7+SoVLYFfhCtbPCBvJCgg/
AhwoknZW4a2ODg+H+5w61v7j2BOQB0ib6Bybr7S/VZ/esyK+m+PUp0FGe5REiM7l
1wHto6omUE+PW7MmCHno2laZLktrt1zOfEE2UOlKWUrZRItoL4yH7zrEuwK/TWAC
+3lq4S+5Xt1JACPqKj2Sx5QS2h/ALJkKvyXANeyx17BhSnwFsNXST2tvyUCTJqWS
JzkHaw71B0O3raVV4M9ukoU3nv/SqDhbpxYtET9zWDtYUBoxU3vVlXDnlcgiBN3q
Q5bobeU/3S5bzgMl+2q7vftqQTr9GlXoVT2odfKK9cUZnPBKvefeYoUmN+1N7obl
TjiUK4X08kMt3q0vGPksV13rFvMdU6mCR1E/CnZ/SiG95gjRGHYS9Ow9mP3jCW/f
wL8bAbBZN/iWRC2JseNddXa7pgh1TrtYZ+JUVB2sYLoSBQ9GSGv3zGD5mZ4Y31wi
SOsjUX2FiM25vAudytx8Ez8PdKPuy0mwqCmex0gi8ZBHOdO40fsMkfGllHnxAYfi
0rpxvntPfEqhaOS9lPOu5teiDWc+aEWc04MTsz9wplqOfpXA0gqkqbN++94Prext
ZaNqSnRZAK+XV74TlajP3PYvA6w7ueCaGfHC4NSbrGnpy/+WHKBNoCYQEdq9+Nsb
lFygBKpnriO8g64g0JUASz5nuQoxOtKmpB3mhApg+FJI6xlexY2aBM5v25yKOehh
wMI0a5RV3D7VmJ+O6QhmuzwDIxX5NxSpTP4IXdvo845U4Ih/m62ltTPSu6qMjSL0
7D1DMH8v+F6XFv9QTep8BKcmmcAB3qdP8u5h+5FkpAbA9yBwvFKjfXCd+DVe05wh
N4oCYnt3kgXgLahO0XS+N27fzNVSvIQBWMo+aWTcxPGINuyGhyB+/m18pE/qtfmM
n2Ji/tcsojJq/HeWM5jCMcCxS4+ufiFqtQXjpw48RTv2OBAl9DAVEhRO9LDehg7F
N0Mhhg8vQlytu8f2ul5O51QTGD4qSOOKqxx3ZBHJ5Jc3GEJxJ2fXYA47Q7aZ4dye
vi+n12O4jA8YgIrbw1PjabrWFEbSnrfhnEa4l/QLjDJutGoacPNmudD52kHMw56H
Ge4Hv8/j/WyI6u1XgPDcA1rcG2e23h83zsNfVhxqWSV9AOkj+v7l42ehtKYfY+kS
XWnxoPCDmtVsuyQhXZ3+3fQBj5mX4tRFsTx7B91pKH7NI6LwTOij4g0JR1FJAeF+
xqTLPv4SxgDF3S/yHAbt1IR7eUCdFNk6TXSjtXXX6QU2aHK7f4lcNsgdPDen0Ejx
REB0uvhGE/YCrrMglyGMwk4CvMhs3EyAtXGvIu1KWSYRyAETZmsbJ5wVqrXREK1i
g37+YkH3rumjyCnXMsTAG8sqkfMltQXyIcRDaSnmobtEwQfIu6k9LqdQBI4ojo6R
iKZSq8Y674Qd3Yo6xq8j9YOAe4bC346VSGo1Qo1bvC8hSTwCKtQd8f/P+zPGbbXX
c1AGNFS4dMeanZqL9c++lVjraRSViadQrjf1suOLGsD103cAFNIJqj3tAGlSnR0R
uS7OGYb9qMjcM7pxz7GwzG2pG90S4FvzL5FEpIYk5m8DwXB2mynEJJqGon1a4Ni9
/nDA8NBaXEyD98kkg5ddxfjjgysWyUro6+KBvtx3e+O988PLxRjzH8x8sH8kskYx
mCnihyKF3tACsFKqegpN7/XpbBlrVUWPXoERDwqGoGlJ6WW4AwcCY0nmnOgU1WFx
ONZf95MR35viOo3P5LkTBsn6xbeQXcz3CDeQiiQ73WV3JqaOdi6gOX1cxR2N9o77
Kpon3I82Kb6pe4tnluDE1ZXuPQ5jtG5zJQEVis8HH5oSaHC65DbLcs4hqs+vlAyi
HCYlPFO2TY5kbESqYa2uHOWghI52erG/gZNowP8pSyouIfLacuqYmvy8TTAqb85h
wWzBEd1txYav7oK+L+DGtRB6Gu6LuokrmGjVx9PRvZXOH2eXUn+n5/DpmH540CdN
xiv5ee+7gOpE0yA5n+2B558B6aZlGOyohc+OGeMkA4KMU1WoGVyqffBFRxMjkLNu
Pashofm2+HueGpb0ObMST3yZbmCi7YHs5YjikoKO30QK5Mwe1i7kgfq7/G9TO0sZ
4LQD8oLSXJ5w80NXOmzHxQePDtBBWeBx6iFJtZklWjvqHhaOtFpTaoDJRJ+rAFRS
N43mu22oh2EPTWQ271JnkTAGq5efiGw8roMidsgqixMo+skl4X7o4E7rk2Rcfh7z
JaHDADGn66UE3V4qSEK1SHjDLgEInVWxWkTVaeLnGZXXb64ajzQ3qSJf68K5zkEr
SgjFB+cOpUOTYaBKJyg/LVpsOijKKRGWFAT1hZLwDJNvKVHMZFTVZBvXfjQO/vkQ
sne+XgGTQ6FYRj+reHQjo0Z328SfddyzGAV800gv1uCmzA2wtXjC6t6BCkw9bxd4
YRhwCnz9Psvoq3GN9XbHumaF79533SygaIXxpkdT9v7IKMJ0cudjS2+AqliCVIef
DYCME3HKbhD+BCODH3LGDJZWwfddknk5nivFqD5Gk2a3zei0RONvWWPAP1q7ngaP
z24Hq9Z+syD1E/nU8jFghcCvIbR7eNFqpaLlO0BAzLOQMy8+lkqBkWqxkqEQlldD
3JP4buGnu+bDVtidOpGnE3RaDsmw4cQVzhVgiNnmxFhLxwgZGPqEeTs2MomQ2FiV
sIm2LhSa5kfzeaJHZHD2pJR+0aprGVe9VG+jBeiHVGHG6kB3pkCdRVjjm8kCR1h/
8TWpGNGPGpXhCKSuTruhttAAaVl2Glli4aGpZ0ZF/IAD4OsCtcZ0y4/lKO8WWGT+
O7trK2jP8PiDTaTG/MOlr9v6MnyEmhbxBjy0EaRJuLRyXORTpZUKS0HhoUn9gdxl
N/H+V+5z7eKpjK+ingQD75/swwDEXeCUGbgG6AxcTVlLM0y7NeRX9Of9Fp/O3mNO
tL6bvQFoMT19Cg54TwYW1l8b1Q/drJiiu4d4GhIn7HEUjdcRWCgY24CfMOJbqjGw
NAnaAO72+pJ4c0pdkR3nLasdhZVTiuY2YUW5mV65zzLjD8Dyk14A97kJqd1TXIu4
aQ3QDr7Tmp4XZT/3Dqg0jKVl41oZJYSgIzuUlTDzXoY4DV+tbCYLPIsCY5CoDHyq
7+nCRLubM8SGb2uWM3XsWDx7RfMg/Qjc/Nd3RkhlTIX7rdY4ZOnOG2ZlIR2DFDBn
qgESpF5ZMlCAWJE9eqKpL3Zomrc4dYYiF+ABwsF/9bIEGBq98zxK5fWW1mOlEh4m
ciAbw8hV9WjP5i2WVVzWCpYZR8HOcHhZHrA4uKCvhQUHurjXlu686M+tWA9L9aAY
RaUOTxty9XPg1CuVmeGe5ds8EAcmSY4ojxxAgv0u2n2o7t1ESSQpyE2BhMuxIEqm
vxoffs9ikoIP1wwxRlCrQSltVRJ31tDL9+uGRpra22Hw1PQAwhebU6ON1sYk6SRZ
ZmhtLqUDV5N4JxIjSNvOSciBFOS9BKu6LxYJJWRcXxpV8hVSuIi3cqnp7Gk327Cd
vIXjbyrXxIJYHtjYUUZh+GGifwfEVAX4tdSKb2LnSflNeQOpYZrty3KvTuLvSsLM
n3NTfcoUec/IX1auz5R7+9qv4FsudAfSiYr2Gpsm66W37BsQm6ndOwZeMSACFWK8
dSxguO9xlpp9P7Uevzg3cPTs6f2p0dZEmg/davyd9ie2P4GL6kTzrgEi0bLdNT9C
IuaSPzxoJqLUalQ1M5uy10W+x2YA6WYkDsOr6p5Nh6bpiJ0rHl7IgbOa6mjPTY6u
xf1tXgIVqCNtJfA4018VXlM2l+5WBFNEKMdTcdvA107HSEu0mDJrPsxFDEHyh6OJ
qHR45nlEEvOO1fhRzaJIdUqKxLXsCg6OELaWsLn65axoZzjXE4KkjuggrINGz9mO
NUtQt2HmnBRhjTCNX46l0LytpqzWxjWFnbE62nkqduwBk3TP8Ct505bDjvI8/MBK
ioaaeHVeqa1BexlDAhSppDysASlKk09RmD+Fs11kFxt7lwxJ5O6yZrQtj2kRnEh2
udO7x/JUYKjpmjutBD1VDwvIH9qZDRe33C1e8DWCo6Z+IHS1mIvVCv4kJ5xQUZmn
5+eB+pzExWQ88RoDzdNNj7QOdz7QdwdLHodW6/iH2vmTxX5qN74IIwLLomI9LhZY
gCSadU/GYZ4E51UWeexY6miM7qBQ/7YhlwdH8u7ZzbKhQ8a2CX88BhZXXjxFOrvu
iiejk6DfBF3xaO/jJhZg2PAGY81k93e4iQTaTuG060nAeY27doJAGrLIXbmyFMUA
6DPR5vRkvCWDKwRLkmjhW0Wbtabx8vRtUGgFhe3LpeIgMcRtI1XTGBg/YwirAd3p
b6e2Ygc/495Kt2UYXXVGk4LwuWCt+UVbuFDugAT0qMtEySb5wqJBGdyvBliMUBvR
DZMKCkAvjK+qbg6yIbJoUJXtzYNCUr8v+wqYlGkReCzWwMjL3/aNvhMNF2d4akz6
aN14y471AvmS8DeJdoDyyKLgsBanPjlBKCtorgv/oG4mT/D36Hb3nc81VbMuRXWd
3kkIFtNsNMrAqiDvP0+u7hqV9+qjrhwIsvdgiTScVgqhkC2/thtomkg2A5Ta6oaq
xgeFC4s5UKVma0rhJ7ByeZtmntInHWYhwwov7E5Z3F6diJ68eLftop1t36Jh0hRH
7tX4AiBlqnpBhAq75FljVR/N50WbbNJRuHV/kJaMCekF850P4VwxkYncQ+bUXQha
i2/pg6fQyBG12PC21DtF/RGB5h+HKuDLC9Qqag252JOtIoJOj5pTyhQsV0DVZIYr
hRSdA8vI9Pvemqx4cR0BK6nWJ2aSLi7RPA6Hw35pe9doJgKmS5IyO0rRPokgzsAH
GxkGm/nb6TcUWvHy72KjvGvRk6tSwvEf0+iXYqqV9OZTYjyo/8tLJz3Naeo4gN9z
NVWog+5SVAqAjPYLJmXALDcQQbBzis/JIDgaIf/TCbT1JaT7h/I8UZa4aj57nIXJ
OyKyeqHN85kT7bWz3jXY1r+9208r6NT8hD0G0PrPX2JvVqYtx6wXbbGpnb0TPO20
BDvA81M0aEuPpwO6uUU6K9NnZ28kGb4u1PhpF1HfeUFEdEeCSGxF5Qx+MNvSNwU4
/sAOXX4C9QOh5IjZWOT5A0Rz2cXMh66yyZ593Wt0PCu5V1Xv9Co0odFA0t1CXoWV
tiggYYxJja8DIfAEizGfa9vu5XsU4hiQUKB8EAv37r0eRhnA+ei7vsoQ3sw8UTps
ltcMsbVvURz+/+KKmWajMoaC+HJxARy7ZWTbBgKO7Okh2cIkkSfllM5VQz52rRRr
d03P2/nEwI7Ovb3hjOqtZSURoWQab+dI8533M7uYFDPe2pe5NQs1cPk/b6wPAtxM
zk/19mXZnWOWeGMdgklVGe5+iKW8FsJg8VoC7Lf5XmVEp06R3oHX41dYoiQ7ibiE
4HpnFZ/eAe59p87mA+oMRZ4objr+RIWIUIw6Me/ZdnG3uOtpZjuTcCiAx8/HJSyF
bI4mj3nET4nT+ZGxWEJa7bavqw98AUQ83vMia0PSnralyLiX9WCGUtZZwJI87U7w
rM0BuwMJjiTPmGEoXQig5YAdgg4mEhqTBZP+qtg8syoMeYo0E6JSlE6PlY4z7N6b
zMyxn+2SCmjDWtKDmVTp5IxVw2JRLIB4tBzI+x0WEF/yITeQKt3ZH3rtmiO9rjqr
vLikqaVYmbBHriv6tl6HyVxO4gv6s7X+owwXoX9AsYvy0O2EsezOnHxnVQCaZSdj
eiF8/KsfnRqOpC9sPpJyp63NIZykr41Sx2w3xzvRemY3PYhoB9F+FJG2hWLItPnv
7cnfhDuVbkpGp7I6PfCRbFLm/4x4HvKxtMjpY4aVllgNlOb+oxzh+iGORdKWvX83
uz9/MzKxfyi7HxpceJpeUoaOA8DZfV6OPVL3wHmx2y/RrCBf9onXpT01i06Tw9BP
4c3DgrJRnaTjg/PCeUJ1PR8vBDqlmv1yQZH7jlIdsUyXhcfiYoRnDfSpIsXut9Gn
13yoGpdGcdh9itVruWrQIRYp76BxycWInI4Wc2OxRtN0fFZZurepGz+scGIS5sG+
uGbqrKUOUS0UmByVd3UrGeWssvjMDE4QobYxzm6ZJS0Xqy1clULFlLER5xErpz+g
C64Eb2hp23wL2R6naKGjniO7/2Mzp31AsnL5TiopSyqqMXiyk2q2Fd/EI8xblum2
HLV6+rAh1LKXrn5/gOCkx/r8vfyQM/3dFAg5q0aVivVqITj10oidM6vwTcM9Oq7q
sBbMw8rpiRaJqPst5b0mtN84qVvjweOi3AyVg4AlruWZ15sfMIWHvJs1zdBcG51m
8knjAr9W56yb5/edt5/7zCi16i28XJBKHSv6mGQ2y99KFuAV2s9jhR/WTfAepz9F
SaTc19ayvH2FV3aMFvyZU8ImgdNT7kTVxklL3B1sSNjkwmTP+BYZP5cpnW4Itqds
2ZwIqrIcmMT9QnN8j44tWz5FhlLqVu3BR22NFyFoT8SbjjlufRRKXqmEAq4cLoeN
n0pSgRxnSpWjmEC8HL/kFs19Q5eVy+lJlm2wbe7OEC9qvq0s8C/dWrUB6FCamo0g
3T9AG3NAJg+fUK3csXxovI76O3q8We3B4QsYwY8jKsyLEz+l1YYgIwriyF2gP8Nc
0c3FKrRk2M20h3Lbnn0cYeshjc+gBftiCgcRJwqze8QXgekX7HHfZKNLhNk6Etab
u2lBip6lvpyTCsZtwWeQuV7kBSKO3jO0NpXfLwfs0OxLrgwzsFL5H12kP+1xp7wj
Oq8Rt3K9v5tvLake5C/Cv6cDxnhAoDdGLvxs3SX+yoGp76KLZsLIE0HNY48H87IT
0zoxr0DtVjvEk412xN58UewAHStmhdNa6JDbJYVYM9dHXT4+lb9KrO07U+gDO3oF
fccR+zORhd/l75DuWBi103EZDzPaC08xynSrGMCoVIuL6Iz5nufRKdzyiVbsQBvd
qp+A/R3PI6cdshUx8RmsYMIv75w3VcyYDu4cmkxuUBeyWTJjAJpp2Em9vzxt4Ovl
6ov0CPxS8B1RpOm7m4JXHMQXi5vwqr9AH8O6W5hY7+5aRR+Bw/3y8uzoDit1ngHv
zUrKes2MXLLyBQKAqMT8iVGiqjRtQXMqihVZD9yl8PNI0EKxsbO/wFp9AHOAPuqQ
R3Qrl8Ny4ibWMhZcZu8B8+qiO867BTMN3XywCwUOdXjGh68vCLitEO3w27GPFbz3
SEv2Q4qVOWBKZ/CAkBoSBASyd/nudmU2bqdQ6mfsGbYA+RTecEYkHjgf4Kj2YwPC
v5Z5wiHGJ+SbQTiBzPeR4vbch8f5fTsdH8aNXxhOEUsFWJ88/Erba/VF86LUVk+s
XY4YhZmu/QEDBHS6mTwsvyCsWNriTt1Ff9WO909ghjNEraEddJpYR2Bd/aFPa0BE
i8Q+0r5C67n4sSQBo0nL3aEWs0dKYKMJTs7VSCCrRhNckaToGDYa0wT/SHmIAnwT
OOW/qmLtQQcHt3jyXtpB/BspqqI7XlP88WoCdfFzK5BmdcDTpqi1/RGyB+BwGAJZ
4WtEqOjiBHCXgPUhK+AeVmGIj22TNqZl1iPX5XYMuwFOMCWOb18U7jayTidP7wut
IMhqLL0DEKa8CAONDPh8rgCS02x9zoACgqF+Ce5az6eKhhcn43PkN7+hUpBnJbd9
OAmtFkBwDShoVWSQyCM+815WQQtOKYWMv1TZcScbqHHownQY1G8bJFtQDDkF4p6s
Mlekz/BzTzP/Zajr0WTNdwrChcF1CYdWT40lbzKtyK3AqRBNL0eLne8rHwAYvefI
n5BZJhNoAnCkPOD52AkrS/zUncm0yGvF6di6qKvjmUJoj8l/naMW5C4vtR690vnT
U2hPcuK6xOSSeyJkJamnsuiuGmSJESIKv8vbVuuB2XiEt7VpIkoS5SplhkCRmE3s
a5f05ompZTymc4J6wD2/wQfDn+TtErKcyL45HgsFyb51kQ47jAS6B5KKeJcR89AZ
UIoz3Z5IMiCnRkZ+5aUnJfUdzbn9oJzSc8LZJFfZ5vxnJbwxoINDZCmHWZrlskX8
odJXpD7eh3oAc0imJb5OOItlSFu90WGja4GLTvRIzCiBc+Ua4EBVxMoU7KxYvxkO
mZklnh2xDsJ4TqJvvT4kNL36J5S86E07RBBCh3CurZrVuophGFpoGawlIugnYhQq
8JkXx8O1vdQ0l54JT0yComiihQtTi1LCeJYcyYAwOdGZuzUgfOaRZh6/fjQB10lj
E4OGvsdtYDl5ikPZ6BON4eDeGsutjSauBC//asWUjWXLkkGQUhMrMepr4NJFDPNh
9zP9YYRxQfzqn26BZi92w9di4/llr7ZMHKU5/OlBuGBnORAvZP3GN5t4UJ1QfHLe
UGlPijltb773zCiexM+jf5IQq3XxDM4QKom0fwV33iA4uTTBAYv01efB1nzyw/BO
bMaAuqYxgbc+rm8K2rI5qX+RWmIdPGbhm+6SUfywSayVF+Rxrj4Robqf+0raAX+2
4i99I686MQmR8+AWPYhziSoiaax+vM9Z8WAey0s8TCrFcuefV8rr40LiykwEhCmy
oHG/syb3TwUZic4fBsqYqQzIu4JeZxnHvl94d0GH4WhghMwgRe361Kd1GbY4aDNs
goUVXA1ziOIPFUgPpZU7gNlBB8/bXHu/uSRSp9AK4kAbaZSjOV0fr8+N9OWYh/V8
mvOuNN3LmUoVPzmX50PvKS4AnbYumBMoDILtnZ9d1gRm/PXQ4x+/ELKAVj89QpG2
i8bIpEiHJChxFGXQ/zKrtUXtc5pqUX5lknF9nvHSJeYFtnrsMxBDTyMe8fY16a6x
avCjJgNgQc0eB7+4abIx4plV6nkIDsBTPyXaIYKFkIsRJoqVysswG1FkC3LeZmBj
zVvUROSGXt2c5ydEgY3cpNrp5qbVYJ+uP1LU8QP0hy4nQ8ExgRixLC6WnSuRUKEH
gURnhk8NSIV7hV8u749SATAT0674rhw+iodsWSL2ndTdV1NbGHrRjp8dRs+byw1W
pC0dDXN8Fw+lyNstksHJuGrrKTDQQ8fLlGvVV014NEX61OWIqu3dFtSAKZQw/uEI
3xfCJbzTOLUjeI9Yn4M0/hhfIJ6RsWg6bz9/XLjwdxIDUC2+uWENUUHQKHSvq3vt
J9Co0M+qo3K30+sGdcfu1AJjV2nVAgVEE8q3OFV09yHpwvWCuUhoWvzFBTZdzr+M
geq6Ep3WzRyg5HtZd7zH/RRVhfRLpr46h93+HmgY2Vo3fivEaLqNAm4m30iqO8do
1L7RNHH0SQgxHUtdKIcDBZpN5UdytKzcATQMSIUQC6KeyzBZjUoMgAAZF4qUy8hL
e1Y/EmJNNCMFVsHy4ggh8vDqYyct7UWm7yAsuQwHpupTJV0lQ+XGQRjyzgaY64I5
V4Kazw3ME2OMCw3WfWw84RIres9g9PXtTo8z4jN4GO5EvbV/6MdbQlASOorw+rR5
MUC/ofxlnDHnnJ2zpNtvtFoYsvOkSPPtDfac0d42A30eS45ss/Qcf5AbX6UrHCG1
wjXke/FGbtmgRkTzwqhL/2IUi/UWY8TZaYazdYcHHzP2wTXwM0R7kZNYm8a32YND
ZWh0m+6lr/Utq58CLNrCpyE22mtMBTuuRbQnHigr1AoGORJfVZmnjiZZ/EWTgOpv
IcA1tgao7eGXSFkT1N353QfNKVX6BypjuTdKnfMghAofED2N6CNbIw6M5ld+jMzq
W/jqSn6PPD92YtEhIVL/Vwo/tyGKb+lFN2yjuh20U4UoUdn9/drTO/AwyzfUB4z2
aodu685aNs9aQ4FcBUJB3+q6GO78hUjiGCMj5FF+8rdxbl7TTOX41bt2s1TDotCJ
swToLT2VlRYaaQgM+gcvopWYCer94AoS+3rB2QNDN0/8lzon2OfyZe134q+IfB34
dKJw88IhQ4cIxZxFI4tsGl64YfbZFsILGRXQWyxpg1MqlQRYsAytxRJy3x8uuwhv
2AyUbKNh0tpY0umc1T6sTBaoxPzQ1oQgTgMLVe/zK9Lffo7mYi3vfOY9N75L/HXg
zqdKGmQBHa/UJWjdLbsbImYRx79gCqwcIzewzEdfELjCVsHXg98MaDTcxxB13uTj
hBfNT4fxSGh3lVl9EiZHK+JKztdVFVSqyGyliE5VYY/Rr+wzpvtvnd+JLV2y3N/8
pjiYRP0aME3vmXBbXclgdOdQJvfcxnO6SLSc4ySKXa1YM58Cqefi4mMYDnV7W4kv
/n6H9hsVV8zo5Zxy07QF1P5QtUehNnyFWpxCov6bSJkDNJYN1J3ybUZQJJSm2xcr
ILUH/I/DroddDXuf886Je0anEUzfmZzZJ5XExFzdsaSTu8ipiw6xqCqULSfx30fR
6AezHvnAjirnT+odlkrJ6/blPTOhT+du0DzIfDpwRBXTSPShymYQRQhHICwMCYt/
5mBC1S5eVtMBFsHas7099TNedCNBelBQWoWXPVu7csrqhhU1rXwwjEFO5g4OVgnJ
Adm3azX4kXo+ybhSD0kVVuoFxc+AwTGzNSh9K3b5u0Hbe+k+Y6CCaA/vn5PbU7Lo
obsWfBXp+KgVWpxL6lyyJOnN4IDgptzampz2U/B+88mtQ02LBMaVBjQ2sEsKwpy3
+BVWnPWdRhnOhASsfrOipcscnuZA2PbhpOtrAYURV9NQgKXD2UEtVJUPAdiWyxie
T1yDgYyiepdfQuM2cEzqIED+FY3HtF4K2pQ+TAYUFYqkjRwKOmRlH6j17+dAe0hm
R9n2Y1sAA+p33FLzmwPwEEqyLus2sZlFKU9ctZLIMnOth5v+e6O/Lqo1QXBa6y91
UKjc3fAUpZJEWJPvzyHRAUT+YzzWWzkdLSz1twkvRB3Gp83dPjjcK2aaMDrryDH+
f65LXilxQ8A8XI6X5PiFYbfBf9l4qLJapXCmrRMUegzl7edya8RftXld0oBHQIvk
yg5Ysm+EsEmqrfZDF6ng2zMcIbBce/GrsXZT7UBhAaUUpfiHSSvE4QEtoTz6yMgo
lSBp4/xkUzU5DAu4TCd06ik3U/cgM5JrkmtmD+sbFIuJNY6UjbPLRr/Qtqzag4in
nV4Y1B3s7T1wmRCZvUg7kbRXGZoj+c4TxCGkpjah0dsJJcm26VUKO3kssruY64uE
l6OB7TdRtZIxgwB3f0/xfr4mQ0vEk0XOHVWcl7UKLfPgrDBGbSv3imGvKTS0+xs9
WoLb+PMOUhAHjPQAATwe17rPx3Xr74ZZRdDhg4AGgLkHDhTpTg16iDTtx8RnCAVt
kmZTNrhgS4MT7jWiVbSQ2TLE+c7OeD9UB5VYmDmrINBLp9NsvLC6W3o8k3VbQ4M8
sI8+o/xVWuN7aHwUGiblw+m7lUClHQmfPlCvPi+iQZX440s7JHfOB9bg42CLM8lK
y6VEY6jsSttLMP8UJxCpIY8NcXKW0OmrdcFMKW3jVQhSeYDKBpSIDKw4Ou2mItfO
Rv8OvSSFNfghDsnKh//izPbhh1jA8QsBC9KT5k4+91KFiAGogJH8LxYNPX7nEafV
FuVjoKu34v2vPxKgQrdCPyD9LJGc+omUHR6GerBiw9Ps3Q4J9k34y3EGMKVfHgLU
z0IsoR8VMKkmuPUCP2/SJpCa8akDZueaOpVRMVCwvc+lUzLkAJpHwS2OK/t1rrJt
6ueb75sTR177vqIh3Lpi1eKSNyPHZXMWWuLtFYKYG4DpH8GO9jHfGjd7YdgZiJu2
IuXg99885ITEwR1UEZUIEMXiZkxmw+Jy70NuB5WFA7MACMcG/8+I29Oq3K3guCxb
OzZPVZmdgEaJb6Q+c5cqpC5QFg+I/nGtS2Y8/7QAsMS0hYYnJthWmS7hQOkNf3mD
IcXIsD03/zT7wUBiivk6PfqUvYPwoc75lLCJnq+IXXBg4G0BpDSOQBAHORgHNGBw
zW++7UX5TOgtNj129zVPbdk+63WPUE90zNRLl78B4AMpxDKdM2tPdCX6AXtKOh5G
03QoAdjazm/Jf/uwjE9nZSg+SoE42HdwcpZbl9tqYua7fAPMZPeZT/Af22b5QOfC
t4mky0QztVPVJRTixGI5qBl7KLGVDE6kIYgpTORI9DiJLZl38Glr01u4cOMAuLDz
XYeQBwbVChSrMVb58P51CSv4r+agDf08y2goa7YPJ8OwKNf2/BC2iJjbDsB0TUbj
6RY+18q7GBAyoec++P18ACas//PgZFclxSkdQfocwod2nZXTSxJdRC2Kt6rD60BT
0z2natbFSvmFyCZ7zY1SwWL7a+Mo3a61xXUVmV5uEoKESg8/RAGDaBPkDPNUoS92
4IgxpWic0nKwZyNFqQlEuIZlRnU0t/KG6ezpN+BTFU+HYF6zZVK/Qiozywt17s04
VSHcvSjazew++UYr6M9Ifu0YLp8IV4hTT+6i2PCixhxCrigyE9A3glx89F2matSU
oXF62Quw3uS4ubJryjYWlE5KY8GG5ZZCH8pTWkDD4dui5xRvjfz6lDWxipYEdtx6
OG6/0f+mesUuY5xraIvsOrBDKEUA6U3fowJM4rkXfJzVvyz37WXKiUvmFF0Ju8IO
LH+IWcw5R0cdqIoXFI4jqjuz3yPO6GHNbXxKJLBeeSwKZkvLS88dHV90RkOou3I/
nS5db5V2Y3PRiaFARJmN6u/AT5+578l+KOEECMzPwKvh6D+Jz0g8yIeWa8GVBrM+
CLumovCTYhB4G/zF4VidY1bALWYGj59Fo4VDvYnruI/6g/UAGjS0jac7cdyJHfJp
cKN5XqK4o8XJ3TMKPcbsZ5rxmOhmDFLiemyiAfyjZUruBd0KpC2G1eRhh5vXdLvk
rSY8WLGbAofoZ1csyJHUggylFf8PCapKwCJZUm3c1EuKsd/JafYv7X8wyd3TFP3J
jvHyAcgcXBKOp9QcX4gYmvNNWqHaT2rmdBORtKIAGCAyCE7B+dDz2tpqvrBGg/vg
QDpr7ZmAcPxU0MvAZwhkzns2OiVrJ0w7gS285WCw1uZYPyxoEp0EWfYlLvbfBhWs
ets5onuObhho/hNjS9S4dWsWkKUrO+TSwV33aRGMVi6Mei2ryczquMuRipHUteNQ
IcDQ1punL7XQg2G6AoXwhCedrl/vSCUc/WT1yYKPRIOCS6a7VMy1Joi400d712m3
4HaefgraBjx/1XfAE8PKEdCXsF46NKJAkbdVYSZsspGKSj0j6Loy1eAbOH/1gySa
uosT1g/zwJcsnSrDqaPku2XE/sq09s2bSiC1pscHxS4WHussr5FeFQc2kE/fnK0N
BkToHx84I4mpONo0tMeRwxv+SSvYUF0+pSPQ/UhXUXAB643J+deeKmXLJxPCCvSh
DSt6Qy0EkXYFHw4+59+3sJVZEX5/Mi9kESb54EypSrM11RvQrTAykkccMI7cDfi7
mDFZO6DpOUuFncwdeGkO/sEWpsk5LXesmFFede7S2Mv/eBmAqMlLCQR72o/BIpLG
JERccwcNxpE13uOC9MZXxVqhfO/gdAvGQkhsbg9MkUQv/cuE3P2D1CmXt/Xtx86s
ZI36ifOv/OlTMWaWCt5BX7m9w3GjyIVEl1IJ+ylptZvruKFzKOWXbtj5xjVkRl38
q5ezlEFjEzWGR7p7NqxxxGT3i7sYbjQmvEWplBMpfXGb/oP8oKies8EW9WBBP6ds
b+c7s74U5hsIC1FExTFYXoEPlPFz7+THBerlQjMCrq3EQgR4hqDdt4qiOVyx1Qcd
GuXW/QW4XdAqiDM7BqG8VmowvMVxXZEELonU7KCc9LBTkV9naRQGZJEtagRceN+Q
KvSm9BlvpZxe/NfCLp/vgcK71/+8rvzTAp1S+YBuAcIgIso+7E/uIN0yBwPgb9vv
vrXHNp9cHeWmIuvtuSOxML+tfwgD9szsepGUc4FL3on2Qt+XtOhoCRe+1zQlhRjA
JFDqdZ1yB+c9snwyX3bbuUOnv6+rOyCbTCLgeQur/Bvl7UJKUOLByXV8LnT22fs4
wxT07cCa4j/An7kHDs4+tqtUug8h3pIejRHSOrz5NG/yoGUgvlhO0TpuzCSUIR20
jEWrmbXiVonSkmbU0z4jo1ttf2OuR7GF0X1u0ITjTi30y/AAOXWrsJLIsequ/e7Q
Gv3SvztVAnKCJAVGpDlGWEexZMwA4yDbXZk96LB/K1GnqeS68nL0zQCQVnT8Fz43
N+yGTlH4LRQ3SZ1ia9WOIzLEScvh+ZRWomuB4uyFjYTbgqpa3NTG7acVsP8mbtd5
Db8F7NdwSO2T2aJ7XosY70OxfdeZr95QlOKBCT8zt94vJsIDqHu7ZW7vOY/dIcOY
Mto61UFB5GgaAeVYYa7Df+UwsQwZXhT5tGUBWphTzJJLFbASDVvit4a6EeiXHFYx
lcQYAAh9qnS+53pz5g0D1IFmA4OwY18drwCfS4+KdlhzzuQQQK9z74cCExdlJpLr
5sYR+A34/cE67gf/8sJmsT1fNLhcpAfPXjLCJnx/POOU723T6WUP8IJhXt8HhsCb
76ZDcX/xH+pbrzhDML4X6ZXgyqqKZiLLh4VPykPNbTs6+n74ZdcH46dJdErqnwIS
CBDcbuu+9bu7++v+Y1GvVxcbHQAIRbpWkDYdvbCcR2H8AKafFZfVpnl40sVdOAgl
4hzbgbINZYa+2V/jK/+ooI77aeAk3XT+0gJopPy82WJZK8GubMzlnpYiyXSuQ6b2
ekO/FfJGOraBISMZBPb73tJYPPnfNQd2O/1r86CZkC7060I+/3l8rJAjoqbfQU1S
sNY4Z6aL/oPnVIp21le9DmTg8l31Uz7EQHjxjjoT3D9kt66lWS5qwIBRUXAiH+C/
tvLT0GJdtEAsU4jyT7OidByV8UOxB5LBEfdsAVPBuVI8/5xzwvLpcDa8Nh/tqIu1
VriEojMOHRX1dLMGhTCYNG9a3vx5+gLYq/ar+sBdJyEkAQr5rkPiW/3XjmeEDLwJ
S/TO5XuJ0f/MN4QjWneB6aGc7fMWIo+s48gaqY2N8oIhb3ORgGpuevohDu93+e4a
iscPW3Mpca4TNwL+D2qDzEz1O90zy5kYKfA59UMh2ogi/5AWjsphklWf+0/oB0pj
ESPKC3ZI0Wn8kWhauwg4cJfFa88E/jvmJeqENREwSX1av6pyhOmaMWpr+TeG88fa
seghFifZT53iDfUQ/TD40us94Fc7N7jb7aTueUcEui10L1vSungBgpA9yQupe2Dh
gROAuLjZjixWd2BFXutGvTdAU1VUparhCA0XmPbGX/yJrR767GFYTfxnFC4RkWC2
SmixE8PJJ6H3aVCyLJPOeUiHvtppLjVouCCdXvs/vPkXoCADytxahHU4RisPpsXO
5T+2+whbbJIpaBId4xfAKlzO5hHuAfJnBHrvKZYSSxhDZ4ThYJ7335J418rYqYz/
7hcYy+cBzMz0GNSc1ZkUk3iV0FNmV/pNBumRFk0/umn5AMpuRtwV/EbR2I7V5XGs
35Cno4in/u4OBvc+j8sZmQCaVh4NKiTiRx1vxo9kjNMhGB6RqUN6z+EUOlirsBTK
BgCIINbDBuo9AaGsYtnYwuf9SopL78s/Tz0WlramdqWaOtOWlm3CuxsIdyjLxF57
714CNL3Nu4k7JkaT6aj31mvkB6YYzUvU/WMqRi/G/soWctIvhJoHz0BKWkyGdTja
YaWYTAEcQ+ZRyFcqNnLU6wACWe6tvPwKstyuGmRUSmR/jkH/2xoDFPi+hbCI0OxP
Cyr4hoelljHE31K5whJ92fVmZEmdoHNYHRbTXc9tQkGTMo4sKkkAu9pW3daKmm4g
eu9dCGzaEhVYzfFXmX0Yw7dZc9C2y78GgtrxF9FQ5nVavEYB3NmXhxRHqzO7M9nd
FVxHmpqz/Sz9f9jOv2jFIwFgk5sWTviESGe9TRxxJdnCgTSaxeJGpRSGXVogp7MO
V3ffgtnHHBvM0kg5mCD3HEL6tSqgyJxRSUK7HPkvUalqYe/hLFP+mluZhlCVqMMY
EHPwxpki53K8uDm8oBq+4HT9GYqrpZAKrSR9HbCainWjMhmtRjJmOKK0dBe2y/1G
Xrn8XDdXhgNTYh6EN1Um3SmtYxKiR11UBhWAKPkvFwSzTprwXurn2NnKPyCiyAcL
6a+wzzD72eUIPmMcmnnN7S3SLANqwwO5KsZsAovXJioLFAX8LYUjKHmKH0+/Uye1
Z4tQZCSRq398e+VYdcu9ahK6edYZclUjnzXmcEwoa7trgc+B3TBxoaVACCn7WouW
CN1yLlNBBztGqaqLo3E8t44avaa73d+avO7LQqltjGdA4hVTC591HG6qoaYtQets
UIkrX0SPaI3sqc4Iw1m2HQF1qyO4Aym+JMLsg4cuLXn/WPjwtfLnE7xQX4GxHSs+
HHMmGZWRJDf84dIcwKXCcc3z6UT2ts/11lEVuKIZ1WzlVb0ZLVQsEzdh8mArbh2w
tVZPJmxslwhNWRxzjUUDBMT+TIdL/nJsIOedX5NEVR4s4wO7wyR20k8pcNs0AdJI
0pPNln6aj8031IZDwk+07p65uWNBZLCCaH5RsEzpvxpuvKlTfSr2Lhu2txKe+uLb
/x1ZrbKQ4nw44bc/g09wC/ouO5+um4FEBw4mQP6MyMZikWXmyaB2T7EApl+F+3D5
UHrcmkJsW1iMv3645aUYshs5HWaL8NBXyDcsc9M/ace5hV2/SNQpBbKJlM9cQF+P
UCTBxGAt2X83Z5zLXJaALb/ip7AqB/5BFNTNho9OQxTveLyAEtLvkBD8OqK8R6nG
8JfMnmMTisrGKFtmrqAVz25W5o625kIhTm0nC8v7AOEhlBYUJA4T1J/gK8deta2O
D43mtGbd3eDnqBOrb4TMpXwm4SYEN41FPRQU5C3cT6Taz0rHn/64ALpHtcD0bRM1
gQc/2fKCEU+4zMIS0QELaSt30iwuvCsH92j12+CINBgbNcSODVhqgDB3/NeIr/OF
heYdD0FGNe170ihPYk/Oulusyvu1blam9XCwupafTombwtc1+hx3F9rFquwpFCaH
GWYOFRhcNCL3JA6/Z41l25maddXrbXwX7TsUNLGtacPz+ZI6zyH7ZmYz7KaCZCdH
XYT6JsnqVgJoH67S/SvdwSUtEtTkl1iDCB9990nvHqq76oOYCwVr/dAncgfwsftN
303nNWKvlaVOx7jqNfgEapv6D2Qes+0ouG3B2TYkkFxlBpZNSledA3ToDdjLrJj6
ACCEaViGk1+I6Gpe35yYQuKWhUMJYFthl1o0s4lhl36/vQHnoiPRwdkMszBj45Ma
Ydu0iUI13R5gTWWxNADW/tNFrQOCR4rcaCpLVJu/IE4QST2kBWwZuVUFLWoaNYIb
C8INw5gfFB/VJUoAbfCxtEfAU+P2NdX9g2lU1jqvO7rKyO6y/NflJxM6j5hZHm2y
8vBU8ZzsRpQCiZUIWA6fh6wIJphaae8trtLKw1FDISWVmovuwVR1vyO18RDjiu84
PvTAhdK1DQ2R9gNqK3wmXCtps4VXeFvR5RZwpkPLu0olS+h9cgUSGREsDE5Fm311
P9j2WY5y61VFwCF+AhKV+hyFB8U0bHZrIgjdFE3KQkx270IpBWeOZuapKv9FdxXD
SJuUHhTHgg+01BzLmG0u06tE30hKMzEPu3pXTrGboA6IP8m79jo/pM1Z7WnE+I2J
YIg61ezdUiZLMH5/VuEZVDOr0Fyhoc46A18VaC7F8OXCHcd+SkwtD2p5+yYBiohP
VyjbodcCcLRkKIw9flEbiHbi4DnZdffOa609ugenX/WQB2VMNvl6tNP6xagPuCuG
palv6dRDCZHf+traZoXu/g0uzzxJiDcSJQoWXBdzcRF6AWUF78aa9QAIRlU9z9IL
FeuMUcw2qMfJ3iadYquopTTD4AHGERILl95up784VJdDpgOGejK2DTKMtnxq2gsP
dZfWcziYpoaAPttIJrGRW2Y+RuVqO+toxG+9opwFdyDz+eU8mZQCLi/Rq1bPllbN
pjfB+U1yLKQyK75EHyzDANilfgJX0mMyXCrk0WOvBiX1kjt1cTp/ruWc6ZsxrVuE
fkLK5s5BnoWdqcJ6zHWPcf7yI/vSPxglq27lFKpfxnpPN8agdhFOBl5Obkj4+j80
JEWr1J/JpvikNSl7YXKuTJsnvXokZQctBsw818nhO3FRbsf048hSFk1h09smnqx3
vAqsUV3wWEKzqB8S+cmyYI20svPnjmgfLYa4L9lhzUtyy2nqJqhh8k1B0YFla70/
Z4UbPHS4Mq2eSupY3BWxizn8MCD1zEwbKNMxefhdxVP32Qr2bUObbkghiPDazXH4
GfvShsQVZY6jcTh1Nig6PAhNtMC9c9gK5zfgpiYfqP40Zei4oiDxRH/d0j5wklWj
v15s/YnTAnbc7zuyvd9xkBWOu3xyjTFT67yDVIjA21h0YCHjf1oqeLSH7xTysCGN
NdiVrLfYe059FlIrLC7eqLKmeFHOEKc1cWPdaPbUuwPlCZ7O4xJ8wst/3jOptMPu
A/Phuc1xt+5gE6UiiNYjjCyCKm42LhCliMnBkSBIFaT85hfFcnXrmNNtIiKQwxIQ
jETuUajukpLfq6HUMLfZG8xLemu3kJEyP9uA5/FbUTew57lVzNr+pGQ2F2drqsF2
s1LaQxxZSc/GeQm5fjF6iepK3Iigxd6FQqoR8F6aXsk4PJ13PghCiwaFPlkC0FCq
UpIb0bp7xQFFryF6EU8hnrHKxtqoErtcFvvZqoTDMT088k0DpTtWGYDbAaI4ECqN
QQ5zFcDAhx6GyJp4lj6mq2Rwptk76Gj2FOJWxOHopC3ui45ztlwIG7+u2vTutOK9
KqiMByU1BPSGKVbFyARj/NOre4HaOLqXs/FI5g0F8aA51TWr2eyRnFmJMlr3U4yY
MKArY+rB5VqTlbH2hMA2vZ0SmzEiESbdGYEZY/GXDj2yDabyMF/uEBxQdamWBhmS
tROSBZo2460WLs5dJ1X64Q3D3+f9A2oIaBgiustmXI7ouKtuP7kVaW/MiRT8SAQW
ytZTcYk71lyNZcw5PuESG52gF8mYwncS7ut1FYB7avUfiY58wDIhyAXSEkf3XNOW
+yEazFK5gPnRuN86krqr2lONV11BWTqE7l2j3gbLV1YZO9tnkCBgzfaJeH7NNu/w
n4GxkmNkhLU+L/HKBlG7uzIPOTcPvDR6IBKUK1aFKB7hnEyErxGXBW6/uFI8m+WD
ROqdYUh4qL8UnrT3HL48CNb9MuDirBNWz668Vfoc1TzFFV9giWSL9WElOIhMTS1/
84uYUaLRMStay25+VmTJwgQr7g8PZppOoIxWGB39ttCOv2H+9UnOZll/4CNzS1ly
fNsKrL5gqEKdx4ElQx5gGGfwKJ1ubMfqZ3kt30OH0xr3Qv3AeGP7mJ/PtzsqXNbd
b1S/v0NsK4HqV/BtEq3yjbQJGvL2NWodSSKxiPkvnYyMw6kvk50Itw4cHwRMdShP
3JBbO3jFcFokUzZZz8eLmE4fhjl00NgTt0mnIQ0vPXoz6bMZXrP+/LaW3orq/EPj
lmbheOu22JU2M5RBxcJx6ZsE/kfJp6+tpJpOsSyYLSoGxvdlS0mkclrGL8y6Jlbm
JhRb88+FzD3W8dTemtHlJPXQ4S73NfiSQuUYJ94J4K9Rkx5ebW69A/kIEAwco/i7
ArbM28zUp90dL8A9ahnL+61SgSN3nn999qF0XpEkHFjE8GQJOvvIDkF6WoSniidh
U1IjeslCDy5lkSlUL1bRAiVzuWu8jag2W7BvaLGyQoGO/uFi3B/smtV6YaAik/gK
gKaemwrgk705/g8iBGPv3OdDLsuhbgww2tUTTA7ettGfxK2s7tzga1v5AxXxVbmO
VNjiByjELD7+pqZpjB/hfg0Bf6kl8joIuJe2zTi/TWaT0upYmkxsNPurbDNs4nbU
igFRV3xC8DXO/hlmlJgNNMmpG3IfCG+2CXbt/oGe717fGlSmXU/N2AvDnacCKq7L
mokWrPz+sNC4tY3ir1X30Qr7nXpd5S+s9ZNLtp2X7vAejKspKXgChoHmtJsjMTEr
UYIObA6PUFUV3ORlrm/1raJBjkcrB7qec7akfVGu7+Ozre3egULsCTlw01iZrU9N
ysi145tlipb0AA22620V+MTlvr1ONlREQmEUbNtaYojYJC3YJnJFVySbaL0k+VsI
KotPR8SM0d3RtGiIcYZepZy1STfinkOuf3+u826YBSBX7Bec0iCdFIGvfLjNU8iE
vFxip+n+NJePoEbeNGKeECKtDOYGPCQ9hh6ELjKyNH1gEPaaD7+10v301Ks/YZOk
K8pC3JpWhsc0NPYAAfvly8WjRCPfSw2pvDmBCLsSS+4UiIAMr10upQPJMJoX6yT7
tykrEIYpjJI2l09yj2/30vfGXZ+nihN/2bjva7ITDS6aPVIGurge8olbQKJ2qYLy
/YXvl5QpJ5aL3LIdDk9IW3EfI2E0ohde4kKzpodsmY2Jk3P4t/0VBax//54oWDEs
y7Vh6HAfm7XSKPRXrqo+wxlCPNDiWQBUK1paB0dcg0dBXVuMVMPmufgPNI4flv+r
NmXV2/L7qiDOiUBAnPRaMJqx9Qu/IqS8ef4WOG6S0CG4nWI+mLE8HzhnK03qPu6r
lA79rj21lW1CoMJD6pb+ppSrLmFAQco0MzH4uzU01ldh7j0Er8bcxO0Pi0BKbgVh
jQip88Ogifbtq8EnvmuNKqCKTpz6poLdK993MbYAGUu3yRVP5pTXnA8a5FHQEfz3
X9GA8ybTan8NOd577hKU31CUsOOBBSOygXQ6y6clsgzU8s7X9kT6fauDWwHAouQI
4lnrX+D64ooYQUWgF0J/ktk23QKOgm7RBH2z9oAXXCDH7SEEj6GHqirRSWXa9xVg
CE1VToqdc0mz5PWUdGbIC8Dmz1ZiNDc1r3Yx4xLMHIaqmjM2eeBIh6Qsk5RvX4nS
r84wrlKqQ+vAEmsEE6qOnJ7Wrkw0iA+er+Z3TueKPTTtjRwvoJR38Gc/Ikyq1Elq
Ypi1DzyPNwQbZZY9/pMLtXrmT4Rpd4VwUl5ANLoX50V1bbJWd/rrLkik2BYtOvdZ
UpMMRMnfcJhAxmCBB44UQQ8FfTo39PCPfQ+O1Q4ztrUlOymPtqrV6kDXbg0llNGp
JtsNOYYWH/Wut+lWE4adAdbUIjipgRUWEuPHp7izHq/kOM8d16gjUKAUeXKYVtgS
wLqCZlOSTH/+6LC97nJGCzyP45q6EY68rYlaYAmPPybJwyn5R8yHgVpHRtKVb4ue
0TU/C3Qw4o65QdAJMGqVloW0kNBMQTdGu33LyhEnOD89q2cnagwtZ2xo2mtENxF3
c0YAtmX96Awl7infCNmBYLm7WV74ZRCmVr4vlkeeQYAt/K8BmPQmI3DAyLw04Ml3
rgrblTieqPYxAYkKy8sgV7GNXMTyJadgLa7wsiLb+T/NeuoPfpnfLfC1zDNaA8Bo
fjw1fq+YcdHKbluIGzrvjCQaF24A4oXMAUCl7B96n3SQ/U4bRPRX6tksn4Gf+eX8
Xh7KFkHrHOSjRjcUAZxJcdfubCnFozpOuQSsXjzFbDNzt8qVz2Lobhn8/yfN5FJ/
H93s97HPEZio99x9CaeHzMlU5AaHCbS1dGGQFbQa8dpqRZqzMtImxTO3c7ix4w3q
ECzwWcFQ6V4xEf5CrXYPW7Yfj4AajmYhvtWBb1vmexeXjq0OCVlQ2KxuuPvLvMj1
Uut4hR1bNaZ+2/+mv8hxSk6zdvp/MUZV8HfhJF2jbbrIWQdHoEE5i3fy5fZJer5f
r85T2wwBLn/Tn2dt1T21seC2CphCjsnsr4KjpMuNzwZCMcISIl7rLtf22bEJ/rhx
Drol7D/dRAtNyk5Jp33qyO3U93VO2MXhBPwTDGKRJMDcw7kgCySERLNxOMi8PAPy
wLU0Hk49kuxatGZK2WZCiNxPAFfttQ30wuK/2f8L7biXM/yhTCwTRhI+r57ujH8Q
Ix5bSQ8FWDnnyv5ycWDHWrUbDy1gW+K1j+w7GtqO50bT5mvMtrCS7VLcTF4HexxC
3NHVhZm9/sEhk0ZrKb8OuWaI3+gqSIyRzWZOBdjQboZGDv0XSnfSyZpNEEq5vxL5
tdSPs5AL+E6gNsxVEyq5H+P9qBT4D5FRzn8rQFDOaHE3iuGIbERQIVYAqlF8lQ2v
JVQY1XON764pbsCm19AGVO2fiY4mqp9Tg05h/ANSw0Cs97MoTSHg3uwrSCsz/7wB
RXqEJw3d7J1DBcRs+oV2IzfnAMU9BKA9Xqba6k7oHv9y8lBvUR0uuOeEey7ThyO+
0iXg4y1lWdmNpA7iP0k5DAOHc0AXU/kk+SjOMRQqjHAjpaFz19jSPwCBXWz6lE9T
dxXoalpdqzxdxKMYYgHDruzNDWP4tFpQcYuHIOogrTfQ2dOxSRSG1vO3nGjDFkJs
kIXw1zJUa+y3bq3UmE8BNrwE+aPupNu1VH2P+1Yi1SQVT5de99HhfCij8afyHJs3
l5p1OtzDAwsJSXBVTdJjpd6ShXrYaTfqshtk5i00bgRjmdeEfriTMMEuGROPmGx7
OWuCBLNQ1nfVo6uLkHFs/aZ7e3M24xqbAjcOvFCH4ugzdMQYI6QYjv6qILQDVacr
qOAlprnxKQC1VPSGJSbtPtQA7G5KvMtcpBcbd3uzSkdxMg+NqRlCfuH/o9q4dMVp
ivKD22tfYLk89KtULqWZsUjoQALeliI+fI4JSMKqdVZ2p6NwUzFw2aEYeCJ6Cv5R
d1rcgtVhLZ4Vs3Fp4q1R9WtqQ68drCq+CZfD0kbXmVmh9SZxEjDqBaUKnbBJRmhp
eXJGds5lCcRLYz+5FaZM7Bzjp5JTH0+mykV5v8ehVE5vNFLDXtU4oZ/AVLl+T6ix
dp2jocbds9A90lmPpBq2CoxtPTH34oylizwwq8m8sAtvJ/EsGKsjP7k72bc4yUi9
peA8lygAUKsHtlsGWq1pvOzmf7E0QL99aAwXU+pEab5CAE90+RFCNMSegYirL3ZF
UhnTmOpvFXOHBw7D04fK7mNELMDeDDonLAyEnq9owta4q3XwJTje58g7gtI3OTVY
ehAK3eetPDwIu4i3Y3+kIz+IDS3eUxzAAWqPaaZ2ZMKHaG4yVH20WgXy9s8bcsv3
CW9CZsRc8lj5o5GqvG1lBFu4GuE7SyxKOkURSoptZsnqPKuTXiL31WF0rW0V8gwj
5ciEkDYYH3SRnDWNEhzcZxN1A5k8OzEYr8sN7anxyT+L4VtZds+OJSEPlPtYzt3h
+PctFzoUnhYTYBjwABh0TYQ9zZfshms9xugGBduUjVAfy9W25vXkH8xzQpdBOUmX
+Jy6CvL8QqBTAZyK7hkfavV6OlltP+/e9cK3mp+ZqAFksXX1E9URQyUXzUUZyPl+
yPtU2wlE08107in9iCLpn2IhBNiQzScV0qw7MP2TaJPHuXxNBhPtpglC5k77cHuC
BFiGULiTI5h0Pdyg+uIW1EwE88qb/ywISMzaDIDscbYYHqYOUV1IeAzFSoPST7UO
JJhTDweAOhZm0NPo/fPMpqnF6hQkDltP0BivcoHDx/hYx0EBcP7InuV8MwXQF2Ox
6MhD3qlFNZUq6xVfZz+/PsUzv1I/DeyxHxRIJOT3zpDOZf+T22eF/1oHuCtaMF4q
UptgDfhhzPbrWbp9tKn8nD/xupP9DhdurzrK08jbtfS4TKNWTnrGNtshryLmKuDd
2MB9AQnkAAI1jg2JmPRqHUk5yI7i2mtAO41ATIjatfRry7kyW7hb6NlXhbwM5/mu
iKmnobz0b4BHPstxABkeXuEmqMK3F7cfUTclx8lF8SCZIwENhBQF+UPjDy8GYPss
nFibcJlfXjOeGfDuIGrJNrUkJUG13uFko+rforJTMQ7Rus3d+7LcbHYT7nZR0V2o
/pXXW+lE+SNB1AHshwZqHp76jSIuW8f6hzEUOADHvqFw/Gq58A5SjjQtk2SDy6zv
BzPZfs0BQJClJdixH4uPiYgfKHUSuwf2IMaHpGyxTYoOHaH5hpeyGNVp8vMhCYHb
DP0kFBgT+CjvNULXkiwEBJ0GWkyiTtUMrojL2mbvAG80JeZrMdo5WuCNqtFtN7Eq
Im6B2yMAO/fwjYmh1rtGcS+6KVn2GaGcrtr/mU5xvwAgMXK38r3Xv78P5L2xapnj
hyzbe/OkVsfvDywOxr1Cv22PEQJovAvsdh9i3TZBNOuJekG85W1QtmBQwx2C8++V
4ZrY9FqXQ8xVkDTs89R/q1DwtQC9tW+7hhNrh7vkoLQIJ5mlt6Xfvt5CwJmXtZwP
1jDeoLth5efsMDfg7hgxh0w7gQ28RpKWq6T8kY5gRGCBb2Q5I/0w9wzaU6YyXAGU
hPWmIyItP4bfGoim7wr72e323Zcs/tH0zIeORcyNsV/8WmaoN96YFvRRgyilhb2s
pF23r8fraCRXYjuVm9SN0MOmcfYIGe59HAfBPZ+dAOcCRe8qBkoH97oFtH6hpR/4
DJ+ONVhHoqQkWTdnQ0wupO0VZ1S72+YmJFN+NyWMT8w1koS/Su8NhxS+7zFFnArv
R1co+RhYnW+xeKUVy6qstuuFx9sEeEM/45hTQ1pHGFaSBIVP6+zsUL5Vepq3qscs
KRJUZFI47VdzpIz5NLB5tvSgEDCbeTba02UjMHmbvUd+R384cxgPGzYPC3f1g2Rs
OH2CrK4f3jK+jyJ8M6DcUzszIM/L689Azq6MBTavnpQH4Zgu2AuDmN+UTivqrMQn
yIk72YYYuhS5IoH4Xfn+0UvALhdiAIsXKJGYkIkKNh0GGdZVhRv9cc3LcOiGDt2c
5bs38ErHaxmGQpvf6G/mduR5ygNBLZ3KoidAgqrmcdUs2VAaHuIwmeMMZ4aYQC3j
T3IsEUt8kDLjvzsPOp9eIPO+2fn6TcqFSLrj/wIvj4JH8ufEx29aqQAfjL5MBbEQ
6i5RCq2lSxHGJXporPmG32DtUwxnyB9ZCGje24XcwSMKyIntDtW9W4yRl4XDSPA/
bD+xmJLGPvsEeUyw82sjlPDkSqventErfhqH9OmhNVg+xQYdOFl9cg1U8noEdY/U
c1PHBbw8zKYFJ1xt1AKR0z1DN5qXQApOxzKEt0VOg1nPnZ/03VXQQPpn10ORDnvE
WRs+raFbesVyOCjPOCcSjAVuQou4If+ddLdxOujbt7nJcA14v3nsAz1Z8tmVR2os
1+4/EdS9y9iNu4x2rPpSI7MZ/pAkchmnuFjzKI/bPHo6yL6cnoM0fnl4lzqFW5PQ
2JhilN1bGRNDvJE3/wf2J/7hQBBYoC+i5fqBqt1Dv+x7aqy4TTkKuh7rdGKFg0xl
OsK6PyFRm7r7L1D6+X5blZbn75v7BUyc932uony+zvjGw1pmmEtmju/XQlWaK6Lm
ogGIiDvGseOsW49VMLtraybosf9/0ebcUK+qYyFTVHB1gotC7sBCxu3b2FcM7piY
xOu0+VmF85turZxsgv9PIIexjFf3Sx4uGEkMjP8Btbcm7DmMvz5Im2x8bgsUxtJN
zy2QN8yBwKZ3X8j6mA9zCRuNIDpEGJePKF1yMOD3KfrhxShTlZgQSaxQUjCpm04f
cbcxnFJyuMlEZa40jvYJ52mLlYgSVKCIHNrGYBd8F+vvilS2NLytpX9Htre24Wa7
Hd0ZosNhVYgy1wQak0YXfIgLvUcIDkBsmfnf5oQAp3o5jAjD8W0GfXBiaYnvtBkU
CJNG/T/Y63FRThHgR3eloMJbHIamGCzW6/7UBa5HVUA8TG+ca4Nv8T/qT6dNCNC6
VcWi+Phf4WhkfiXAq5rQcsRK6F43Ar8x7V4X8hCxPjTOwNahItkEbV1UkO+2/YeK
Lh0Z3uj0Cc7LZEw7bnPi1mFJaeTc+GtKmkriYCyQ7JqJscJg8Unv86MLZrSJUM66
5HGxoEUPCNwd/OfVnwTEF7uXQ+CvIe7/zGjq8oQZuvPrdTGGuzKxDjtN9YFQEMQ+
xYAOOUTB+x2N3cSHwdPDXnguujWMeqZpeyUdOj45t/f7GDymSqq71KVp/h7+p4o2
zlopGlJrc/OsQXO0klmPx+f9qLhR3MEWYv65zXuhGTSCMOkL5RcIp5yvxoGT5AYp
7zS6rYti6hHQidZzCBmGNDHWtgR8pf6RETCZ6bQ2VPF/Cz0mKMnS2DQhlE6wGJwC
9ya5O5jmbN7RfYA34Vs19JLGINvkAkaX+cM8fcrY28NU2O8I4GX/G9t5YSawAsHK
tL5GGnsN0PZxvHXCJE+Z2gkSjwrfgTXWKHfmm1P+ceUWWRN4Flhp49r3cF1a6a93
XO32Y2WMGPy8z8jNksEUFxJQVbhScvz8I9ikKQ3oGH1nkiGCLdyAMrMdlBbdha8r
0cKxL6YTEhgYobHpOeFuEazqtfSn7gmC3oG/8aQm669ZnXF+oatCuOwRUc7nabRg
/POmUJyuphiRu6g7NrRFRSiI314QZO8J6gNkDS9mLbHVMCEKXT+qFyMdr0xdQil0
oHXw5C/xWQ7/4+VI5o4K3OwZXPS++9KlI/194pELGFS84IGogHnXqzJyMVg5RxNL
maf8U9uNPrWLeyEl9nncMBHhxYL3v3ymQyU7MYUhRwOYGz1WUvniJXjWnt2U1JUp
LW5c69xjX2VbhGm66n/CP2d9tN/UulPbPZ4UGSeMqhhTBi0SppBc86J3MBc2AxKn
K3hvFQNBxUUA9KoGdO8VZBAUqZGDhl9ywIz2DwT+5mFPa12Tt/zucV/vL5TG+n4d
f9lG0Yn7UJkTK/MmWP+arz4PqnbS3VOya0G8ERxgwkI6hMKNZM8FzEtCdKZGBTA9
mx/ofC7YdPwzOi5B/PQvHi1f4TUxCpD9+Hz4MU2cMrJkstrNvFyiS6fAptXp1M1R
HYsB01fYZbAhH8MOBIHZdInRzM4LRH5WS6Lwt09zkuc7X4Ks7UOU+PqeBSE4wLqs
DrQmSbxJeFb+TbMhgmwIf5B/kuIuaKOkAsII4x1xJvOTa89toFI93Fgwcc51u1R/
EgK63Bp4zEALHd1nBW0z4yOOvSGdoSZg9eGiIansvVOMF/WocltMmZ9xCachuruU
sMCTSuy2yXfLdRfHrRBuWdqNHQe1tanF2kCmuuDfAjPTEBYc26NB9gpkz3GDs7JB
6bNN6Bf3TMEVwH8Kw9QofMG2Low9smBsS6w/+mgJsvdIHpePHtaHxqWT8oEw54cp
i2Dta1cJzR1sBERcE0gFsTpDBOMXsMOs9tUgRKLFYOrw6mV4zq+piYdBUs6SjjVp
gZmtSgpeXUzSqetH5OCFxO5N/zWVSuyVIgdXxyJaoncoQmaNObqtguwN4jt+sffE
4P4K1WwFCs8F5xffzjE7NaYRFXwViutuKedX98/cqWca2PplF9q6MObk7wC8yOEU
IxHnsgMLaErp7tcTf4s//dMsFcIs+b1fLVeImBdi0VuKF2Um1FTO1iAiWqT+cvJc
qREg+O22gT5iDrkv/V6sXrXa6vHLFxPw612cZa9/YnZ2SJsXZ9Ukxv1bupt61ftk
ygRntXZrXuotP3HwaOXhT00uMXqvBJ3a/leIqRBx1G28GmIWK5y0JJAVadEufMaG
4T/33faJBPQjI4ZtpCXVR3ss+SGBnPrHHy3ni5gclnPAeHSSuOE5lrG582ktycZr
6isCqRajcT7LsaUIib9hPyB7uCw9gpgvNASfRZxRmIx4raVe75tntf+lp5X0jnF3
t5f6NrZD/+OOxVYgCKFrI0FxzFYB7oX62SDQrWV43r0uv0GUeydw1s3eG72FXolz
GeIXGDKUp7DeErQ4Xrrcd+T9fb5RgT8to/vn+3Py6deGR/tt1zXl6VJO40Ok+pcR
HUk2jBKL5V0E32Y1Syh9EBHAVf9I1I+0X3RdX/R21BcAGkyR9mKimYYV7Pz1agK+
e5S/k73T6Im5e0Vc9tRZxOvXrtms3QGKbmNa4r8pfj3X5+JB2byceLxjz0K0RlZp
RWQwf79p3Dd0BfKBAZ6qtzVPYFG9gmMTLrc6havYpmexfOtcyjqvv419CauApt7i
EAwV215YOHWIxOq9W1xz5JV7dc9kdo6xPXC2FYXSs5+n8QMYiiHaviT11tgZR/Bn
ej2fFAQ/26cJD+H5JawuEJBxB5ZHeKfrlGss5af+Y1+7K0MM8beLPaqSgsvtfIXP
7O8MXiNyrL6Fqz37xc3mXGWXS/ygOYNyH/PDaSkZfdd6i5i7wYKNg3puDA1vRTxn
dWft8UiHIo8TP9RGA2irdfyMc30AWtkGmZzDAM99KE931D9sIBGGyzxN/CE0mIl+
EoCXkB2jALkrLObFMT/5ssnGLNGZLcC+6nHb9Ww9Nwaub2ndUg85QVbcbs7zlPrx
E1vlaauILKsfiUQ1Fo4bYIfqKnCFPfl61hdR+daGVY39nIDRWbnEtE0hmIh5GxMX
qGpkTb2qlhC9eA5JFq6IijP8WAdI2KpPrWAiV8lKddWmxnsoJldglT39Wy+uZ4mM
C72gBYeUWn6KKk9JH5KMsUJGBrBMrwzMT0jul2NT5hwrkeQyGdN1uPofVpEskkkn
SWf9E5HGNRO56XYKrdmhTMOptvD6gqfdJcWGQ4AbBBiYZvebsSpUyDsek9CAos6r
zMSE1tkD6ebU1QjdeET42DF4rTDaS/egH5letxTAiTZK1YrM7GoG6s+uxpRojpSe
d84x7N8OWUx/XZZ9jlhHRadTs0WbmyhkWH7ldCl82bBJBjJhTYFfJIEZ9Oak5kce
oT/JcJQMPDAntmbHK+Vo9X7d8HJ+JB1jhS0leq/Ptk6WXILQ4FGIHXuLTk+tf0Ot
PPGhMK2TQk8McFG0SL85jVDqrDJHBrP3WDpOKd1eVIiwENuhL7RXSZoM8T0nTjoz
A3NuMA2G5JhVFGnqUGK/BrjRpcbazJKnaZF9go/XMu6HQvqR1TFLlIRrKfqfUiPa
PDStpKGGSekgTspOFx5v6GEtHMeomWtGoegVwxI2e1ezK9fC2eDIiAxUZRjILTOj
SM7P7aQ0V0nK2z7pytlnwyd1eQ4nDX5uYLezToF07adXCq8zlS10z1QM1mSEKZcM
XG9TlozmCSMLkKkeWaplbqlxX8E4u/FSMsgogBTo81Wt3/iYM7K8F7oW3AjGy/h2
vugUibHSwIqlW1xs/66FZFE/Ge2d4pKhYR/G9F/SIZfXBhy7/bbQ9OlH4RnJiJAV
cz7YeX5+uKO/yxHYpEhX5o6UiPaZEUNoRnBW1bdPjRjThWgNCl6AsQqB50pVvbYx
vcAUwlujFzzx84QgtrkOueVaeheaTQD4kDAdcIlZh51G53MvTBJctHyYiMNPS8kT
LM0alphaUPUqMhiivah0iXPp6653Y17CxLT/ZvROIsbTm9oagIU+natV1fgw9nZF
qMqsLdYOC1RV4lvdlXJujPgFz2beXpXUXlL2KyXXou9w/EW2T6SM9jDzejqti6qV
UE4kymnigc85g0wQnrgP0JSidnfgS05/ecLei3+AuBEuLJgLHliU8s7TQ2KiJrgi
p0Edwp152VoV79lP2v8Kmmlq0byPkNIifFAFAogiuTNWCW/DsCAazai9XvuIGmYD
eKkxLlhvCmZNUk+HXzZdbFvhgGVmT1gC2N2AQPYJy+Tsbc6gJMvUsFMehc5zqQH5
slxrDNhuLIH06BoOOYY4ZZkoiSt2cCFe5+Ea/ylry0VMORWFamREdc2INH9KCJt4
HZcHffoBWpURvs1ctLchrb+aScU0EgmpMqLQe22nJJrtl0GGVjc6ivY6YxZvX/YJ
dzxVkBgm5b0Cz9gyKKsZ1a7PlUhPrHVxpDjp/16v8JdJ5g0x9zdlaJmmMREVy8jY
pmwGgnquBMGrU6BlnYZoTfKDz7UkLVXylB2EmOd/jmzIOT1sqRmQLY2Bdms5i+AL
gBhk3o7cSsK/jiSlgv8IADQiDhtUb93Onbcqs2obcWiCNzMrcxHUcfmKPgrJD24Q
jlaKvuMrEoIGGZHJiYvg4xgqZHcX+YmDqbB0YaU3OW1RNoEyf6Nel4Gg21m4X8bf
/Ri/a1sZZDlEmZWgY+2Bm3h8uVjvQvycnkItteRgE7bj7Db3otE518rbrdauJX9P
nvuesnpOZQC6V1lZaPyMAzsmFyLB19SBdtjtjYyI2UCiNum8rLt6tRoKfCHJqbpo
D9agCdgQQmHsWe+Ia6oqCF9RHu5bEkEHIYwQAHKMHQnBRb2xs+oPDnv7Le5bxtOC
jLanI8uDV8AyXsJDUdewl25xD34fMd9kllp6g1iBSq+TWHjPRJg52omCsxjf8s+S
AYFUvZwMXAttW9O6zVcmk2GlrtUB3ZFEe4Rd0der073bV2DF2mxlehjY/YFfjEVY
V71uwadjUV9+5dMMrFkCnVKmrBiL9FkD5Uqr9FB1dOxfjXwkh+u2yE6h09yuvVW5
TYcP0j98iMSPqt2KlE4mcgq7yfYeXJa/M6s+dld4jWLN8EXu8b23/onzYp7nLyN+
AqltrmXsJ3y8AAZYq7AMP75loM3DCYJblrSczsxDB4JMzuZiwIj7p1SnvnE7Av9w
TiiZVyNrQQtep4HOovGrlCftB6y2GPPwXjvh6aG3c56+P6NfMZ9Rys7MglJRMS3x
C6w8sIhqJ6Sdu+CMeNqWgwLtA3/2FE4/p1nQzLCZL4cQyh2hMuQAiUzRbMYJU8U2
kGxIcZS35GbmfTYxDL/DwZmRhx8HKLYkzoGvLgbpl8SjhPYUj0LhGRdP0qt1AZM3
Jx4uiOG3HK4u1KvXsDF64Aw+VQQGzKtifBhJ/OcDYffrvUDw0AuRpQ65ZjlIE7Op
OzJumJuMwY0NjiCevh9vUJNRIUy/+Ax/i+n5YC2SpJXEAi8/0hVg45nkVuzQJgtv
Je6VFByRKcUUVmar5sj1dI5iWt3LObP3/eMdtR1MFZwxLav6Qy2XaeRdpeDvC5Nd
c+bVVosZmU581xymp5PAZ4PpAh84Wyhh7v0LOTnI64IeozJKWWwoyrhR9ruo1eeN
uxAmYywjHjrH7IQhlQlTMrBMwYIpQvM5w2qKgDaEsN5g2slgN5epZ0g9xGoZnZSP
xZo6EhFhc63vEMW6NvLa7ElZUW5Y8Oe5DlcFz2yqkR2hPcIYeOAHd8PjcrFrvXzN
FL+PQLOIPpVjjC+ouUJLw/O2niGAP9NyWaqJq9CbWa6nbKfyLh2rJIseR/ZEs6Z6
1BBZo7U5lXC1GH1kLa8KAUbkbRH2ps5dz+tVo6lg4gYp+jZrV0wbWSM2HgqMAfSR
R/uCeRx5S7VH/frJTSIbyWTQ/y9GPnZb3mDYjTWKVlXNi4feiMGPaRIbRYDapMRA
mZeKX9o+FX0I/aNZK2JPNZ0CI0ta97e0LyIxyO5TR0xCJS1/rVz2JDjcAExTERNV
vluONQDyyAbMymAyCG+s9FBObszcyvjXv0sqxnoV5vGytNYLttb19AejSyX+AEdS
1N5Zvnwc2AoX4U2M9t7IipmONB+HLHZMqhtHHydyqMUy9E8yCaqGhh6HyUdyu9rE
J9bEM0PygvHKr/D4adP8zQyKeQM3dB9mWZxwv4Jij90QLVoTmx+lDue0jPciNCjX
xgimjWuoa0uGijgcIQleRICk9ZDM669SO9M9qNrJAgASxw0GEoo3rUigwu5zuDND
obgk+DrIZfiIsLeEt+XKorzJH0cjObB5ZJ2i8T9S+6ospq5S526i4DS2zl7BnRMY
dVMtf9kYlekatPeq8jAHL7sd5hbwlGQoYVn6JmWA93aaH7GrwvsCNbHS66144hQp
wTVvpxYg3p6nWN0Q3RQadqzbR37KwOC1kx6HKNbKq0l67IwslNknghVBLttyfhwZ
86A+WaIAhmpsICTuw4psFYbEr1Mh11VnR03PFbyCr0UqTHzkGKyQX9uJ7CZ5DNKT
ERRVXJ56lwwib7a0pN9Mt1MG/s9uDrQ78kUGoohT76hxs9r1rcZ2MnCg6VMNrJ7X
0xVETnORl2EkMeBzpmxC7lp9ff8GH+Wvirx3yVlxbAilGacCvQryiCpTAE8YIjgl
RNRzmPuRaJ9cQoEFxqQU6iQVR7oFciNE3atapr5jmIW6F6sayTxaJU7H7D6Oss8Q
kcRObdwOmWvqgMgpMTIjDsUod3k70yEGIy4NZvGgRxrw3tu/m/PFZGYxNMxOD5a7
sksDc1dzf4a2GjjXKzYDh/wdGo1wqHBUYBNA+6Ds2Or9PraCTA+Bc77MGJ1TLNTj
KFlfca3zoFXjrZmXRMkSYZVbexaukBu49jTaAnOMYWAEfCyrXsidjsjbXSziQ6Rs
StYsdpIT+JEIyaUaOgZj+3vvnG5R/mUOP33lWyVPo68RoR0R6+pYdXslSO2FyAwk
az/pFd/t7oIdhBhysJHmY9xDSF9v0ifYbmagMaXqAT05yr7TwqButPR1fCC8kqwL
B4GM4iACtgl/hih3MZzLlqwBcmcvFDLNjiOA+Hierdm8U+WHjBQuRXrpJMaRsrWL
1gr8xGt+tmQKz3end3K2vd8JzmQboXIbWc+Pd4sLQ3C3MDnrB8p6rKU9C3btYl2X
ti/OoOqpAvKy6jvETRJOTdkxNbvqwDiK9c2ooo/DuuP+0/JMT8vB5/UeAZupopHg
SyAlnuJ/vxsRx3Gjv0JA57wUMTP53OiUR48NGDuLSLF3wlT9RyEccSazgKFB3LlX
FsTxGEdpJCDcu4Z3LZ2saweqH09fKlffcKFioR6K9VX6PRzIISopifcF+bnnMJs9
NH6VeHQcsFM53HbmC8njtdnll58ZvYyB25nBS3QM9s1zGMwO2g0oM+CJk+P43QzX
BilIZAJcRaDJxh1H0KKmaoSSKu5Cnt7nfFB6M3iPI/P4a10Jb4H6PmKGB41gN3pD
5PvlqR96O2ZT4Msrxsvk75WGBP1pxoSK9fWHVXx8EsejIJNDUJCIU9429J8UiRCw
JnRc+FqqO2zIAtg8M2zafg6YX+LJjyKDbU9n5OzLxI18VWSKiKg9dHryBQDEUqOI
2n6T4pbV+Q2fIG0vkOyX4h6Fj8ozWkbyson66plSImOmvxWO/Br3yYatOMrn8Os4
h42lXU6EgsBVLNNYyY4/ScfiH1dtdkH2mjnWfDLCke8i4c1iKi/dTcKG9ziZRpQu
5BByPJao96TxWn8bSp31CuZQaOFZqenofkyr8VPGlrl7Pela5NpfZI/53V83+nIg
8DH9hPrH/ch7TNv5/7s/gVtxYV+q1chuYz5nSc/j1OgHCrymakXblvWW2YNU+R0F
RNeMvU3+D1VLxsA5yplPlSp2oz6SfntBrLXE5NC+ZY27JG4ZeBwlIKXg+0EraWQh
vSqxO9JMulL4LS95feQtPMKwz8t3yAA5MKU46CQ/O5nf/hcGVZZ9YrCZDi4p78/N
lgY2StEZknN5BD2dXfHFWkWz4ItybSse4b2kDyrY+dhBvu3gbI1XToAUXIh+m8t5
NjgzKw2bXL2pibTruQl+SyiFD34wS9/J8O24v0rVjHG26ht6kv2+peJZVWk3fBh4
UHZFa1HE57n1S81b+p+gVUMAAccxBgpcwzBhSoRR3FL64Y8M+4xD01OTw8la5IyT
pIHr9Qo6pPBE9SmnP5qVjun0Zxw1BHBu+jSSf3wNZPjj4d+bhbWSDAxpFKAVJFG2
LiKCb/K9bboZpZnyr3KIKDdmv9mFUcCC64cYLKyTiJfJh7q/3jxe7SIWNHtxmyFK
ekOqUKxdmWMBv6XEnupoaLlTqmrYCW4noL1qCKiDFfHnO+QFHjcOpfph6mspWOxZ
j9u57sfa8wOr3y8Wc3gVPZWJAp4FOxYq6y8+kRqrkMAQkKc1Q7RkY0hyjvEpGFZo
Btx82ls0nCaZP+bqwBryFdksBXCMsoVLcEzkvNgUXiJqDXWQGSb2CaZI2V0RizCx
sXZeq8TGwA+5lqVjxSEda+Ce5Rue0fodp7XwRMZQH3sQ2/GE5VwMHYC9lBZwc303
3CBnRfpJGTVBBUI1yTBHciE0NjXX6F+C7LCe+M7MUnJtzTTZOi7Ws5uv7PPQso81
ict78E1fce/snYI0Pezi0mf4vUkBrLdXUjJYlYQMUBFS8EebHHLWy6BhGWrTdYwe
1vWNG32EWVNMBuS0QwbreWdac93SBrwn+VawRUhFkWzaTrbT1GuBBG7m24qL39G0
5siHlrQjze9F7oiB/OoF6kjeiM9yfSw8vlTuclEeayTq0/227hLAmqIRdYbYDrKH
ZI/svveeAHX8dhJOARYuGPCeR3blymVN6EjXJi/PLV9nsF8t26GJ1RZ3lOxIlYSv
h5yeAu6qdmYdEDkHPUZquWuAdp7rETv64jSNk6TxDsbNs9kWIj0mkdcPP96BBaKr
b8mst+ELdAeWa6McT4nLSYLHXYEAtfu9Zx100haWI7iMbaFW5D4OAdT3+h0utKoN
Xl8ZHrdrR0FYb6Ytrx/2LDltcCY31f34HzenF38uRdBJ9Jp4l/8KNoyKRrNEsHve
5OiQRBC/MrhhCwF1f3VmdyYaEDcMsFd/9R9IjuWdDRoyfE8yb+n8ZFVaB/mNefcx
AvnE5nV0zgwLB0txLImXphxrkqFpKWNC3y66BtQMuDLnpDb156BG8WHm/qTOROOX
d2NrHYuhH1OCJeq41C6luVnN8561TReKk6xgi1KsTBXSu9Lpa7CXuCydqHLjrNu+
3Lv45JF9w87w6bnCBQPVQtGzt2KkcDSrO6/Eqh+JoN14u88D8F68G/LmCTyIT6Yz
udS1z8EjilvMJIm3/0Ol+v1Uf629qQ9V6tKjqRRZuULisHvwi+JaGPj4obVRJpnq
W2jYPOfZgcxrrV9f9m9vy2wd1GgppZBzRc2kv9uPjmaunjtZHAs24q6B8PM651Fu
6qxoXxmK5myslUtzWZF4qDcyPT84Qr9ekXfWcNso7lhC1+yp5EUfZYZL2pPGDL3P
ztZ413g07m8nxuu8olOMaDpMD3+giw5uM5s7bOUoPD1kLDeAHDOZOTnuw9PRHuwN
Hnqzz//AWa5Go5c65skOPFtYFTVYvti1r0be325BSSnO5nmTp/ZnRCRAmgIrQkE+
bxsc+QN3dnnXorJadAp3k/HdIYvfeSjG30MD5QypevK6Lt3ACWZqG1CX0VgbsN0y
TtDcMmn7g5zaVXtzXPFTU5+NiFXGAQmfX8ua4QN+Dx3jIUOB7tBsWkALNA2+RFHm
hMvmfUs2yAEqltrsy6X013dWCVDkweARReBn8NM4IVVRQDgS1EY/no71ntTjEq5W
YQUaphgBuTAEa6m3TG3+C+s2fO7UeSMifc38u4y8r/zrOUHJM9SaBsW3ZfoUBCDZ
rR4M2BbZTOOttCYxJ8bfW7b9hF+imo3NB6IqTfR4WEczkBo81ZX5kSseGUg2hEp3
f4gf88/gGy47JWtN1fXpTscnLgPgDHV6OAzBe11xKYx/qnmcb1G2pkN1kcKr/Mmd
Q4CNkW6UwuzE59S/XaaFwLpbZQ/U2gpNzUnfiil5tSRz//vMzr/+Yy0FoAMuQL81
DiKDrDIIzYMARUJQXf4CrAAf/FanJHIcf62ZfmYl9+6jhq3CyuWw7s9ia1pWU+MB
9ArttT2YF7J5TQTdQAms+X2k+AE9a6feaXy76/vycxS+HpFk8xC61IKTtzpLaodj
6g2Lbpnik6mfnPyrBRGt/k425B3susraXQ0uUfGNpODsdHyHyQUvNiOM/wuKvt8R
VjS28D0Bhbk8l/LHMw9xptaNv0kW9FnJ6fccAIBCZZ83ZG00ck95KWTF4Q+a3RqA
bN5SlUVsEzPgXG+M7Q73xGVSUoZ13yzltnWblGsBxdmLzq1KbCC4rdL6RKDOHW9W
iBKay9QcieGqTBpHmvH+7cE17VRhVz4hqX5CpMrBYZJbxJeMbv+x7WAfgeShdVdS
kQdSAuXesbrrljNORGdULnmR0Dk/szN9BnVGQGJqxpbIZjHM3FPUkj6j92CP6Fdv
eLFRunPQi4VPbayPXtplZMhmb8D+BRJ6LOZOVBuy5pNz7tLBIu0yTTrdqnqksI/b
BseropinOXK3EtuxLhuNwD7JIMXe6CRwH8N7UqWq7aurzjWpCSQ8BNIH5zZvqaj/
owGPhWWlr8LnbneWXB4bO4rNFU8Vm2xheIlaH5xtNFSlDMAIcJwNqdAMsvOWI5e8
DwZOacr7MKBtjF9nUUoRhoPGSGeEhdPmgoW2XOjPyB9xS8RWYoAtOtLkw7eC4RKQ
lHJ1TxipV45WAafzuiEDjabHusczxgK7+XrFNg1slckgJOsrT/LbkzuJSrmGIFIw
8pHmQZvR7Wj8gfZB0yTUulGrn7YkfN26laMZRIPxK0GmZB9CwPrAxlDs0AuC7CEa
BxN6yZqggw+nvT5gm+fL1A24DnuGwKJ4nxSYqUvT0txs3jepxuWk8LN0+To2Yc4m
Q8w/gGiY5Ugu9HN8NwnScvpz+EZ7XcBF9epX6V4O8tMvwl4H91LsoJGfYdozKl+D
UY0SXChCJJcO1L7r5krTQBdrTFVF1QYfeYmYSeExaYCoWnzn9hnjDhkwARfUpEBN
GpUH5VBdPflJmu0+Dcq3AWRyf3nKlje/9jVQJmw99KGsU8YWj0ckqknQpnE/bGvJ
YFNUnw2plQHOYqmc64ejFK4h3oNWGzKXbXg5JBAhKu6Tol5gV9Z0eG82I9X2ATj8
govXzgLTEHmXe37HWmh96G8BbrwsySDCJ100r6e5Yz/CGWW1Ay3I35SgYu+69vv0
N+fCxH6j56RGcsRUuZ5zgM8a6yIneDj//3MPIPAXY1UddbByby8yAKHjV56+8N7B
ImnmFw87YtjeooHOge095ykTjfD1GL13Y+ZY2V9MGtrGwVQqUOTCg6Dhc63ZkPL4
APEPnXOSv4fHjLNFfxoNJwsRkLY/Csz/6kH0eju8Pt2pw/kHxXpLAMfLLtoKZBDI
uKD5VsvVdxpttYNwjERb+DDSQabrhCJEOaMItaSRICBzTiFoM1SPORYsmzmFziiQ
hxrsK2VFJ1Jyk65m9krS1fzv0ej+hjhx8x4tPAvuCCv4BPtTCeRRcGIJAKJTFQhS
f0I1yeLN0DfFv4FeDK4lvPERlRVGLsBZuiGFPAnLsSoGYrLZJXG73FvHMjkJX+1u
8lPBkicdelGK5RSYcWe6lGHNdTwhR98r0ftGYaasrWtg+ZUw5tZ0bZtqdA15dlFh
lyHPl08xERs36D2QOTzNkSHiSrXpaPHpQlOeUP7M9tV3/0aQ22n9cjH1ft1G1b9y
NiV0UxF8m9rbkZA7zhRzPemJ4pBD/dJrCc9Gbogm+n9fYaOuYvi4Np9UET8++oM7
ZTQS5x6oDnIQGlaTXYgsf7dGf7E6/3doKo7dR4iNwxmeEgh/6Z3RxXpVMUig+ZhV
G/Dp7ISJBkua8NDSPnGHtE+TVlM3uQkdnTSrTn3rc3S1f0eq42lmFD0G5ThETDMm
7vuMDHzdlZh9u+yvqmzuIP8po0yhffqiJhOVfrBF+teQbxsfqwW5NI5cmntjdxLH
jjM1zsHSMZzbg4QsRneliK3Ux90E0vBOPoxNIrsb0KWckOZKg/02gHCAV0+rXWaZ
4F1ViSAONW1LeRd0x8jnwg0x63pQWSMuBHGjVsHLFEQNrbx4xHVFGDWPsu9rDSX8
53CpiUz7fnN8lXAXIUVgFaBYtrtOw47pXVURCP15cHrrNRZkW1BhuwQgVtG05I8u
4Iho/RtgHt8oPBNoepje5bMI1zSEPvkdGXmo8mBJK2lmvhMZXo12Op/SJ86kwSqt
vDzxZhOH9hB/LUZLTdQgalR6JNO24n1wznwaYTnScWR53k2YPzSCu1OaJfNcbxne
uERIjfbKPJE4I1ZDe7JOTC5oqlP5BTvTntRFBWx2Sn2yEbEufN/IA4pMZKLNFL8v
fT9+T6HgL/BWMit2x/OCCBCsaTi2Q/UdBrbrxavSUQZpz7abP+yEYrqOa9EUAws7
C531j/nCHR5FhBBOtzL4t+27xYFSN3wv53ApG3u1no7ic4IH810W8uAVFz7ala6W
CMrlv2fi9U6U4bGQ8iY5dmTIzEJ/ssLbhavd2nfzOTbfsjhGceTAJgZ+Q3xvw7er
8Td8a6oPOwqV8Jmj5dXI2EesfVkfdItiyvtCQZquhAghFNah8vS8KY/8mdBAz0/j
AM9hnTUQqo7JPfT03Z2wGPCM8ob5wvVZNv+pPJkUdzX4D7H9nS76gPrLBWSLFe1+
+O92aLL0lWFgvkdj89JofnfEaNu8h5snCxSX6HT9EUAf4Xwosw4hgvzJtNISsYee
2mZBfmtF5EqeWYSRYkBPgCE/aZZrS/EyJKyZ4Nih/MBC5H3gJPcNyH60ftzccwfx
j7ktr+2guUesprO2pCH/cArSxqONNKs5PwBLzXVmj4XELOtT5E+M7K7cmFdu1mas
jcJUxAJ+zImLxqYJve4Ud+H+uSDqaE7YVIIiItZLYnX0/svuDY7arMnxbUj9bIDe
Lc28NFRudBMu/FdYfJMeYdQc1p0LZVTgwrd7Krf2tKxeQD1GuePNv36jptrHWRmH
ukUjJVKeOz8/S9beJnON2dXhlBnLQfJESg0IWuoAcBNDUm7HBFmtQ8OVQY+2Pk2a
7mvVSuISJGKAJpjBttHL1/IdsOYla2SDLR1RLEAXY8dmh7k/hI4wFGU/4lUliAL+
XZyUmNWwn8EYR0GFl5hKLISEp1xWT/asgIWUlmq/ERUxGKdNuebTmHxeyVaXibdD
FYCO0aB5XWC9rkRIne4vP8+gwGcXffU4C0Xy2h9ffDZ0pGHR9g3omvjw/4sWTwBq
sSzdaE26U0t2QpDVrAuTz6GRiWsUsoIizZb738D0VjJMy2RLfwm33mPlW9fRngeG
XFcdYKeoQL2O5AoGJmPKM+LJqvcHJuYHHO96nDhis2cCdNaH7kiUCA3RoWynEjry
ka/p1A8FWxo13TNL4c7xXsss3myVLJWEJAE4XR4eIWI8z3/JezJqUF+FlJCKrQF4
negdRhx7gArUgLv1GPLyUNnXYEWogoy+mtVi9IufJps44QpDzL5sjeynLb9azlMb
3rgmqyjHwttZ8dXVPzZwXVXlaaYvHVn52RDV8bGpfjYkucWx9pmtq87GT7jdiaHW
v0sw+jucsyQwOtyxfFFsflPqj/z6ZCYSzNuHo06Zjkzv/wccfkHh+CtCONofs+AV
56k33yY5QkmTexxTcaQJUHQewCOevDnFt0o6iudCVlBJIzZuJawUPT96LiEyQ0PJ
nDU0YfTRonhgzg9Ccb0/LWp/iqUkyXxi0MZj+cBFPo/O5ChtacV39i08OrrKqq/m
F0x2pX0avggddrgWucubAML4Evwa2XYhoELKrzldM4L91Ig6J7yz73fxm9eaXIjK
S6hDU4+k6MACGxV+bx0MNOa+x7BQ9gJnnBT09+sfaGz8zdngCyznS1NVVYeDjn/Y
hzH9dEyBL+a9s5ulpoV8jgkMbDpLcog8pk2JbiDiYB3Mm0V9yjoBAiVTlR7Mb1TD
cAHEgQOYUCwXunXNYJERyHVfNlQh0CWl+yuJNVPJMMwRbjTpp6RVIIgBTL/sRFwG
dXeMMCDKDI1XtpQqFtY0mf0WjzAObMPhGRNIjr9XufD1k15wFhlRGz8ISp3gemye
eq5ONvCyCgpBpUMeZqs3jaCzUW6wTmMfa+oG8vgmQG/Tp4awBo1PFAn+aMPnSPeP
m+HD7z+f4nRAgSfupJJ5c6GBd6kqzbZJYlipktQoLS86quoJZCTVSocoaaT9l/4X
1VeaNGWsoNzP9E8pCaxnIW/QMspM1m6gs7vAFjAeZO2OCDkDiAACwo4RUfssgFQi
epgVAVDGPsKQ8fK5q/TLJ8GO1bvqISP94CoPxSTtrCcgQtboAs0/XEljsbr1y8Rw
ZNVmgG2IHdYPPusLbBaE945Epg91HOADQGyYnx59tuNXLiSn/e++37paNEOS01uW
HiRZ2FeiBPEBF/7O2HyMCrxCAAR/JEHUQP6DLor+nowSfiUbmWJuB66c72U/zk8x
4C9Vc7sknI0JrTC+sM9rln8rqzCf6Gu8016njxXlKJ083E2jOLC1i1m6jxNeAdtG
NwX+uFiBGOea/fjI2txksqM3wNbLuat8bGQRf6ixZKrgW1W5oX6D8Dj4tPRcEuQr
tphizpVefL9BC5cIez6U3b5Iy/8qEQCE09PKHDIY3+Mo9M+Xe4m6u6YNrkBcdkHP
CvOTwPIBczQhAR9I6fuvZ6OolpabRPui9+BIxoUMLIPwd+liq3h53y2AbAjDS2j3
F4jNEKItOTmJB7J97Kylg7sJ4Vzgot1xQElC/smlv5dkI/2IrUyc5cxhqlT6FPHV
3SYTB7DlxBKbb78ehhBcAqN7RgKJKv4DYIuwFmUtvqi7e+Hw0/5asD5VLFsAftGu
+44Mj3pC/qmOBIurmsn3b4sk0wAmE/8Ty2oDcEXEi/ebDhhpYi+gARiXCrnR7yGq
Y1c/c1hmH1KW3R/ZMyqGjsy5El/aE8u+cGBoD/izfZgxsqkRN1PX0nBHeqHWRxTh
Y5Fdn6wkpV/5apQYTs2WUF/Da2Lu84VScg0d6/6imAgaDfYDlGjSysKtn5M8pQQD
KbZv/ESltUadPDO3pLwr1swlzkEX9P2SqGePuLhgAVbeDp7E/ob4h8nROJHp7XSX
Us18FT3/U73Y9lbjBwQ508uHFczDIb+ZfSvis5FEiW2LohDZQksyHCv9hNuoPtaW
7rtFjRJ0pjjCTqMZYzt9kaosVpLphsVqctjQMhCmT8kN60lnxE0bzOrqsaZGlnlO
gZFZeIuOSp0uUfZhm2ug558QTXE2Wgv3CQD/xzHXUpYIUoQFMmmKq5fyHXSYnkvk
TKLUkbbAAePvoEuWoDTb4Jo1iNzju/R57ukbhidzAwxn7sAvdgTvkX8hKQhw689m
iu9lGNh4hlP8AFRE5fzt3fO3hr5YiMtG9qF3rxwumog4iI7nblmduPG38TiUYHB8
JGBL3uOrZONKay+gGPQGPikSaHiAyXwiQIyWj+Ns0PG2oT3ve+XKWQ1xPwLMMiRn
Zc7fu3ZwlrySQbkU0fo8Ls5KDLOBVAukC+mtFoqIUAd7DH9pPCP/r6ckvdmNOrmu
BuGiHJxH2gPCa43GmWhYE9BYKMROq16Yo3a5ADtk4CiyiIj+eVQIKNnpd/4hQzbR
oY79JBrxnCVTpTvYHTO7fjq2W2Qlx8OSz/fD6izAECQZ50K+1uPswctFwC1nxGA8
WZCLYBhHYoVqlcO1VTqzEiChjeKSEp70s0mLbNrMBpM/chr2p8PMIryxV0+zfDud
STKtjY0XmZKSvdzw4XNIHS6v9K7UiXlmUQ0FcuebJjEg1FVlwJXlK/2+W33K7L1q
Wt4xg+31Qv05h0UyAZ0gYYNds6hfR3K0Tt/SU5Pwto3eTkq5YjpIR/OmBZ4vtgW6
jccPY+OaT5HhnDywUq05N6/dZpuHm2cJDnQBxQdhqDo0ReAkWQltMkbI96yABe/F
+/uueWGCkpUPE3cJ/GeYPm3BeZYlaRYjh8LTCyYmo12FNmxHv45jp6y+VOEo7utX
kOnYc6WrqDDURaa5kH8oPqwFEIHoeUfvTcyXq7OvnmUkSQlgpF/NLNZOt3R5hrCV
fYEEXtPwRaLSTKG9Tf3Jddbxm9fi9R2zURmv/zP/7Ur11vQ8bQPFQjt9+SQ1/KdF
5RXMZ3Ax4FDeKaoeAY+GMBL2ZNnttxPghdQmgC35kNDz5I500+QkcBvg/aKnak47
dyv1HiP6JezByvmG7IvtTkhBDoYT+GwiyJiR3x25ZKdoBf2WlLp63oQxjJmUbda4
TokdhVECEnNhUGziFy5rQXNUqMTCNEvOVmi40Rjpo6ibYMBuZfrC96Bq896e7XOB
YZjzrBgj3f9qdOk09ujBx/GLFYKqDyhT2SWCF2IBIXaOVv+XQWQVJJ0pYr6OdYEa
g8fybt2M5nMSIbCFiwqp1+rMlmPnEkslhHdA+NOimq2DvV6Gq17cPt0fVnqnh3jm
DX38+gxzpIRSp9Q7heDv3GAQZqBXq4bTwzszPqe/HbyxuB1t0OZCDc4aychN65pE
HtEP+Tu/uKnbMc7GqO2zkgS3rLWdf2M7t2yk08ehmkdn4vLM2GrgzP7Y9+gNE9W5
2Yg767SQ9unmTlX9pGMAg35O72Gsvu5+YhTA1o5jCQN+SlvZiBmQK0/+cWycVQje
/GfyjsLeIhfPOYN7K7ZZ2PE/MHms39I2XDZh4SP4x/8+AuYLhKOLWqtrXp76eG81
2Xl0nIEngGrkUm47X6YajnMJkh9NRQBOC6UgZTlQwPzSn34IXTwSNL+bMUjbLCBb
EkYgWxxfmUg0OCxKG6YnoKZCM9AnRGmq6cbtXS8ii7701xmpPD1VNN8XLsqbCiwI
ZVDymcCRQP9hC97pCs1EItRGpGWmYaiSPG8Gs3SF7Zy2Qs1MkxoZau6vPfGQu4wH
2kf/efDV4HgrZdJf8EQKGwqubHK2QunuHl4pvDOG/UsIPaPan1fnwRHWzA6TGvlV
GsX/HOPr1E2sJuV4wYdBybM+WZMm1yuBJRRQzAfGmdHh76Vth9T83Z3DmiTfIEPN
Es/rxTourhQuo40uTXzcV0WYoVnYZ0CbTE/NuxkjrigNCx7DtnysutlZd7jls/UN
LcrpuF+Z1KdWcaL/jhd+4IZ3bJmMBb0LWFmovxNGrY6LatOhyoh+JzRLp548r0Pw
JGTQGIR4XojCAtvn4NRsuHnsaMo/mD2huO1CTencl9iZoMbQYfdzVNcAtLVTyHYX
4bVsPZKfDx2zbasofeVbUNNQ01yqwmfmT0GuD4RhMIIsXLqjclSYAA42jeJzLIm8
bYUNswiM/LllX72iNy1kNdBKFBJfygvW7NzWA/jJwei5QxP2el3BlNhsO8N8/GVH
hGDnyE/q1qvIgYPKXfEUVPuxJfV7Ad9j3mmEF64BaqJBjor7jse8nKg/qIknmeWo
T25EWfgHi0S1tkglWfzHMEwvmYetSftukIiLVX/H3FHEGALKcwKLeXa7FXIetlFg
3bAutALKEVLosvn2gEJQhKwnB9BNzo8BWduGDUhqTS5sjifjfJ5woSJZiFL8kQDW
xtXYlpoepcIv/1YqPYA49DpxZOwcX8rMIVXyzJRnuXzlZbw1c0t9945eR58Ypvnm
PIvpF98Pf6WRbirB1OCVhLeHTH0nkA+/ysSW/B5uZmOgs1BxeO4/rJ9Rvg2usiv7
MZ4k4v24nGFLyxs4nRHsTv2vwnJbYV13itMEoqwylg+QBxgW20vG9i9LZNsxJaTq
qOH5UiELMKU+5/9hqHFziurIqL582L52K7z+3vmWjz4Dqi4F5JE7obPLjtl6woY/
HpoL59L2x0/n9GYm6GCIjaJJqAXWTattOpJipwpLZGu4D+IlPleki96rkcoSLSp2
qbyE6R1dd0tc23uUwbZta/yyFo1SuUh7ALrAKuV3kR2BkfJ+rXot84oT0IsDaQuK
ofOJHNu9MAYMXwSjb8N3tO5eK9ivGb5hnqe+ht3zY7FTzGBbmZ9gpAs8JxT0JFxP
inqOzyk95OjNjvEJfqxohLWJ8GgIpqRikYacsSUJ+gXpT/9v76Rqx31XaJ26wUXJ
oKfIdFPQVMfjXlad70fXpVN7s7bqNALuuIgMIF9u4rhrcMvPLbGM5IgnPvPcIqsZ
xu73NKWVweXTWN58Rz3NJOEi73Id5id9vVYktVog+QjKkUaXF1y6yIMamYxo+UO4
gN2H0VOKvmYyJqGBKatNJgnFLVuJ2BxC0RfK60FhJb9uRRa5skbfLLINaxP+fOtu
sV97JWI7vGgaoo7e5IvONCiBqPqZt4z0I7bzj/DBxlW1/v1kAc7aq4YQvfg/AZNh
aQHmov18+WJCYVLH2wlQhN+I9xXMqqNuXIeMRhlA/h8SWfB23nl/WTdYqZPq9ENn
2WgLL7peep8/MT5EHPNRWYzka8kSxFDNUavnm+vqIkstkz1szkr8CxHMLoWZ492+
038JVzPtMiBg/GwgU9b/iomRFh9U90C6wSDiseRUOGXwwpjH0XZ7I8lWFHw3lYUJ
ZlSsFWUVDXJEQQvsOu3Axjgu5HC6p+aCtOTBxRPbNhbMrwlLhAhJoQpsRiCaJWE5
nrXbsP/SLsVbz00R8GCheT/Z6Z36IzyCHHt5Dth23xdKDOW93+WMe4FPbzKF5j6s
mH772hTIqfluDXdH/HP4N3mHyCTDYp5MlObp1qdEyPSpl3EQCP8eAGser9BfHCuV
uWIVfNazj0z2WiYkWJABcq9q4oBFjH9ugcgQHbO4qS+nzWywJnb/oS//HcgKHxZD
c8FAIRdx1aU6ajqx4GPB78JVYz6/6yMYFiBx6EKZ2NZomZ0JtJp9AFZhet32l2w/
p0KJIOX5Uga+tI6bEkp5GOSLQzFmfaphRljAb4IC1HZDygsQRqj2Evn2/B6+xJcb
ts2zha+tUSmifBRStNx3kmoye4pM2Gz6xqHHMI8jgI/B4rYMa5zKam+Z0k0271I0
FWQMmf8U44w0gvNXEPN4/HNTNczSUuZpskylCZ75zizHwk1Ik5W0kh1FRTT/TWPY
Q1If6i+t4c11NaYxYGA2g2KC+A8ukHhG7XRVfNnjuyvrIepsD5l0fOmyuxvFSwNF
tutV2xUTSNIxOi5sjVTKJERBDmNc9cFF30qKHfgJcwJh+rN63t77CYxB7r9LUz07
D5ZErvCyK+mIIPTdwfnY2iT029+qI2jQojls544XoIhctIxduxCgFDotX0orJnaW
FCwu/+I69FPdhFPEjxREbi5q/k8qwd/qAkvLrVcaqxZejSGZr2ub5p3mMdglTccA
l+JUhFdGZ3bgUL8hiwl7V87ySg4RVFth0EJZ0ki/KzHQ015wU5WfTidL3nKROkHa
gvGfmiRFTXuFBxbuEzcl89vJ9Gg2/VMxO5OrvMrD8SHHRN5vxcjPCbpQCR8kYd8A
axoVsQVbz8XpvI6VYnGHmtEmUlnARmfYDoATsTfRg+ENn1RhXvjXirXvigSb2C6I
2KAeKQWbZTEXS8HuZ43NGz7D3cv3uIMxppgEdBfRtuSC7wRJ6cKev2CLfcVGdRJQ
uo2aoulhv9BOwQhz+lidOvE9emZ+MmTKiid8qScDO6xvGMBcTaTAKzLTMN2vwd3L
sxry5/vgQ9cTU3hC16El21UYkJk+prd6adaP2QtjzJq6qU2WzuiCOphpsOcCrl/K
aJAsYOdUkqtbpvlq07iSEU7acqV58MkWNe27lPvwWay/wpVJj4Iungsgq/IKGaxh
zN/40jlCC0iexYp+5dCCEfxl9x9i1jZo6SHa25Q+kolGOhHcnB5PUqrcWjTec5ng
PmLabLLVH7d0HXP/orqU4t87j8sr5nyBVvOseLdukNQGjLtNWOPRNIKkD1JoRNcv
Vb3nprrkDGsylzK4FvCFg210A3Fjdh2daMeelNOj39iep8IoA6POEbU1s7J8+nB9
r/SlruLOLuWYnF0/2vx2pPou8+J7a9f9B6qpGyeFLePT43YdldyGEbsOYtzr/Km3
nXz6lFKP+u7vq7PMgxqxxv9kzU084wFms+T0IxfW+dyGSQbxkqbovqOx4x2JU+EQ
av3m4vG9mXzcrim4GaQaozS6ppzzeR46TIPAvFyDfo1Wx9/k3kmLCdaV8gRt/VFq
ZBORd8TykwlgbOWGnWFv86Aysxnfu5BStmt/lvIg85KjDIqQpbqvOfuH0G9aqFiP
pqsAGTesy37psLeR/8o3LbzAt8bnHZ/l2WKHYOFrL1MdRljruCblTDDZntUrWREO
vz8BV4NgqdxYrf45Jhr1kk16DusXU6Zxa27CpHglhIPOKscHPYPqcJDo1vvqU8by
H0KQ3Qz3weA5BuQUD+h2a/z+HnzcJM9GMTle91gnh42rJ4SXZTbM41sWOEbOXpre
5URDOzWvQ3OMADB6lcVE2pnE8i3FFIslRpxHKjQqPBgfyYSu+tqF1Jp9yGLzkbKE
m3MR5M8vDLVa3klPBvp06W8DEt7bBDbxSa3Pi69ma/aMTKnXBHvn04ayBACjfd6s
Ynekq8WvcZZnwpgQQLJhGWUYDdqncW5Bmr/XzkvGEGK+BOR5v3qt82icLEEsHHXZ
/FEcSUwrWcfPWHiBAhBo1TAYIj4zunYc3jAb6AFkBRmQFgYlK5mcP/Wv7gxiFBv2
HEGzhC4BPDLGC7SquX1iqYo6/GaqesWaVXDXE/l5NNZI2KZKscjnYJ7ONRbnSj3V
kWq9FCFD77dmJyHI58ybvwE+qeHb4Uh25uB6/glY8AaZgz2dIKpzAf/PhbRffNO7
k2tce9bVLrHd4a4lXw6fUnyPy8CGtrwtoZmIQNj0+fnd682ieploOsdic/ZVbs4x
EZpTgv9e7HceiTMcBKPVSo5J/paBCXxUTDbGf00S7pnkBSe0DSaTSuSk4brmDlJo
xDObJVvx5IyJMoFUnKYh7E+eW6wz4jk8ZGF+JBa+KiDw8vkR6YvHbXcREUrIsyRU
goO7gXhH6WL2m8+yK8dnXjqv2PKWzHtQCYDTzrnBLTckkqYmmfhdVrsqlolJOv2B
GzfeDA75r16sm65J+S62qPdGlKGKLj5sxLwywbI1Lpljgf6cAg/8WGQp7TvZZwCz
vfqMKGhm+bO+rSqKnKu8KNf059xG2kiJQVBzkZLoUXY2dxvbubpqf6O1JNpNW4Ot
f0381Vv+d9HOqNNwbWq+BOHQYxVEYrmg+0knMxr2NYm8wQdpcG2vRL4jhLlumlKO
E0mvdo+oAUQnhmtWtFIPQWsYMZ9l9HAPxbXCLCnzP1imH3tBLO604m9YRt9C/K/O
Y61SFI5OILtcDN1RKLiPXzLQs9WSF2v53E9BFEqS9XknAfxWL45lwDzUHBKOEpw6
DndecAaHvTqq2n9LQ6aOGgTVT/ZUfyLhSZ8382bLt6L8b4sm1zdoqW2BJgVZOgyN
fV0prF00BqltVy0BxBy4tLBFjZw11cM/RKms7m8yHrGIieREFJyXPhoZDAO0khtD
0bQl9Ogs6/ekmS3KHeFt8s7F7i717e6p++6jzaNDSiBX8DC1y/6JPMBkGqfgynJ9
2vVzvZCeqTT9TQF6emTnlJKMC/zRHM3yr6xozGV9SqhbWxZJxORqpUu1LUcX0MSN
49F/aW6+E2Ej6VsraaiUYL7Rw5DsChLH4UIUPU2blQRW7wSpQy+/ztWgESvZSM4b
WVtmexDE2qGEY9hM+Pgc5TsnIdhRcbCbw+uqKDVvPWVT1S6BejK8x5+FjTzAiEzI
kOCscAyFj4dsjD9TIf7sr1maRa/rfQsefeE7aO6jeLsM5BuwVimjovrv6bqsUMc6
9kMEy0+rbiMG36jJ+UhsGMmB+gQbL+VXcAER9yuTKyQbZxYuuEOXETy5jZmvgfZD
gwVFAGTFRLGuMPTlNUqDuUT7Al6w1uXEu69GxqW1pSCnXyhbN4OJ+TEuzzYvuks9
30CvRZraiWzZ9HboL3bRWrG7orQSncb5A7FCG7Ww7S8IfByNfsxllfPLk0abi+rY
JAXdGQSN0XD5eaD7MJc/KjCHhmbObtRuZ1XWEf9P9HhG5FB4N7qPTQ6peFM13UE6
xf94dNGnCLNrCDEzKW41x9nJq4axKOj28XSIKv4BxIYELqGNyVZkkUxK5ue16BSO
gtUp3qfGtz+pHRtMH12sTWSn0zofY5qu6rA18cLDmMrWA/zRdRdqLhYX29U6HkqO
6pl7L4iL4l1kb1zsZNbj0b5WpoFIsJrhL30cAniffqclMdvO9dsW/hn58JM3Ybo0
/WSBqMk/9dgNH4ak/2K29YpEXfVRLhzzI0gFB2Za6qdk0+J859h37jl56q6lXvIF
GFgf2nJyWz9lVMVFX9HbYpv1w8rRTLuRI1iuXIEjW5gu6/r3WIhd74GoLgyhxpQu
ZnDs9jDXXx18Ac3oAG6WPOE4GRB/TxTU092/VNsSJdi+zkPIXfCTniMyQtgY2LT/
1VsLsNqHNQ2YL1MWSDgPMmJhhqGXsULrIE8dKxS3WCX70DOekwBt49l55ypzNdKN
NPoxGOV1O1UBRXBQ05qnNmTa28+sHk58X8q0ZeTmB7bDRf+rCPEmK0LTa/JRrYgA
+nXrl6J7rbhAxcSh1SuLh3gejnsDzfE3r3mqI0vJljREFFXHjAtVXS8nAldRmQsJ
15olIrX+r7kk8kMewA01MtpiwI/MdN8JG8Gcpq6HG67a1lcEXCrzq3uQll60XiOC
krfC9D9RprvS1mPC0Y/tAbYQwc3kI3b8hcrEGxksbAS7SevxzkuyOElAz1cKEkCZ
BLTvI3tdX2QYKh/wpAXPcXtEAsgAnzMwKbTiO7rxy/XAGhgWMI4ZEHvD1z19+pw3
Zj9vuxRj7a6miZWEP5CY3q4kQgI0zfTSIhF4+Fvdg9VVPB6vMBxMNDCOd3PwIZg0
iY3iucP9XSkJarxAwJ5xvpK0bGBgHbVCkZTn1PlZbT1jwa7edSBYmvJFbamRsxu3
DbX2rl/Bz2SEgsMz/u4TX6/2IprulHpyHBvpVQv0V/TayRAMYltz9xz2jIzp+hCL
K6JS5NkCE04FreT0eNCNblwSgIyHrp1yUXG6tB8D4P+s0rLBwE2nbMCcVrWsTYfF
1uc58YSblyY7NOO664jW1odIRzPb0STdsqIrDetjO6VXLr7AFcEEN/vXzBHF3O+N
BvR4sl/zuDe7L4pcwNDrYFVIncYvfsAqbAg0cGkdBCTGm96d2lc1DN13xdAnFgOl
Grde+MgZSXN4+QKkr5Ok31N9ZXa7OjQ8bifhD5fv6TncSgNRwpnIXsxGkxiZ3a/+
mXC0kIXr1SptCJt5xCaxdU+yNPrFFduapUX9JWlcPpz82fd/MsU5HmPKxnEbSSro
0DpKxZaynY04dA27Y/htJ968q9O8X0+cuJVSU0cQkaHzd6QZrnT2DtnOuUnpkphQ
qs5lZrvxElcQ5YqH+UOfOMkaarNul9viBpfCsuodAh51m0JbCS4V6g9WMJYULfo+
ut8iVqacm2+tiJIe2pVtxtUQvddY2jdzY6tSZjqLaJUMa0vKrmDcPQ5FyPdPdBUs
RV/agnbaodjKC6qPR2g6GHIoq64WEuL8AwGyToESF0eEE7xV5Mk9SktKc/Te2dBE
Muro9s6XrYk7CKkRJcIOs/+cvMsq2Qij5g8Ioqn4jGbW9zQQYA+WdLqV2zkXt92J
N6ozeSCNu5+DweMq3JUgVUA6bP4KfPrRfexPw0aMTJFeYEjMmVLYfTWYIC+rQLjQ
ncirHbFGnXI9vMAt0erX8EsOBxq4SuCu/4LNlpAnM6SRpTibRNrmPYspB50zu2nx
GmaKkZxR+EkuC3o3XauBNhxC7cpVbvkvAUG9yXSzjDSkUCT7qqJKWgtBn2Px4g6q
vhDdvAQhVVgjSvSLhczqpPEouJFZ3I3CxwchevdxLwLp4CO5C1dFQ91rffiHIK2M
X0LhYdvvhb2cX826ZMR39Fjy4kVO6Nu7t4qbPI55pC0n8NeDWYGuRV35nqYuvw6q
MxHS1GrnExTs2XltlaPBZtG5dOYbf4YJ95QQqR8bdc23baXxMv8h+S9FaqWwI2ng
K5klMOVJ41iwT5zNvCRLaXROnpET1oPauzwpJ7Nx0uR4ziLXtFwbo3ENQ0TkKvW6
Q9+QRyIhF95YwoSwgEdMDWGhVc1G36vfyHMWV8NtaGAkIrOnw1I52ajrHt3Neexn
pb15QV5WIonPFg1rMST3AralMuRPIl2wl3K8n8p8sSi65BlUr208kspo7dROO3/X
Jm/CFlBlHffeWNZX2+cbyfAtg2ny3lC4T0AzYOBf0RP43IdJ4SP3wCvJJ6PhMYJg
18d+BdPA0UdaLXFk7Grju/4S8+ZtjKqOr52dht0DM0GgWsjwnlaBVSPpW4wBBqMb
VI7JeMKFjhkhETTu8+bNNJ0fyGAVocl5K+IRhy3LDD2A8PZyE+Q6yUeQZRwoaRcn
2x6b7ddzzKDmJfxtTipwvOQ3TKRvm3YOUJ0fMEiquvQmXkp2hk8m1adWr0c/ajtl
gboFIVQ7L3plZWLr+tNQQpXVwZBfpLnk9NhjWzmHZlfQxJBpqZYO/bDOPehIsNHl
C4NsYE240oSi4B1NQakRqCJ92E1oda4CilJ1AIhbBW4k9KtF+ZxEZt+eqWy1OidT
DjzEbVGid+7nFAktQ7iJGVPS/WzJ06pd7ERRRueT9R14O/Wf5avoxI8HxcbW6Pdo
LEm6on43pfVQzmvbU+LjZj91u/kVOvhaHZGu54lsgrqsCHn0LOAx7Y8tFN61zk92
Vq+RLX1+p2tddJPIQi8BNsF2MSyai7myoPV9p3x5FAbOH2fA33jlzKtQhgcFqtRQ
tM7e6d08aLUJBA8A4WH6ZbekDMkEwrBmJIwj/D5c6VTqfTfdiqd/L/qd1K6GLSff
co1vJ5MGOM/f7zQkMnQ09T0YD3mXV7lksftAkeN+2tFyTiQSxpzR0T31KfkVlEE2
ER62O5KeSAK2lPtW/vACEijgrBZ7GF4yxRPpY4r0WmmzOJWW9YsYY+okd0jw0AU8
10BCfvxC6OyoSxKUIfG15Klazx7bPWJtVBfvtPThKYpFveuh6YUFISTyo80MdNuj
ZVm4BNRaIosI3Lzqa+vW/e98WUX+PvrjqiyLqSsbXbetGpTEFE7Ipom+K19l3DDr
6r8eNAuLSpBR37B3tDZRCQJIx3bUv2yZEGc2kf5dBFHogQeeiJcfXx9O1ak3mSA1
ZQHuR3QA76qNNpuO9QwdBuGwAgjEeeKqyC7XsJHzZ4psPm/6G2sMeNJIDifJQbcf
6Dvv0zHbR69XTg10vxumjGm5jhQqHtipDleKy/MawiY8a1CntOuCG9TYVFwq4lvO
c5mvWrEhbk97wxWK+g3KUeL6MriLjxErYn3cnc16i0+Lecgu6ywmsl+zXXp0v+Zh
OVB6VTpIYa+boQTH4uUQ9miLHKknOn/ZlXMXSV0a1DcNU1GX7y307dAW8AkdDHZ2
Quvb/CFMku+vQT/gQD1v4YKyyh9QSYrwrtuipyNtsfdD01dQGLuKxo/3Va8WmSSc
hXthfVNofQ1XyPUn06sJwUg2F7b+bAqbMLQn2WmSRK1yeHCVHjsim2lc1u3TlxaT
tAyxF2MMdra/Mc1SRjz6lkkUif/x+Bx8+7+GgYoGETVfb6bg1Wvf25fTQe8bLQ2y
mXT2Ltxx0M8shp6ZXDLcwycJdUDBVc2HifkEbcBGEZLGiCJgG7mA67pgOLR84LFp
cpF5HWy5zZXMuV7a5cirIxV9GMryb1xvSd2AIQpCYVrMPZpluZ1EScV+kylbDpSo
gU5y+ICXDITxGYRqdLkMTEDqMzTdbnpTBnR1xhzMFTuVcZES2xbiF98dTwVF1/Mf
IJzChIbw52yyfgZsflo3RYHlzMTotU7AbOv04OQLDpCtEqnIMAjhjP6wgoBYz6y1
o9+GDyS+KRkqIvYeu0tIhe38NS9kjse+6fXs9uQ+NaWOCJd9Ojkw6xbQR6rII6Zl
l79hAmPUVXXVhnLU1Zgijefp6QbqbGatch1334YK2LPUHjc62c7oWyChbNjqoqE8
+Pv1Zw8ioKSim8gujvjOJuUEv/4t2EwHCLKU0xSlRmd9OGy7TTAQ1/LxXulJ/6f4
EEdXNXPvGrd3rD/zQbDGxYcMxY7Rpx+tSo80/UW6KbIwbBUfmdeocJ4Js6Y+Pa/v
fgAWw2OByDG/HHfxICmC3v7lqALEdLJ+0KM0ng4gRBht99tjCgyz50PvzAikahHA
A9XieHLplfT5h8n8y7kbOrTLqrqdaRsv6CgLTeUUCF0eN6xsm0Sspp/u0MS11Hax
HseQN+we4pHlPvQ4VHPv8dySnh41ArIMyEfSVtcCuq6MpBEKYPZ6HqapLFFzz0fs
zFjeZorqXG1L//UvWQ7kpatM5BtkkSVF86Ll4GDzrwMBybCOcz4CspO2T86p8q1f
TR4WeTFUBIj8lIBYWALpQ8tjWBNeaIibXsD1I3Gql5iy7L/jVct1GR+z80RkdWmZ
2y69oyozTp6OecgWHw5lL1A+QQeBjrasn5D+G+bBKCp4soTaOkAaPqrLZcl5tUl4
nYm0YEC8oVBHIeBrFHU4yyzia2j32I7WvGcNnftdsAne/7qxMBvB+P1FlV8ZdS18
gYtLABZsGxP9bygGFce+QTep1ETA/5vFi6JQ/jOWu7xQAjM0gpnLMGd795fJ319R
kGdzgVC/yII0/ESoO+0TZFSwKfoHETQfPYXuA8J2Fz/mtewubzDWkjQDshYN6spO
l5wB6/JHeTMlFubIqrazUrCrlFSPSXKvwwClMPljn8CWd6/TWIqcyjKfbFRQr747
dzw0d9ngPmvD29juxlKpHq4YXtOGzqEjQNQ7gdDLeoKUoJX3ihTYx7/S9GYhNPiQ
t450NmyB+q02qvh29cFFT7pWUNRFIYd+WJngJ4NdMZqiTuFDW/rIcuM9YrpinxAi
hB9r7+ftTAGiEIx/Ts5Lx9fzS3FYdCok2mAI7ts3Q0BePZNV0MPWAenKb/Xxgbt6
YeZrq1N3Zdqs54Q8viPydGfF1HW2OMZvQ7R3TEkdsowJTcwK/qVhY72TtgVcOD+V
MuHE1Jjxx4XmoGmFo3ixXQ/8QJSyzIAJbTdMB2zclox1t1Bdo8QQhqGt/fRsHlL5
5fYlCArGlTULTUGtQNfhpYwJxbIjpfZfZyXAviCn7UMtMEX650Rt91yL4lScJbtG
8QUvXDlycm30nGslMURysfuCWzxNQ9zgK/kf+Ylwf0qSArUGCZ6AaLkinGENWYsl
Lfh2f3rHzg5MsW3hOwTcsrc1I1lDhIrHWgUtS/n6NEWh6sV5eyQD8DXzy4+kWTer
hKTdP3+nJSNcQkuTdDy80swY1EKr+Sj25pf2XyZdAS+MU983yUS/g4/vWeKmwz99
qsbBJ+eTlXlmXOSdCnEKcSZ6x/nU6v4ctpGR6sxHSi31YHplYRhv47W8M546keJ3
u+3PdSKaQi1//Pb8K9t3Xpsbgcz1A5uJ4Ypg0VpBSgY2CquT72MYW4p+lbcF6DPi
+90hdRe0gWUr1qi5hsNeCbLGszwEpE7F9c8VxkbGHgLrHhAQXwbpV7TedSkWKRlO
x+OvOfo4EvbJqs+qAlOOrB2tqLpCoNhDNh6yiNfn++CKsSKg7O3mgUAx5x7rQpZu
XhBt9Y+NA6DJ+pI0c9ZxSvNLPeJIhNoF3pakS2H94LZpwpleJvyEblMG8OCsFyqw
oHNO2YPHyrm1q1+b0ftVXINTMrljAHKRnNyX4utLWleZ9Uggw9DrAyxpA9z5AWVy
13vfpv6f8gownFuw34co54i/dpewUojFJvQKpcLxWUrNXkh9Gev27YnKvgJmBTop
Ly+dbR1yadzzKZ7q6WQFZmNvdJLOFxbvOcjfTJyz+GNRjRGuvS/TL4lVTWAsK2ks
gs+AaQbVA54E7df4sq18HTPTwKFjsnfjtChu87fxPcCqC4LUrloHPqFHySu9nBxU
t8K3TXMzX81gnCyPSJ35lPTIKYmTHrsCyRg3mkyPTCCJaEZoYTY6ATf6XQI7iNzj
tL9gBtdAG2Eb+59HgOe+UReU+mbVt1uiXMQjH18Sef9V9JM7XNpveqKLMiIg+JLA
11J2VPLKWCwQOGVCDMOcWeIb8qVZN29hBWDCQEzRN/eAevPQmSMZFDt+6D90pvO2
LWpQqMiPLtsL/Em3EwHvLzRyXtvcUV+i5mSt0gdU2QLXwFMBIiv3AI1EREoJUEgS
HoWlNlNc0wv7myROKhWpwiNQHZty1q/vFvkCb2zRuMJSpfLR3dxGSu0di6wOoMpH
TlZLw/aZ49K0qGOJTESXdxLEBgbPEigMizO6YSqvrhIrVRVlKGlGUR3+vPiNgv2s
naYV5kSH1rAf6WmhQMjlfokLJhHJUPMUyQkHwJzNsMGkVZhfAek2oSvMMpqnmM+D
0dLL7Pas13GMFARcgJOwY9gkJDtUN9zZXQAGgJ6uBD/vijGhRL94C0qcRLJspf4l
JtdBSYicqtYtnt7KSpJqd/FOWEJtN2Ya9S8FMqxGx6Ko6KDqKxs/tjTBenu4WRjF
O2urpFCM9nTKmykNmngbW4y4KAcn5e9H0bJex6kRxbw0FXv0S10CbpQytqHB+OUA
rFIQ/oXjTQGC7kS2e1ZOPfir5FaaB4CePhmHOcgaFzeN9/Lev9AVuZ+wzrmpKZEk
JtPJT+mK6G6RtYLx8950J7N4ahiw45meGlajRD+QxGpYXCiEUFxcoxpE4fLkBdIb
xlaO4AenoRtlv0XNdAT6L72DaWnCrS9J691DATkqK/tN+zgbgz2+a6K1RT4JGXfA
aiExeR68eduDcMfQbLYKb4wdTOipo2Fna33f8CFq2UWt5HGtmeSJg0fJVC8O2EHD
49ovoyb596pN/bBXyB9FeoKcn/eSHf8be6h/WHLoEUEycYNHmXRaEPVDXNdjx0cm
AvQHDiEIKUv0rxoz4zgErwPBNefGRgiQCuFbgzm+oQnpbI/vcZuAp2FvGzy4shPY
TuPsXTmaFVsw7A/ivJ7BfqV/7QSiCD+qMGOlylCqYC57APE142xIErNbofhxr37d
XxS/yZc8IDqD1f7OG4THmybb6t9OjviuRS92aueT0RhzeGB/VEhZVP+HlqHJOSxP
DmJHbHe1pzl9KVCCUK29GLHtXfm0XmlyvXDbwo+BIe7YlPNFPjXwWMw8nPBwUJUg
p/cTwMUpl6VEtWEjvYf4xQ9z23naNVzbnLS8F/siA1L5j1SfxoqNTuNdc7ilIC7M
dxjaiUpOXIGRazTkd9WeAR9056KQpAn+pH9CM3wzDfiECoIAjfonAnV6FLDzuWPS
plT5yoA3qeVOT3wMCHLogtQ9gIiwBOd+gHuMadiKu4NxUXlGx8HA6xFdgCPBItOX
1+hyvpBKWJRN7kNtZTpB7voRsD+mX8YIavhLlLEDNWqDvWQJkAwsPuLS8oUPZXy3
RZcba8/EBSbzzl+aYLBRnPgp7P/Kje50IzSCbqKgrSvqpsAgHp/QJsHrtyw8wbCz
qpHSsAkvBy5JKKnZPJMquCNeU/PNhkFWJhL/Tj/rAaIWW41DrGsled/3M2dWqtE+
Anc1dXv6MTg+l5wLJniFUKtrLKRCSSmdy8CQM/XVRGfP6bSuhdcqbk3Nengwj2tx
omkxpS3keeN0gWOPJEX083tkOz/uRU9qujSp6x8zSSZmXGXNCgtL+ZhFAlNScrNd
n996L9G6MmYSUSBB930aoXZ/kJF2+fqW+88NfUxfp+f6XhRP/3ED8jwF8v+AMXoS
UnsVNuDVCtXNFdm5r2CL/miPv3SBI8Mki/Hm7UV5bs5xSUfd1TZAy/UaCK2N04Ki
L6Wu+ki2Z2Ty4ocdPnn/xunFK8s5nKOhf19SZZpTtXHave3Yti0ZZ30tcQ1tSaJm
tPb5/RfmdJtVvuj95YvnVU+otOoi03g9q60a+1EyG37I8O1da8A8ubSUZcBkLsHB
20HJoaw9K6aP8KWivjEhiIGbjdz2ytQM7Yly7Zqkzj0kexvMyLfzShXWHGLz7gtK
TuCsoxBxq1tWUJnXkpAhxoBYQZZDz5OR2uybJ6VbOmuA/6JJhgctlOvc1R5fOBnf
gMPzkz6eEWtWEeJNMcrSV7F3xI+tpYsldSni4p2xygs23KGS/6UI+5xwk0itMkbi
yXEiX5CCd2+rrketuuillrk9MARDMxZincIWioFQF1VOebRVxCaErk7Xlu7/cTSw
h6ZvVILtjvGFvuCcDpooSnxaL7fqYBiqkbYgEZQfYGMMu3q3Fvwzy5ogt/d4OSGQ
CLQQme/FouF7XW40RGYM23imzZv5fuVoQTgP+fDb9FhKzCeWPeGaRrqAE4QUebVx
StSbT9n5DiAIuuomzZ5MiWLqc8y8b+1Rinhfqpg4nlEtSl3P21Hl1h+b5PMCYQpf
Zj8WQidWfQqDdH/bCRPynz2JC14+rWbDV74MivYpHyW8QcBRf/sXA/p0nOzRrf78
YA7mID9Jspuyl38H2bCVwFP/h4EbCyOCC+Xj9eUwkl5bcy7onH26YoisFkyePiUz
hMAYU27YvoQYesASAnDGB0kT5UKD5keLkgMMa0u13cNrJ5V4hjxW805GGwSgyL22
MMgh1ONYdaQSICloy+5LtHqcUtD/EPEkp0gHfjP17RWwTDQHALg4I14YwPhK/xXT
ATTQrx0m7safJh/BqDXqzD7wrmRdc9D/VKbe+tQ2l1MDEkzR0YNDoale1Q9Lbtgj
mxLh3CL4BEjM6raJs3AJYUOs2DMkYPKTX+Ef6GHTf++YHiSsVSWtd/aeBlW9kmgg
v45l8eOkIQIyFLAIYdKJOQQBSc+bk0sLKJD+Foz9WDk7idafDSXmHoG7yN21ft/C
e8ghM2X6TTDx1nsFstYAc53KfQYm5Mu3YtfA/GMlr83la9wp0XYZVhsvCJQMUQns
9PY32RbCzmdVbGQylK4LSd5rFadaKORZ46oYyOCSkYPamXc4at7Ab5gYche7C1vt
ZXBstOx0kJPjjawOYKNL5CaN+TKdq/o7kghf5Ci5IckHqJcQF8zOUxToQZ5JoZ2k
51lr3lpe4i8hw3u5CxAvBgNKQe2KUPY7fimwY5fa0z/e83yidTWxOR3toDYXhx9L
31d52sDznoVJl3vWoKI0XnwUSxHMXh2uurXLtQ40yC/vSRAyZM4cGgtjhTSRHeNF
xyXPiZBkoedLNHgP9nTUIu2mbhrr0QsAv+4ieElsJIln8itTzVzmQ5vaX0HWM5gx
7CmHJhYWawWORDwc3gOdRJSEceDZJDLedBpxpcUcLR6DmJPiA7+80ea3T751T/zY
X8rFP0veWcUFMJWdwnSI1rw80qZm9ZZ3aRDsJoZQq6ZbKQgBF5UZUYqrwF8oCXuV
sDQHcrTfbfy6GGRFXUekjiisC38QTVSb+QZNQ1rzkd2LUsgIf7OkS/psoiSYEP7u
71gk52ScqJWDH9qc2pzdgsDg0RYstmO59h4dx/yWkmrB0y4xxF5N8bBOuQujBbVq
sJBFvYKkz0vIkh2UCe5GIyWHpese5F31vxrX4cndyJA8nB7hOeB+7RhUiNIN/f0C
LyzTJlmT13Hx3zgZJTo1eufBtFZthULdDKw/9lyTtmKVxJ0CUwDkvBx5HZJek+k2
g+ZiCqepxYEs5sE6bdjEal23me2mp3uHl3IguGLW2f5BbaMWZ+Y7mQfUNBYUpjli
xg9HnsbJUbPxLeWMa0e7pJh6nLoJKwTqiSB2i1+M10Zl32k4nkw0mRoNoUhepPKW
uDj0DUGfCSOt7uiKt6a32anyFWoK0o6aPMn1nQIOVxAs58toIv5DrMAFvUGpLSTW
xZXsC7nMPn/XZXdwsYbkQtsEJEynFA1l7/xfBBXESFjOAgWrWS2kozOmTA6radhq
feIybSOiuxbIXCjZrKMy+Sxs1AwBRacDRBlMWWraX6LWe1hy/Mn8jIc2+RS3EmYK
a6Ku5VJfd6rQojDD7QmiiH7Y3ZWLe3o3c3L4xrcCCwG1G2/a+iwo0gk/JG1TDWmj
j12XdGZzIuSpaM1SkZ/nLDra6zmaGfZrgzkrc+UNzeuL4FIKTuY8b0AVvovoR+rv
CcRUhLgfgBsFogJW6LDVUXoDom1JYw9toj/WE0PVOWMoCAv/2VctELNlajdj7hPb
rG43naBg8tnm7Ux9E7/c2Oyu/SwZYrKd2hnMi4cW4FbxZ5tWXcwutrjbtIAki4hI
Mp0Jt/x0Ybu1ojhrFXzqteGrkJIDE5BrW7mTY36IGJCVWRqgkXykQ6IKCZhQ4MEN
rqkhC085rXEPfL4+qKBy9qEEx+BB1absRIavWvTnycn6p4N4aejG32YWywivAhmh
nP7mD+b4F81A72xy8censWTj/mBcF0oNNGFOxLBy6WU4pBw77C76u9u/f2wshLgD
PDw1f/W/NxFcwbgjuJOtpJBzxbQ28kgzxG0ckmwH1/kl+UspmkNU0T6fJzWhbohD
jmVR0pF5h6Yi4oXoUJOWx9PQHjndxyVlwUAoS/3CLeFCx0ek5/Sau787vI1KQW7u
u957osZurQqy+xmq71F6iDH+CQ/O2gt2+0oYMHAeQP9OmhfHZNMgBHF8mc5lGRg0
sZXC1gpqrm/zEQ9X8pCSzxvwBbxS9BzjNXsU/96abu+KR2nMJ6e6GE9NQFrLt5NA
EDySINtSUT0lHObnl9yuR0+fEyjG1tXGWPi67PqG4yHSR5MRae2BJQbJVaJ//BpD
D5iH+8mw4D5r/t6gpByxi714hJDV1vBdW7uNSndD83WpUCcqx6Tc3U89M75XlQ1b
J2lWqzwObd7d7/bDC19awtc0iFuhAj31SUaHpr3tnRMjV4/L1dqmIwp5t4dcdk6Z
x3SnBAKnUtBkIr9mvgpK13l2Q6tDzr2NaYSXN3Ax4lY9KThca5yI92wfsf+wxec7
Lzcf66fjmoHj6/ajrjF4BXzK7SVDEfJwv3z4GnI0VAGqIZChcb8M9dPRa++fFgyQ
2umkt1Ki6BufibBXNrn2NMzEwOpMkNkPIonr16waG0sTL6xs/dYpJ+c5L2TKNLtF
9yF+HoUIabXlELZgw+AA4aZpFll24Gp5q7E94n0TQVtBUyxICcZQ20QBEF6NTj/q
ID85nzPlLZF2aIkTWS8QCtoAg0gdcqDhIf7cvylzP7tcvHByZqf7QUxdlZrQAV80
ZiS7ya7O3JBKefDqKH6BuUQ6p5+wKeLc5NtJkTuwSzhg7y2mmgy17Xdt0JyZUNyt
xui0jIA6+VdUjj3qGfHqbFsigAK9FMKwfeuQyy9lRWOzySszEqcYThvy0KfC/Guf
+WQyQEvHQjzeb2zKHDN0dujvuVhfNVMv4qASwDvgy9HchOeVCju8WNbdKRUY4YJ6
TuDwyhb5omJfCCrRcGKLgLbHeSEcqbEVxpN/oyL5dvY4v/eJcId7E6gLYFySwkEQ
LHl8f8bvh+VvTLzb+d0FeoaMr9/+S1sk9E/zSWiWLXelzGW+k26j3yxqC34C+ruI
Qaq3yoNeu1sTEcSRZrqTFAEbtChhfrj3sKy/sa1NQ/FYh5kK7FFP+steK0EtmqJM
p2BMJbxLic9EbRAIGWFwQaz/wfLAaaC9vF1u6iE6v/HLM5hApMtwasrB0bYF3UO+
/q6byPK714sB3VM1Yi66w9ISZ9N0Uq6gUkywxt6wuxIH5/qfsr2javxboxtNVjKg
0jV0F6AnHuP7PJm8NzXa4FhxXXaDQYJjwBsjDUGRtoS4RsPyHunhgHMc8ufFkzDh
cuXE3yuzwdYZ93Qvy7W+sy47gJrqbfrOZNfg7ABSb2QTaODXqw4VOLNNuICrtpfd
OzY9+9JAtbc0k1WWYhaEHszJi1NAGdabFVCutL6ekPGlYPD1wcOYUuhaOAjI3QYL
l6anv7/XrNmIjmPfpwNaKqT0dURqkBiGljRyX6NBZDcZ2wKv/Gnpgm7TAQgPsnTD
oXMiwP7YPBPaF21lcxY6diegqvs025DQW/sFLj7/Kf4DmkAUGSCFOyiyuvXq5J0Y
rJvo74OZSGkS765LcwY2bI9BOwasJryyvMU0f6Hzam1rvVFPAXY9k/xuTW+8CKY5
WSnx0Jjakq/fmOS3mzMlKRG+to2K8kRlKvVjgzeomXzHh923oRJA4uM11khqH+EU
35+wmpsNpVuo7vzaSOWzFDtrf6lXa34ytycGI2Nds7NKCFowCnE9ulXslxEhOIyL
bi3qmIpHs5ZM8vk+va/kVAxJd1mjlueMYVLVvedJGXf1w+tTDkg/qHraf+2UcotY
aRa9Ws1WR58ppwJO64iSup6GnIFB1pKDnuWz0aBRO07HHNj1LeRDc1kz/CUzaqsE
t22JislGc8Tl7HeZak4cC1yhEFMmPZWr5ekxkyT0G67oPTFOyDwOrm9Zee5TrnI6
PDmbapDyfs8eifMtiDxqxGF0ahJdsqRWtF10PcnPwN/cGmL7NBAQJSadFkR7vm2n
Q8BGIi0LP/lsRwgKJgUiV01FLpd8+RkAhWSNu9+Fg317gBq8fVov+t8syO+0Etyk
u+2bk9zK2f5Yo81gGpQC8BNPDVU6nWJEGV6amHFdePKOD4mcsZIbOoiScm3BOKL/
lqA74I+bo1iRcnJeMdNkSsf98fedcSRhcoLuPe9s2YvcAUBEYqkZoI+8b9YMwiJ/
C21oRPCMHNyzNp1g+gSkYuzNSeifXmasCihaecL8YM7/kC66RRugi9pJqVri5lui
9RQ11GScQHBWxqLWbySdAvFtBR0MTceKQ/C+JWCOM2G1hJ0VfXLxNJr0PR8iUq/n
WbB3IKUNx28Y8Bca0Ts0egut4jIWljq5TyWIKe2KneGgB01Ho9COAMaBh7spABMU
nX/5I/RMKZQ3IQSwWeqhuuaYd1guXSSjQ7rtV9t7ZD7t3EiARzxOC1Z6D1B3xncw
PN1sPaBI4afqv8VG9zUSjUiC+UZitZs1Cvk+4tzJBATlFXbzgQvsNaX+l6vO9mbS
CHcRUrSQbD7dKJX2GCnUV9Gg1WOeFCt+QgDnLsF1lCJl6bVJFtzVETGw8MZJUgs2
r8VBBAHznHzd7fFyurQyMp7XW8/Nf/s6wZoFk8VERX3niPrWqn4LquA3oATlaba4
O/qEzxZl/CK1lczZVY0mAsGBqyXFB+7QTCHB+Kci8EtI7h2yZ4c/kwmvcIohShfy
EcupsTsbI6XjsA5iSA0ZKf5ABJPbP9URT3Cq6hnjJQTYHzT3BgqX3oqBa7RoqfDy
oRaZq53hjSgqyxgE9q3NZx5v/ESySwyRBbxP4N7AMgAXw2V3TEPSN4vP9SuXpRh5
QhoNHGsGdY7HixW2ulJkCdBPYigORg3/Mi6VHHXmcHKXfSBPfZ9pbJDFTQy/fx8T
pgzEhssnLxgBNV3rcqIUZLlPTNM9fJaW8LWQXZZ8wLgTcx46e+Am94xQ6WymxZ0S
SApEP7jbR6kxwW6O+n0Vlxmg2vrW3c+axSdFUEcCthEPVcYsCvgwtYVDx0AS7+Yy
HuDaD3Jw77tttFVDVuz1zTQt27pjvoEqaxZ+juObouYktDSX3oANonwSiYqRUysy
mySF88tlDJwhtqTaoMV984kG+MwIsdojWrDByuw91HmOJPux/nFyt13OxDHK+prP
lNtoWaQpiS7AAlOgRNeIrJBgrTS+XYIyhRpIhilEZu3BJ2vfjGBPVVQNIw5aZlkl
GGGmBkyIK3pDhRxOOSVQ+GG52aJuIX5QOHF16uEfIIAAxyVSPjT9eCk9brUWUmrr
KnggHll5x1T30knZXyKSYR4rGgPMfF4AsEUi5ZZoAwqLxTIWtwxUS4Oz0o2SiiiV
MzMYtThkoGPiva2aSDa1cmvDnCCJW8CYh3si9Y8CHxGRLkXP9Mj9DaNF6xF7exOW
gZSJlnOYqxG1Ppce+M7sQke9cEjyzA0QsQ0RiqTxvjgLmPIJg6706x/e5YfYO/86
vgC7lBnELBs2hYdIWwpLWrpLP7po7Xj1N07p0AA5L5MIY/Gw27hQG7K+24tbDAZe
zrjPXT1ckK/zu6lS4aKOexXl+XMEq2mgPAyRWxJmfngiBBgPYdykgS0mSe0VKlpL
QVoxvmsafonQZkeNKVwyw6u6RBa+x9kva398d3TOI/QsvuMsVfq3mUPFse3+bMth
KgZq/5gg5pDh74xBpaVD84y/xxEUwbr6YEZaRMw97NQdA6XoZyGWyla/5o90cwW3
gMX0OvjBWWYOjYhphXaLGYnmbO9Uz2Yl55pCnEPoHGIyrz94/Vqr2nFzyZJ9eX2v
nTOGSwokSUJF0SMFYOVp5TbNm9j1vzxZQdlRDOnUrcw5+wnWAKKF0Se1dfUEP0I9
oS+4d6i7XjK1mP1hayG0OaGYCusa7jXuNoAoIYpjYQ9if8Ef40Qb5GjZhUvwNWqV
MkEY8ysP+6lR9u5Y9KG4ccykFW2DekPUEYnuuSnWBCEuGPVxSV+ksDqEvuWNZvzP
R1P1WDq71gyF8RowtF++st9jSGQ1Gx+PTnUPOd1VidVTWVSm0k2mXg9v7myP+eKv
Hmw4qve/w140YRjZWNaL1TOqw5LCV/+MQ8WcNaJOPQvTjHLemcXJZDHc5L5/neyH
4wSmV4PgoynN/iHwBC2oFT/sJyxceWS47e6E8auG2OooPnmFW3KVl0uHeft9uhkI
1DO2eKLXldk/oiaHPpSa3nTui6p447yOFeHSt8PhtU+c3EMLAoO7hiEHa4Y2MRL3
TptfKpSjYiF3EHqRS5On7OmV8S8eTWIIZE+VuE4h9Tlms1MP1ki8884ogk+ZQ5xk
NjhiSWHSFY3zQzvcO+IYJPXwI1hkpSQ0PwnMjLYxHknqbvazfSrIV+K/IBQXgMh6
q5zKjK/c6xUbZrS2RH2UynzGvMJgvmMdjU6TCymOfiNvIfm7wefJiVN0gva+W6Jx
GIAuUPSGhQMf1pTc0hFsf08W6KydSXgQJtPv3tuzT13p3zDGWrQ6nvZx4h0rpOaW
yzqubzH65u62o3840pdVwdbCCDYaAaZVKb0raBPUZU4o+dweB4Xixcq9PHU3aaXp
Bfv2DGNbS4ZfZ9ltm24EGGeqNLy3pk6C1k2+A28yrRtIOahBO3Xmk/SBRcRdPH49
TSeN0cuv+Ano7QJWrU2wNlADb6yOdcmrUjEjMSEVJcgXRe20VtcaK43Ef4FCbo12
x1D2oovHXm1IZTUPuTJNsvkSX9aHXgblDZha8EMmyzxqIRQOgLWzYbsg8gAdP+dA
bz+XQpuZAbWSGBCXydCMvQItGQy1WsZdh5GfgAW1XslL3JxU1E7p/o9IHTToaWdu
lRggIS+XvGY8o884Y42G/+FxG/eeTYmRJRlg3nJbFjbrVEzb0796+UM8RFoRLsVX
JJJehOBxclWYIA9cyTxrS+Nh1Q6PkCVIL+E4bbfDG0Aokrv52vdiRaFVVwrvGv1w
oqNrPgpO8RY5HziQJf/zI5HdMJtP+Eqj42GwMPWlCH1DA8InZroHcvPTLVXt6lvD
ZkpvAYDCiZZvgXWROQ3aEJE7SOmdxRJNdrUxto/CB3ApnzpShgV/Eonqx8s9vpcv
O+sXVVdHf4cP+5h5VrMyuIJpI4J1h8/VIEmXJs1k4MBG0pDGQQQaMHT8KZze8tUU
w12a3Q5UTQDYcAohM/cCmulAZjfmnoNdX/PMzB45yNpeFMcid1cd1mijaU3av34X
ob+tABWJsSMP0mloAg0GXkP8PWG1z4LPooC3q8HV40qBFrfJMF1ldvyDiOBUtzps
HAPVlrbtauXDUR/fvm8IAUsELE7ziw2w6X7z9XFTTqyqZ14BRAz+JDs5voFWqoGs
WzcckfjeHprO3wBIrS/geQdQKkielFLAljQMNvFBI9S+naw4/g+c/+fhzc57LqnC
MzngqZkpipEJKoZmSMQMeFRIlTYqwGQ4IOtyDZ221S4MV+1XbenqLH+dQXYSVoMp
beEwp7d5rnzxqyovL9LnUInc617NGiYI4oo3SrD4SKex5kt98HAju9fcwxYn10wP
bIAPMBzz2CC5TK9cm/9oVA2P4/5rn3kwkjYNTqXL3+s6tJ2hvYzbz1AU50miV7XU
QDWHiD2vmk9rLB+GInikUh5B+0k2cjxlh4L/hIGO0Uawe7+V9tpBjmDgbUisiz9m
aLhGFJJho4cuu+uARC0zsCdfxn6CvrqlU0mWDQvyDiSGouU8j+V6O67QiC0IzHjD
r42fMJdFOujlsoLGk3sAzhkuUJlZGU1KApWUroOYJdSnJqMbNf5QmlH3fz9GF1oJ
gLnOYmY6y48x0eFoDwwZ5bjl968cGasyjm9xHhgYtdwEIoeqWFBWq6tuUC75/CqN
twdwCVi/jPKpwuNOiNjaX8m3IJQhvBTisJLb5NOu7fvn7+I6uVdSU0orYnlwISD2
XBjQeHpsWCghuCd/ObrZH0E1Lvqja5+ndisCq46Y4t0o8C3mACakkirgYsHtj6u4
BKvnloXHgeQO2B5NeOj9i2JD/TdEYcS5JWHiJ44TG+9Zr7HQgmv+AgC8IB+i7lQD
37bEgatbi+9Yt8rkTjlrA2PF4rJS3bbHcOdL/VGrxSxAyZN/Ma1lheVZ/K8Fzl/v
R+NA1dFEuEHSqwTzpE5Sjp8RJNBiaROrtTMfdxAy5lzfwpoUwG6+H/9FmnIbwSAB
Y9nE6n/CD9x8jWHkJjlPEDf3jS/4yUMLS5s76QaQl9P9HZcfpWtpIkCgLUflmtJ9
w/czNvVrbLjtb7lVBeHEBNxHb8t1nl7HcorkZCnVV18eY46qp246g5iGI7nrETPw
g9LqA7eQECtkDIcACiZeEmjsG5zNIAnYT5kbaurVkYCAac46ImFo6c3w393tgmvh
Yofz/mWsJJ478MFccEkZg8ukhAchc+LZ1rxIRm9maVVn3++MdHTBTpYo/kPyAadf
suYN60LSTuDJ+/xMGIyeW/v00Egt4n1IEiOee9R4otcvYyXmQwag163oMHVkMJMP
9q0GYHmR+1/bJt61qm1YCk5HB05a5CppEuq3ecQnGfX63qVBHDglCIJFaz2HuDqY
TmMgzP7ns9JdCUbZW8MzL3RbH4FhYSY8rJxceNvQyhfxtYhiE+D1Qm5P+aPpZDkS
qCVQdwWdP0Rp3Dvl8VqAeC+FcQ9leggNqkMTRXN9kq6FQ5nPOK0bI/HthRlpVbyY
vsnK+4bjoVibGZ4WbnisalAKcA3+3f97SYj2gefw/g4VIfCENQz9KAEDniuSg2l8
0DosJ+moMR3NHlEXsY1JbWZeWTeV8mn75vtCbJzJwQDMlu7Auy6OQnxB6Przi01E
7/ZmxniXj80VUVOvzjuUbcmSeGhA3jICPDxEyNL9y57y/Twaulira61o5KSj7cqi
6/mx0hJJSyX3J0ybvfqz0/6gv8MFRUhXW5ZFXAZixA32Vco6ABUO3CKWiEO7NxOO
/xSxtJdBdUy2tMyABcoGaRsj774uJ3Iz0LZg/D+A8861g48wOpEzERzxdKbZbHnt
LZUXfpVrR5LRokrB7eKxykydpbGcCpIdvUa/PLGWyYEosDyfoD+XdxEGx5DMyI5c
M3uXXDDif9nMxMm53aN1cnAYPbHi2BJKvZjJTK6Y9f7KsDgkqP1Qs8887j1Hlw6c
ne7yrRVNOtjlWZruTgaRDAyAdUohvS4r/9urdJGJz+yBtmm4Imq13OHt1MRXu0sc
e8owDuiCRR9rpwkSp5ykjAnFn/CdtivP1aB5FCjnLkAqiXVZvykfgJ1wYJZUzRCA
io2Qxxnm1La+Zf8xM4kOIlQE5CaRmwVtAMwOlMrDhVwbpZpzAqRY5Vz1Z5aIrnFj
ndhqgt/YSjlmcB+M4MVooU4Pxh3YRzEwFmnbM4lliVIIKUJ7GGYzWNSkHS84SM3o
n063q3t6WE2QjdQnewYZ2ytGrHgWGXOBIoc4+wHZlCE7HWucwkITHbC1Q1trKuhv
NxzkSRi7E5gswp3A1xviiVeBm8Qndx6xvSf8v6hhk6T9wrUhRxUAFIe8LP2RudSY
iegneFZDHqlsejpOchoKfn6BIp9uTk6dnZkvVAMItByHQH4u4+2Lpd6oq0/Qn+pe
CAyXqrYLXoEnXvn8HoPkISPO+zRpID5cneN5kXzmp6tuicSE1Mo58c09mcq7jiDK
1U/EtiXt/iMxNnB9DG6qwC9kyG1VugnAEA+lKOF0kR7y4TX6pUyTYD6Zt80s2ntr
8lTj4W7aHhBDxh+R+7VZezRBnjE1NtCYYTFFXiLnHoHfUMRGl6c3bpm5i4Q+1FuM
neyWBbVG/TSe4O8KMgheP66bmcnMQ4aE17YN7sO4RA6GMalzzeXQmPj3VizrDOuP
W5YPOIXHWzddfOs/M6zMn+Uih4OnEo9wo4u49K4k39FomTQ3Vl4pbhy+BeZ1X72U
lrIGIRcFWFaflP8BbNjv7KP7krLoBVR/lEQCHnC5ovUEc73pvj2lgRG+OvxXPg9A
nz9dTgnvIGHBD170ZQlHPzHsgw0gjxF8r3r3sJU1p98FMWky3kiemVm7L3nOgj8J
lLluXt6mZJdf1q8SVQJC88JEO38Cb0clNp6unwCjSy9IEHXuK6gLxTRU3sVHKYeg
ZiZHLNyFCNH7reBQA1URHWB25SjpJoCSGFuqbySTLtOvKwn3gAfMeoE29H1ZOc85
xmFy89iv9WbDlgHtWrQXmdAAdwESM2IJykaZZHhLhiZPUhMlS8XdQSrBGvnHWCYd
IIbGFxuffhNp/ctxbJT4j1IdmidMn2Y1tMfvYeLOOJR0VuelHFA9ECFxI3oGwAIh
WJePEssYtMPuDyeRYVDtHGoxLesM8D+a6YhlxZsTZklk+AraJNmfbYW3fR+JX1TI
RLzgNmc/LuO5wrMFHaL+tqKoYTN/ctC7e2OVPmjcp+hb/7pJRtHUEIz0BFW5nJ6S
c+pZdN4SPtBG3tUewtdIBNAX3UCnn62XIUZx9NxB3cuGERsSPcJbhFHQIvj13d/c
5Tq8ofN/P1JdK4eUUF0LdxeoMKR/fwPNzpb7n8tIa026ERbPPb4vLatqVN3CClD2
kqSitD8608pq9lhnOdE6IxIiZwlj73haaw4wHNZTyaSNBX53qblDfSnS3Zx3cPpw
gNR1juXSmvnotNMuEwcTk4eAvXYgoNDBPwy40jPxx/kaEZJKcvB6y3Z9YjUd/J1P
oixfC74XYiCVBPoF9c3HwRhlU+gWNVEWJXThQRTkGQ19z33AuT8BYqpPBQnkJUx2
VE3nSL+mDE6zE6raeUor0Nd2LOX3Rpjm8ZTPNZxS0XQy/dRHTsT1xFZt+/ET1sx7
kHaj+hVSrjxe/tiIKuEL48e6v3rYwfVJPlvsQVdRbG13D6epqfM4O3mJZhhVO1Ur
d/HoNYbuFYI+t2CSp+9kOpfYdWeYXMwYcSVhSmCXxKEDoZXrleCs4/uN6Zt/75J2
uTxo2gD7L0gxHHbzU7g28hZuloi3flGjPU7maEb6DH2gAfXuBp4NmxaTO+/3yFlv
Rzo096HXWND0140tW2RSc1rdMnTeRSBSvzIyk5u4XbHunQ6GoDG6goWNZWkgdKtR
MujyDQfAICz+ZIDtbHYI72hVzWWXFqqtmap0tW19p6pExBt3qhywh4LFr8TnRDP/
McpwT1msyv84UT52sJ9LmqcA/FiIq6Sg1op3wDIDltjLoO2QTKtP0fQDKnqPO8lf
Ja5EnLPtKQ6Tji752U2mEQqQ/82suUx8kBzYdWcdyoWvulFm+ujWzlpwmWSaf0N/
Bu41NDe8tv1Ck02kIGyVc6Fj7DgBf4os9RvgmdCzOkJGJuOqJAO0h8wuG7YsmsTa
V84BNTB9Idh51v/7C94KT+DpYQyyzqyozJXHNiMf8HuIyXmDy8zCSitBMiEMlfhq
uAcjZK0VsoxzG9gSu9xj5PPL+iSuk6uqm9Wc5BBGStjelrRR6kwSK6Gd0k5bHV4g
w3BGQufo+lreOZhjvetDC+yG3pqyg5il+vwxcFMAcjmFHSv9J6JkBOM3ZylCgrDw
4ulvSmwbADdKXoteR9/SDMx8ESkXeFBlHeIWqt0bR2lPU6tshttQZx1Wf7VxRF3c
Nc3itWN6wYsa5aP4beUfJooqyqpZV+GeaWieJH/k2IBZUyeE2f1EXjVrJIwPhKmX
Tha/2ZOJ7LGyxIUbP7BbMfqleVhrnAOQTjd1I72HfS27T7dqBGroQOsc6SD7i9oW
zCMdcJUMbHBQxz1jmYxuNvhuWUzBaARgwS0gHF6PRRm8tYjbwuywFI9GPLCeVFmo
30nwhoJkjBsdaKoQCgpuE8FYv4j1rSP89cH9d8YeyQxA55C2pUxtp/CWkfjy54le
/9ahiynZxxWSiT9K2ake4JH9DiyPrjVVBpc70KftTJqQdVJj5vZZH20AR9CTSKNd
LZRsV7GTm22YpZTcdn5AtWfTS0/lHhPYdVY44Bsim+Ai5KvvJSWF5/k5r4uUSpPr
MsVipcWa+SCMOPmtUIxWkYzfu3izuFhxKOp+aBqCcw3QmA25D5V/pyRbdguJkart
fHd0uBtRLZ7j5BW+otN4PSK3Vwawwjkdgi9P5kdO5SFwfMmKw33oF0WTGQN2INtf
bNZe5xEs3EbMnulCBvYUB19NIWhZZ9PbUbn+tTA6p/g2otUH1VfnJfoOieqM/ElO
yWOT0guPyEMFv96BV7m290CxEi95g2TKmisvnOBMa9h8t7T/+hh8GrdZhqI/UcTN
uSY6sTouEebJrZZvzRozgnDhBE9ievArSlT5ff4p50yznYXamDMMM2sAytqKc0mH
xEJDQJ4Yo+g0wPQO/+eb2K/9WWjvuW2oe8Iae/n68PYk5AOvJz6MEzZVxcxnbnym
bCDGOP3VwTiIxa+1TJZDEQduJswTG5ywdbtkofO1xcgVxNsiAbbxVOSmpjy+GF65
xK4PJGR16XgaG9vzH8VI6tR1+KEatWuW1vpu2JIWaU3L47O25QTuxB3KYBumq4Pg
IREA2UBraIf97SQzrLDmOaGGjgLrr+EsWF3L6VaHaUxceMMiTY3TCRgopIjwMDMF
3KP0ldKUtg7wDhAwUTw+MctgGFRyaOUzuo+LNMyogudiViBowzPHkeBk4ZBukEaz
RPzky90y9O7Cvd0i2JGlAvVUXwHhPoVLYfv2Igr2SFKeuuq22Ka/I5k1OePMSBpw
xgjq2vINM48mFxkGJfkwd/C4tKpi/rKSyos9nk14XHyvvLnFLVbTsFa3+MLCg/+P
J4A4Sv6NiS0ZZnB5DQFdQFRd3eIxCuZgxCzMJeHwcwCGmUXil4CnXo2NR1cF3fDx
nnMPO4mvbth6H/miaECjS2ysrgxK8QemK/lmdDUCP9zUARPn+UXfQaCRU2q2F99m
dkTAAi3qxjvk6DxX30dgrnGgis1Rz52pwlZaW6d/kdMnLgSejVlmPmUUh5kdR1HS
vFzrSa2GTcreYd6lEZQJKZxa2j4cA6LthAy3G5mDirCqqvGpNG+LLE1s63ke5TUx
+kUYtJvXtZ8+c+OBPpO77s6aDWTwgHm8US0YoLNEEpc/pJpYmBBO8iUP732qATzS
VMoQBzL4TwZzkcgdCjeC+N1Vnly+UcECzYb+wJJBKQ0C1K2teoBJ5KVARLl4xvmm
EUVknVMbul+vfSLKgj8et0vAqf3/kIg0KV1uGoCBYC0xLBxmtusPDbrPBbrKxq4J
m5COD+Ygt5MTS2nChwAJPjxg4LsUgxSYwLBXnhipnN+WV1USm2CLZ+EQIWfNz30m
VSW5eMbcXbN0cmhFFp9NZQHKEdzw3Ww4HVxPfbElGvA6KbDsbefod7SinVQY/5zF
B7iD5XFTPdCEvZkGMKwT0OEQeAbcwvsSAd0+010iSLKPxP3Y0tcY/d6Z5lnlTbWq
yynN/XRRB6es8dwLfN33eF1TZP23bLqx2I5zDKVdD7JE5QgzoXQFAYdqdoTGPIUv
2lfn3w54C1tZKT+6DcAYeeuKeC/RWwdGSAPa43SmzxSXqbeuFl5DF3mHAwbnbdQe
I1i+qUgCICNxg9DmFruA6JxjsthIqz7k32E5Wf54lZXir4UNp5yJ4/Xcq+rmDr/+
3jZ+RSy+sfKe9Myv1Cv7hrkzDYNv+Aw6Q4BH+xVJQKdBg7wDij38Pno+4Be+5ymo
j3W1RSrpzJd3p/KzbqAamurHk1/k4gRYB1wE/DON1xqr2EBDIwSdDGCORnLSq87i
TZPhc+ep3udqrx25/9MDyddI0jo3IAyIzcZZCvlY6tRbudmEAtowK98UySjU45BP
s4h5vZWthk+L4NOEDqjmwCizQpGD67CuoGSO0ACgriy3hChUAJ/e6TdvrJBDV1hw
SO+s7Skhh/rbdUgXKmw50U/JLPzTdnAvXRyLA319HvnaWyAwlYBg15pGHSBoMSd+
4j6xBEPD6XqErWbmwywQYKZw7y4KrJLJds6cVCuVKTD0XCEFnLO2G4jbQF+IAMCe
1VMePtSXUymDKCh8ax26uJRAMXhmcabSr8sGfgpr8LggTc0lzf2NmvOrpj6wJbSi
LxuOmINOjUyVWkNTPaVFAyPvf/zuFDvqoXMWbZq1Bue2MMzvkb0IkyQIPoAL+iAX
1KC2td0Aevg6IZt7IMnaqgIApSWK5xIWjm917K0cHkUEeF+TTevNmzy4fFzJUV6P
GxveZgqSJR8B7UGLh7tIAFjkowZ0eO1HKsDcLtUZ69a4CIoBngst2Mb5In6qE6HB
ep7hLPL9LbIBtOxLxqOHCqNX65dJ5UMxysb33ux+C2vmYs5Xrv71Q43EcwM9YaD/
vxr+un68yuVuCcvEdKnEf59SF3QFzCmhChi5qfLfKljQH0cvTHE7F4tycnsdzASk
L+jL0qNzXS0ttwxeB7NQdtZEhfJtSzeGu5i1QrTlj7s9R03mxKN6bv5oNsAS3vCb
7oT4xhB9rrkaUc5koyc6+40AsHNiLxSNx040izOU2ApblhTvmX7SNmGXKGb4bos3
wcKaoBuTjxiS/wsmGfmvhiGWGwqK7+N9vAcu/2hJMoRXed4bpDOjg8QT9JJdIm2F
OW33RDJiLK5wXzuoG0Mw0Y9aWBOL/1FIN+UcTlFl2qyfPdrR0J9ybyft1lrxvsWL
TkuoLLus0Iraa4Ti89XWHvRMhcCfXpmVZQiDU46wlnu5o5GpgjDP9E/CDnDThPky
oeQZv+foQM0+Q1KECpvVDmro6Jn4yInoMlXljr5iQ5S2L1a3z3Qd6Jst+7QRuUrT
B4O4J7Lt9Ut2QXgRq8/T7M0+HDA1EEveRgWYFXsWjEypJ3UgJRec8OkywxXcyLo4
5VvGUHkoBLFeDCxraQgWQcHxbF2gKI4N3jyKUzfk6YJ84gSkr3NBuapn+WX0yAmg
Z6sQ1ZpV/hGWKUFaWo6db1maf9EsrcJ3Lk1kc+mrWpYvdDWbf20OivufFpe6bF/L
vH63fKr8ESnz+gQ+0j7m9PB3rEmfdSJKnJ9rMc9Rvh6kuvITkl/TPe/7WTDXoCIZ
7AQTlJvxp2+vxGNuG4yEGBP5eYwOSYCQ6Jnebr2fTk0xBjUPPkUc3ZvKSqsvDkII
1AmPGiwgEspelGJlcIIcg1ULwh6iLCKCLlKIK1A+3t2eOQwVvqYsVuwXHQn5CNiN
793aLBpr7QuED79IPMCJ4IHcUzBgGuk2G/59arBqjPeV+y9u00oN378yVkXkEgIc
myGm/Lmshg2CFpXQmQ4rpgaTGKGB82miAuBiPThRQp7oJpSSW84Z9esdkUbODN5S
jQpaFByQ65+IkZIqOCQ3IG1oTJLhluUZTDhxyTTDqOAHvfIBDPPsuyuBnhm7fYt4
FtxDJLqG2rPW2C/MAwMJMvWgkZ7g+urcuPM1SLfmRzHHSxHQLzRnIHKRTolZB0bK
Nwf61uq4ciAsrYA9k55mo2xA8VB/xtrv9nsEIUGBVJ0f7N8bZZvBTd0beoZrbqj+
YINlASYl7DCUxYmjSKTV2MFUYkqNVVUVX6CgCO3BlPwsvD4RJZumlAXjb0XXcqIb
ZLsnwMREOen7HKupbIHSMSKEnNCxd9si5alllG4D3stGL3oXOmEAHDS2SGS99MQi
UTqTKHoJPqZa9WRqLIEng0PF18T3sBjksdoPQZ7Uhz4jIBCZUMdBIVWYC48X6rtQ
Ju1q4JhrMAP/OvGQX9SnuC7Ze9GqYoBw8xe61clVzCB+7t3yPzIdag4JX4uIS2SE
T7RaS6Ms/GhenjpBUnfO7vizyBEd+sti2I1wYd53yzx9WhbOF5HRPZGFGPx50yvW
frNJRsVdh8o0KdQUGIsmzSjYKHz3HpB4wBcqNusWcQr7LPcjicrPKNJ4oGWsdvrB
VmDGOgYLFASTkhGdbyStWVSgmNW4hkNnBaqoUVxR4XLo8X2Fq2ee0rmuEovr0Ahw
/gYgxY9Oj7JwUy3+aFNMgNAY0VP3kaqMznO7iCgIBebuWKS1u7gB+hH40nmSCDX6
4LPk2wNmpHg0P+ZYg+DWFsTO5Xz992dX0lVytZF0Y3gfPBwcYLiwkkDnwp5Zn46J
uNpDZ/pzgJcKKT55QIjSdsrkQNXGzH1jRIXIemLujUcl85Jb8aRH9Yk2cQv+FiWw
6Zf9WOdbUQIbEzqfTSqx0xcfBREfJVW+BXIhkJmALn2bpD78cwI3FVGni27g8hKH
eYv/G8OB+o8D3UD2YMD0k86FfGE+pTtiWQ77fBLwvjeV35dBlBfio4CNtMC9YZxl
4KRHhmcjSIFf/ezXOJ8mDRTNHKK91nHWoIYB5cyPZx3dADeS0WEhU/9aVYGkL3no
QTA+wwrVvazKhAQK8vZ+WcYhJ0XoyxE/xP+4UmednJp90ExOIKbZIM6kNeCSS9xW
Ue2rc8rs3pUWatmYfovf7jd9Mxq8ZovRUwwZPVrGCQGdaqif3xJ1YqaaFD8VkTzp
/qPx/tb2736MvCnULa+vI/9YAiLZDALG/rQRKDz+DRDqJZrHitxuj1wY2Ou4SrUN
u0vkh/LeaeSB1dq9cftZ53t9xgOLV9c6pf1bO/rykoDd+0kXcCMMQgxXa9aQHyVg
BmthcTlQr+t+lNDap5Mwk2mW9q2DqPwx1cjjz+5kGGQGC8Hh/6UfE9pMuTakXgSy
i67r8JMFWODEcp/EJrDSptYOs0UIJZ+76hCD7XwljeWCUwLyzmFEznEBAZOtOCwe
M+ejGaoLf7CYZL5xptUZnrmqRmBDmwcQSRAR8iXRH3WYgIJPRktq5x27A/Z9cgXj
7S6HS2EfuETFbtobRzpxz5CK4v/GNIXdP0skMC6SwV39toDmmu8ActkSdWTyh3or
GcD/g7KXMigNYaO6QeUUHA5EySWCJvU4M/ZS4Ss8KFuv4eGpZgC203OuqxwLf774
QeYMCSWh6k7UWir/5qJOX6fPTOeeQI4/F3Q/2DagF6LdEmGW/U7Y55OwG9Ek+0Iw
s6O4t5WlwBM6vK3r9Erc/uTTaJ776TXytTQxggZJkHD92VOeC0gqGWlz2KNOK5eE
iuQXbW6N4XKKMn27OVzIu5w7Z+feAEJmiL8PkAvnv9rfIUE6ns8GqaB0lwrpyKoZ
AjRLCVuOGU//GkKRLELdYWBgl3e/PCjN1AQFZBMvh0OOwCHR2OvwIbs3E7W1pELS
ujaaOmdssGRh4iTH6GWDxdJKVhv+pMYrmODC5kDGnKjIcll6DpIWxs9F11W46Sc/
76NoQnZqcc/TtoDnJbDo3zIxK6r8Jf1gyNMd0mLOsDLOwlU5xU1/hX6FTPOlMK7O
kM52C+Yhe8I9ATeG+90zT3Qsi3PC62YuW+DPwn5tiTbhnmVYaJPp1juPYIn9rRzF
pRw4pcNbAQiplRGFxuMZqriUE/qIVh1BGisF4VQSDbuTDQ0oO21niJZ/m8FDNOhL
2Jc2O3egKurQ+IzX0FV494pqg/7rQxogKMw2/N2OhADBFI2/8XXZapeGQy5z4Erv
+0AKOoayyP4c26fMMcD07W/Mbx1kqcdYHDAVuQkkodJeCzq5UdQMkUQQxJ2yrs2m
PPExu7JRiT64m1fi/qGOKNl009e6pfeyIsqLzMrlQn0gF6KcPUEiVt8hRfTBeOP9
hym4L/+b5dLv3K4JZLEqTfp0hA/b235eqiUKt+E2ftksl/D5PofnS3l4BsrME4PT
mr6YwvPMAqjPElsOEOPf60tXweUMj9USM9e/Ds7sEJlWEjRPv5QE1S/PR9PLVBiF
v/ei6KzBKJ1J3zfRxUYwzBBWr47CvLICsM9MJJTQKLos6WlhotKAz/dlCXOYvt4b
pjHo5ettDAdFeFCKwebfkAd6PNG5OozVddA6Hoona+2AS13oEvIue5OmZuQqzHf0
QPRgjm0/sDxxZwrspBIv0dpBGqz62QRwcvU0LqcoImRwaZWWqoIFONNQhN5ETPrz
DT2SWFtZqUrp2e26DEqp57mJwOJLnRJ7UjtXWBhlvJUHYlEn0w//lbotrPxMs/mn
pb2Y0hj6/1rnigJi2FOXmSYBy8PcVmLVEbLtlsiosP8PexIHe7gQyXUBdULrVNFl
BkaBHwlol/EVdi3mrRzTisQveUYixuuy7W6+0e9AjyZOL2pWeSZ39EAmiFt0o1Se
7+l62t9QT69osO9qXCoqHzHcMh+XPJM6G+bY2k9pjFhJZnU1tKtf0U3v+4k+nAVy
0MBB45EJUnEyHPseUcDSfbvBFG5rsW2GmsegXV6AUJ0N5rsmMzqulnoW/TBGZMGE
ACDPa8RJ9H7tjy7mftHEzMWW8uCc7JDpHpUlSARMqbA8HpRZ+dG4JpFIemjBzS54
WCzRZaKSUV4LfSFBKLNgTZFd9MHq+nYvfcg3/xHhxbpSGXOThVm30CoNyPzVtqVZ
S05TFnxjRK8GWl+dszMPn9/qS5mEgu+gLsSEMeFH+w4kaRkwFA3xNqx/uXLjF1yh
sql0+8Wa9iTULKIHlJyFWsBG8cyF+E2FKOIVXeMGNdgwxqMHdIAPOwHa/49bS6Gg
jCZHlYnitNrFq3mVWM0cb3hKJwpGyS2a7tONihbZ7PW+z7JcTy4T78iSwi93Aabc
tcJvOK+NLvnmVHx5Su3wFE9PS5ZyXcW6LbVNHGBXX6fshX5UcvsRIDC271omhsA3
YTFkPt8qRWnqRbhSuLat23by40gAKFQFCDOvu3lZ0uoMzrDlTmOoerTVriwj2wR4
L4cVyMHQ/jp0149iKek/itH6bn9HhJuaEpQKSzB38MpanNXp5LtC+3CGkLGfyTcG
2QcZ2ZxI5RPrXk/+q4kavAcn4b7XCOa6oec6Bmzbe8GGGSTkHMAC55SFy3txhIvW
yiF7crwMOZioRZyAJNuBrbt2Af0GjKTMMPAl+uuzeM6sYxiieJzCGmv+FQRaZM5h
Nu8DxzeqbqY0EKLePyYqVMk7cSKL6gCKgRQRYSUQIcBllTFZiRNJA5awI8kcu81z
tfk5HWNiQvHvb1z8ZzM9Umch7l+/CKTmhmHZm9kYNN1E+zT7qMiv27cU8P3hZ1wu
k4zC0FoucfUNrnkR0g1xsMZ0Yrvhqs7b88Tsoi4dazxOHJV0r2806anhg1KMlhcu
6+hwkYbhNDSsNU73Kh2jJ12jvuKykVRq+6pcBS7AtTL24zxrh0v0gGC9OtGVaDXV
j3cLPW3bVAPeGdp/YXp4mSwGPKqpWgvREz+OBuIz0lzZqkxn0hzXNtJLOHZC1rzI
xYVcsBhhsNOWpD0NJPigWvnxHEK7fuJdS9bRBIei5EUJ2BnVSkA4/QYmamiPTjzx
w/xxGaj8wASbNetmCMY0bprzJHfiVNQXMP4QPCtJdqH+hRdfnMn5YtV/Qv3QJRlm
KOvO9OtLhVuwhIjuI8qKrDsKlZ6B0ywHokbBoV0ZK8GlBJyTT6ASDAg3IlReuA+y
SJVtrscpvtqWdt9pUwlUtP1ZDW7l83wfe/+b2o1dREb7KO0P77vhC3hKK4Xr/2Sn
8RXnGfdniKbiEY8XGSW3BtEaySzD0vyyvlx4kMK5C9e+WkQJieI9k0zliB/qj0x9
OwODhuYLUy0sUtp/hxqOiTmFFnU8D9BHTcax2vSYr/RwgHVZXInSvEpBJ7uGRP3v
7vYH8tuXGwSgr6py/RgWY25eCHYuUD4ZPr6M5vgLgg4xoetOGVo1eq9CzYUcim33
b/zKcjF5Qjd0KO7ZRvCzfzyAuL1Gm5lYbir+pXLgAwCctVFqVq9FxKj8xCrhr3NJ
C8rvUfPo7nP5RL1ge9W8SWwpPQACtL6R0UYmckNwRL2fksb2ix8QO/0oqRuoPQLm
MM/5pY26Gr3zI3JVOpkgkKEBuTNXB9hzYhIqz36GHtCQX7ylMCHNEOmjZABo2/Re
5Kn8P7/iSk66AhHMhKPE0mCseBzjO2L6aEUBNiCMbekq9StHeWbjjk9I36akOYHL
/MRQHNeFikhwrMrqP9/iJV3Po0BiUd+Kl+8xpI4yWMw6/Vc+GTaQOZr8t7RlTrrM
gD3LsvbcZaKexPQCItMYoemMpqCGlGZE6esln2AVxGjpCGGfhtlrIk8ZkNvvhJr1
UvRjvXd4ih2GVTgON1vCuNRpvv3risWDTNNiyfoOutNJ87lXbomXN8tsmgJ0CG2t
2Au5rMPdL9p9ojXl71l697z9JwHrUqp+kbWTB1FqqpOSIL16A1Kp7E3anNNoHLEl
VoDc73/UkP9QJoOYdV87k260hMgiyxX9ee9ymSNANHTm0QJ5AlDsEIPbE0NYfOkT
l4BUIIhJGfvaE6V6Sux1sFwGxuxTJHtK6B/1cdWY6EE6RnD0Ydo+UdkWmTnZ2pQm
PMx8Zr6eSobiUcZjuYyo19WPZlx8AMRuJUkQdvR3Shlt2t/yjntyXKWzJZgLRkmI
HoaOHx3qIgnvivyGq5eXoJAuYPeC1flJ15NTwmgjDBJ3NCSOTmzGVL9spCGSEKhg
eGS8PbLBrqMwbV6pG27EFK8oDQHD7NeCqRhemXLjkNkPJX2abP8cdGrzA4iNpZD7
LWJqtbviNydcHrVrUM3CZXtgtAFV7Vhq9oKh3wMyBlDCdL2geLOpHITBqzQ3aaL1
963nY/Zs5Ldr5kDGSjxS/oNaWYQkYRyFVqUawOmHjF3E6qdLlbokzkExKKmZ5TgP
rqEzy6JBIGUPl1M6jMlPp1Y2x/syugofUakqmIaYleZBQOcnwIcN8ga/9NxWnbcH
5WUcQXAJlOjdiSWuE4h0KQ4S14C+HbuK13IVAPylwo5yCfiVOcPw5aHZuq6RzUef
DWEHqdlFEBrj/hJfRFeN+mUboa3PfEMP/RFTwZD5zSheUGpR5ethigro8xZLFuRz
akVhb4FYxm3TJ0+JD5Z1YRDvPE5Tdclzqto//Wt68AwDzqwS83L+hsILEO4aeeDg
3I9vr9F39raxsaO3jnfZU3u7mSuRAocmr0ntRPyHfPOYX32u3ABOXCRGpWZ+lzjU
4zDGBYA/AdqgfCHJOeFXzrK9P0hmSNl0l3q1yR5i1JQJowdjmCu9xY3YePCZH93b
aVTs1DCnGPrl6EP9eepP/Kj1EXksVjJuCInt8ldvAcC4Rw0FYp2Au3WtJFBXn+qa
rf7NDr7VA9nVrW40rtKbMpSag8JyLjiZQHa2EM/HeM/EQ+MDUjAT6Li26LMibiH0
WvvHRMyyMQZ7DsVH6uYx8y5avg29O3+3Mq7jxWqHBuWgocSjDizdxSV/h8inlG4y
1Gt92xOKzHvQ4rI4WTb0JHH1t0ZV8tzR5VST0GgOTzRp15CvzUt2L65tv4JXh5Jt
/bjTc07Jm7Rs/M8DeLFmv1DP//eVHUpINc6fTMXE/kSBQN2tzaTxCTSQy7r3QIkt
veiPSXtoRE4yWiveTt/3OMx4klsXw2wHjd8D+7d1zeRsdKrWUEBIxC2ZV8laduuA
iz2jVenKPpEZURtdVb1z3aJ0w3ap1mK8N5u2xqGJZhuTyc87ujV9rvVhS50uOCjX
zZ1wbqq5ATf4wpAViVCJCO59uxUdfqQMKosUTHDP6PnUWzistbgVIwRIsXDVzpik
+b8rEkZ3uCziU4v9XzJZpYAzMfdzwM6M8bNda5xvIH7R09FV4eI1b/fkN9q1waYf
ZUCFtYDeDBHEzhIkvAucToV7hzYQtpHdX1e5VtHSkZe3tcK8CQUW4Ht1CiiR2FO4
108ykTcQVPa+GUeiFn3CX1yPTuwySVIEV7cDw1twzcvWxte7UWkcrC2b8A7dF6Dv
M4yDqsZaromfBkTzjmJcYsZrPVg3UXAtQS7q9N8yPVgqdzC+IGk7so951aHNXc1Q
fZ3elBI6gjaS2GQ52HVbM7xBNpcpcOxxDtO7mdDtOGtdJRm9S0zI/LbX1OGbhz8I
w82wd4Ejgok78yCRDbjgQDD49BHRcBMDXkUyusz3CfWW6SYfi2V/UrGsAbPpZAkJ
lgU/SbqePMaGmCLQpGWMuZbuxqOWUGGcJXRnZr7E+oA8PJ37qefykCZ6vufJKcUZ
LEVcMrM2iORcQ+1xagjCcrPjuUq+Vbnd0WtYg7C8AuC9AgK6MLM81ABUjoYvIldp
aMw837iozyrB9S0HEt9/dscxbxx965XrVfuAyNWxc3FAs1A67lSy902c50eKVWWV
sMuxyiVBlrtPSrFXuQdfa1Yf9QT1j2fCw0myyraKzsE569ln13xoBTRN1MeZXbFt
HTdiQDsmhUwad5aYaX0iz0n2s/AtqBwwuDxxYRFN4YtFe09jpGqv5J0FEVAb25Wc
7oRooGt78frqKTSUTNkn64IzNjo1A5ZuEB7wKdg7mZHsBfrHRbfY4C6dXuGsjyR6
Dv6Cbss1gHqqfqCkEa4qyn0+E6hTHKpUI+RVi5tDl9gn79/Xq7boA1LvlWcX3qYE
4WmAxeijo4m7sgykSaU0IoOdOlOyZTLGZQ+MCEfVHpSOdE+SzEI8GW5TDfGUqSVA
4NFGXwH/9V7zTh348V9ZlsAVLpguR3XDk/OTM2xcVrGopKEtbag1M7N64Ji6BCoP
RCoJ/sI7DViakl+zw47kByM54YygAcp7FlM5k9O0ughw6OC4W0aZyoGfRi+NymRA
4527sLijINpCVvuDl8sqZQ4VSbUn3JSQcEUhxL2lzldI/kTvXhUznjIVZK6ZLnKp
FizYMo1F9iskmV8wOe80FNK3Mtz3iKaR1hs7qhS5DG+YC2pWNjS5JlFZyQkm0w68
+Ov4eb7YencbUA+eBlG6YPl5d7XoIqazhrconAHu3vkeipGv0+H+a0AEh0GwRIGB
tiVrxv3o+qqzIWy+sbOeSpEtn0Ws5/bpLn1V952NBTeRUIramEYE+dOjr/LlNm/C
D/Om0expdm9r/HPpUCLM7USDAl2+5Mu1oeZQSp5uDnSJSv/SOPIJtrPHtJ5mzppT
8sOk0BYxc8oYeXzfUxxdE1uOVk9io/GKVUG4RUCjsaz8SJwF5UFT0hL/vhgKa6SD
Ln7ff8Jgl5KKxiS18k2KqkgeRTQztJ4Psc5MMLrbzDHpw8lh+jS1RuIagfttXPv/
X40Cys4h3SVG3+xfLoXYgVRWqtEsYjFTpdjC5nFB72xSWY3XYSirwjOLtSKQQMxz
HOroPfESGynRwcFZAPTqmvK1s+LFTrjVIx3I4oq1O9O8+1u3UEYuwub1my+svN5z
ZNuIMu3mGVAIndOZuu78mZ8Whb1ySbCNjkdIETATejZYpEhTT3nkwOwJhCa2xGEg
Hf/gYLxKtMb5LZ5zbOXxDOeRMZakYA/k3c8bPRJMpjInJPYS8uiWXxrFD0YKW9nK
9rV7/58GEFQQFw/qU8jCSrx35uBqTd0652rcK7TdgW4O/xCMSrmSQNbQorvDm13Y
tswaVqFtUzAXk30/TD9zYUztfgmZJy+7KktUHt0DXQ4+SgRraXhCeaM8AU+M6g7x
hki34ACxbZYgG+ezMTepJ4cI9Iq3KTmqZHQMspLtgShcA+AjibN2GQtq2HaJWPV2
66luz3JaQ/30enCYE5QF79CzTSBB9kPlcdX8ZuoD27Q+jkcP3UHE1ziqmmCWFdck
X+FqwxYQHqJ+TLVWEKB/0LQD8WYJWRgnTP+OAK9eQuFhYi+7WAD797UZvHwJLPX1
CtvTphUFkmrb6VkbBpqBf40+V5kuxnaRYIKcSnc7QKdplrqE2DBRiQCMkes9yDCx
JSgD20AvpNs1ZG0ooBi8rvjcNa7ax0QcipFpdWzEac90BvB7nqvo2KHpDRffvX5B
SZ6UwrFXeGK1Kf5dzozTNZdn0cUTGoMAPOyBhkpzYkXVZOTDr+wjqUkQT37a5aXV
pI/uqiGrwswDspASxuBIQDq9/o1R1w5IaYN/LWG27mEkZZc8xS0hXpKXsMhHErhC
snuwNdxbu21pQt/nsvXTeyqXEe1R8rFXYQex6bz+rH8jsz92QNzt+eYFUmvaRrXG
k090far/dnbnT6zFOUZebsotHvAL4KWFM10+kA6FkZu14y87WckXe66n8pccLJ+6
72PgJCjROo5707wB1w6+EnLRwPHQaNcynFma0hxqKh+R6yVRTbgWWPPryCMkekol
oxYZunsHS8sCdpJoBohHZHvd/Ul/vkbJAe6rwn7nUPF8wEUifk93SzDJGzfrjWEg
NttTsXhg0zTsceMDjSpj0t4vny0oIa0bzRysAAaWD4ERSHxg/zST43cEf3myeVyQ
gWN+I6yPhMppjX26IDKAuqwV/NmtyfBR+jUx4p8ey8wQVPUoVpkfj9pcf++BSppz
a7dk4lMf1DdS3p/kyjYD5kCaHmxN0/WMR+RghLfwoZq2yE+CnJAnk4XG3RCp0bOE
w0kjBrk2T2SKgxihnwg1TyJ5jOVmFEiCjpBTEypXRdsZ5CZN1onGWYAZXXdSmvX0
DJYQwF96oa/HuF1CDHQ6rQXvWle8/d04f0ltGvxS1EMyb8bUsbKPuS55EjAxdz+z
P8widYZq/SDIsNOmMi0sLvQUe0Oq6Ydj4wSwS8wjQ9JDvpLLcc8kIHAG4MbDbId0
v+CnOawd7VvfeFexHLhkX7W6BUIRFyoQ0tP9AEDcUZz9dHE6FEVsOIwn5368SkUH
fPnNOngZo25X57wAW4l5mvPm1RLBrILyrdfpDrgKeRkz6CQfu43Z0PCjocI0Paey
j/up01v/o7uyD+wU44wge92sM63hYN7GLyzIsSE/7SW+6sW4RkMdnXSeJKgUzNd+
rvZZ/AEvyJAWtTLHNxVypSOf/puTQGLAr2HEDbM06sIiUELsTHVhTXbNRGinHXMk
XfZJVupBGV6Z2ddGFH/r5zCK0hWEv9tg4dA5M9212pc9VcsWaBjtZHWDZiwapfYT
MK4mO6KDA6AncMfvEGGDvH7QY4Xj1/pf/xW1NGJsSKltG+FOQHsqktyXud6yEipF
x16UhGBiImSlBlhDWJKx4J52D9/p/PCMGNIvzpCnujCTA+ry499We1ZkTVpon52K
eQat0FZ+/hOHTE97XBNrczwY3FVuatGd7a8trihuISXDVQ18lNLwerr/molT/Fky
TYEXjUW+8fPbkMOI6+U2tBkRYu2qPoV8CU09wpoJ/0rz3KdN4p05Bh7Atbge968B
zTquU6SSvE4jeHG6W+gZDgJtRLy2fuo/HvWq9nUTvrxSwklwLfXZu+7d0bE1oVU3
T061Eiptp4wOueKMuZuwDmnL59wFp7lMr76gyUP7qdzGrnsSBaY9YrIfYJ5mKUfP
gIMgBzrIJYziJCPv+cheV5qH2LBiKT7WRsfrwBG2Zz1kt9E7nFSTzYAd25OTWBbY
CLvPH3YsfxgVvsa0QvG3WFEq71zfgcG17OYw2zUsFETtRACVymME4j7eIDkCZrYR
mhOgEnBvKi2jaokVMURaw5KDgURzrHKLuhVdFvMp0q4xTDnKT+y4lyDWXHNSZX/V
fyiTka6UhLBYxzaHKaTm5O4gsHSsUtXS4tIHDJPJX4LHYsr1TbjXmc9TawhXLE/A
Bx35X+vPmI7nhNW8nJyvFJbnvwAZmCla/wa0vVnVFwPuvvf2vmHhL/O0sAz5+CC3
mAM17sNj2LkQEA3/Lh5yZ70+5oBBRKu03C/FrHDW0nMoH09J8B2lXdgZjQQCBGNt
ScDzQOvXDqFNdNidkSo6+ct3K33xAL5hBU+/h2pXZgMULhIebxFjHPU4cJZKmHvJ
dWHQbL83WfibHOBMNEAKwpWsyEHyr9RHVPKOu+SJRE9DgSa628+avd4rFYslIbY8
1R6xmpE9UAydg7Au+MweE+Vfuc3HZ4b5z/a32/xW/vyoqSlPIc2r19B/X9fbbeso
BRxuXDZV2nNGF6g1nqbgbGuUzQKIwrq40XoARRfy6ljP960i0wLUoIukYYcvkrQ9
4WanMYXZtn2ZtJr3ve12DQ+WIg3Z4YcUQHoYf5fpyJMU+wi+JzQFcMo+U5xxILLv
EimEvhA4m6fUBMVZrCF+40H7bp0Pkm8ILd4SY0kt8fr/tPNLa1YmoZu2r4axx8Pg
cnFKGBRNKFqUN/FSgE00XxGrnKWXNtv9S+sccwFfF0JYDPhvPGXbzf+NTgwKFEkR
AEaTiA38UgNGychNoa8pH9v7x0qbwXbp2EuuYpcuRTFDpnjaZA4twEYKdMvYmvoI
9vvfRoPH+dEUN4zQMHKfakdYy1yz/D+D8OySfaxotaBmwIaSlsk1JQ16D/R80mUP
rKcQhlnq5V9wQBjSNTbd6nga5IsHAUWb+s2WiZx6RQCplasy6SNh+QAPP8zaeqD/
eeU0AY1olpzCWfZ7044jHBQEUUE0Uh49CfVNV9Y4NOTBOi1YCnQ6TwP1TrMpCLSz
noBhhXcDF5waYjioPVtinZBErOzj6/0xrS1lUJAom9iw5nkgGLTOzzRlyFe2Xu16
xKPxZZll2CxHhlKsgLY7kLdR9FO7DwbqWS/C/vCa/Zyf2dewgFzsCuQY8RFot860
buOEk1IMPqi6p4dEgb3u64GJMOpbScFTDIiSmbVxYHJepjOJFqjdB6Rv61MfU4H7
yWzjQvxBeQb4BucS0Lh5ySUZxjpZ0AXloNH/anZJUTyeCDkRaYojH30+7XzMkNqM
W0UggBWbfTMCBTZ/XcvzBY9QuQBujzJgLNmlbeGdcmEkFBIpC6XS4l+uftLSamZ0
5CybDObCMsJMWTosfIoKSxjafXloqwPl01RRUbVj8wCDBN08ZYMj97BHDbeRo5sj
hRtpZBrODg/VRpUnLituK8Y/+KFCbfIPwAy+Zmphwk8/rXEwouv2BP1q2Z8e5USN
ojB9mADcUCscHG2x6Ohqehm3/ZXWTg0EnR70C7dLxn5d0XQev9IMKqG/uXhUirvU
bnmdrf+L+EvhjRgqnh6jJ7YIXOPhL0JyfgBQbyWA8gEd9LMnNxcHn7cChUKAqqtR
cneXDVM8eu5n8eY9YvmxkkrBDB8fSye8HYp1RTM92qVtdZoYLr9QUV4gR4Q1tGzJ
OTdOvuAT6zWAQvP/3xAGe5UdpzlBlupp39xT5SHxbsolKZr+8RljDtyjWwaO6KCq
eqvzR7mSIJzBFsx8yWWlMWwK/6u2D1Ebjc7yNa90KqJ21QX18yUA9cP8+pgsTKJW
0DqoZ7AiUuj/GXbMZ2ril1ssJtuALyYQS+2LiMZqrGxOSNgodBCbqzZCxdIN9Y1X
mdX3lFDIbLPV570Tff28akE/Cp+9VTevR4kwLT2EpSPSrOOzbUJU8rwLbof9kLOi
mrKFUcd1AcJiGdaYrq7ucYp1PTAAEBaMx3EOX7+hH4azWQqzYDhirfFF7J1+FTGB
Ts9M2OJ8lMC1POlpAbEsY0xZ1OYCJtMFKAT7D3gZHhrjFWWTW4Wu/sX/i9M5Ag3c
a4140YZW8MSLMnx3UHa8b+/4JUaW8NQ8HJWl8jzUZfTOQNDgDj+QbcCorvYE0OZ8
fTuI1Ql22n7OrrBvQ9jX983XnaYd5n09iQMhjvF0MGDKZ0XZUzQXJi5uvDxPOrQw
M7/JcTepGEVcdpoa7wHmqL72bUvNfGHYLYk75WLiHMxp8tzY6hsJ8PLz9CUUJrLO
e1KDF9J8jnsdkn2eAfDYPjTCbjiehQjrYB8iDQFKnkx8Tm45aBoKScleDpfv/s0G
pYfx/6Q261w45ejBDRQQuYngl4Ci5K0oQN0Ia5G8xNkYGDKZUC17bNzxdO44LQ0t
jfO7pQnAjkcMhxmFx7z/EQNmEPYav1bKQZwpV0Oqwv9E02XRZbTb7oK3QgmI7r/e
+hGsVZdrnpMuZxu8ypdisX9o3Kh864oPQxEcbiCEXFu/A/5NUfH0tybZ+CaKw6R0
C8eNXAs/+JLBY36szv51Qw6cTmoBPVkx3Z8NQesq9m6HKmcT/5tXSwerTh2DutW1
6v01xakL2gQhlf7urk5qwYP7SWQOfVy913/aLx9a36WqjH43TBbEjniouJVIjmWc
0VloZqxuxv4KjORSYP4CGoS2kyyYlfdbXR80oSjj4NY0ZeVeodw2GX6dZbxUqdPy
zzjQYR+l7nKZEsw5+lE/YYEhuUrgj5a9QxKKifwnDP4BToXeKRi9ut+ulFKf70gj
xc7WHI5Ynxey6bclx/YMNuGJrKxvPi3HT4Y0nAh2w3t8XKaRqmWPZFVwlUEqFdEv
eG+9MDRGuhBMNm+Ylv8/ZYXEeWPWwM4a/TlJKeOMGUYrWU052udGp34dU+2FqnzD
KSy2WnIHoSCWjZMNDpLxWPIcbBMia7KlaT4tdTVIIOTYPWImZSygQpXg0TArQoDG
pWbRXcKUvJYGZTdOJpM2ZkFOzhE+WptmQWgjl6vmhDoqWx7e/5EbxsPtT2+JfYoo
uxNPZ0KEnCtzEyfhiOGuV704x3CXYFIwNAfZdij8gwIZF8VrqcwAHPfkoNGUHI7q
nN6OwGe5CJQK8RQx1uJwZ7rhMu6oCNhZCVaiq1TD51Ht9CXUIfImADOKlfqqFSdX
6a5j48nCEkCKfaf0+VnY7ZjE5x2lbfFLaGdOqXTDU3WNfV8OdTcEpNvSZtvsRqqw
b+6580ekxoAqqMJiPNX1djxOEUePQedxVAHC9tmX9RdHs9rgjxv9ZMRo3gGb+muq
Y02ZHzmQnTeruR22N3l55ilRSYbMJEECUxX7s4ZtFSMBXxslNBpgHHYOFjfMpwI3
6gTpsZioUhWLUxUEu1VrqdxHExaVEP3CtaNe4d1P7tlri2b2qP26jRmBj2IqsFfN
OJkhEbqp4DuVBYicgLYpmPrc7YbddeSFkYZf4GhUg6z/0p0EbITiuM8hVzZx26Kq
YWW0CRcCcr6f0oxxA32PWZrxGPXqTHOxkx6MzyQx55mNKK1vJ8SWt0wnlLq2xVcy
MTMy1Yb6QHuzVfVbK1jfiYLdVpvSbgcanEt2IES7+to79iUIcoA3a4lkGa4QCRn7
MtKjsU+5N87HLiHFhSvti5T4IWaqpEA3ozyrpykRkpltx3+e1OBSYaTssEdVvCqz
RndvrYGUizbnAGmy+YKvzAWR1VqRboFue64gkaI444yldk3JyAcr2sjCPIFcA1jP
gC6x9E0h5Tfv+K0ecKqwT+se+YXY4b0o2oN2mVQ4+Ok0aiqAv1Nk0Xw2Mkyu0ryo
h0p/Nj+uaVZqRs3wEK5zaChicV2B0KG7VJD41rI0SRQDSsNB48pm2jg6aq2J/ZkL
X5jwtuSaVC5YI7PjXM1P/lE7SzPIpXFTIYt5LJmxzzh8fL2QLV2cpo79x/VxGRh7
nirIiWR1dU1Xf/A0u67JOsAOgw7TAFJF7y6QXH1/I/G3eggn38CxYVBkCAR59Nb7
0Im2y2vsPRyW/SWNbJd2QLulP7fGihr24gpSMACqhWTnKKo8OEldLCOOf7MBv3J6
nJ9jy7hyB72O1Wjx2XOq06dzHnPi5V5fmZ4U0dottRbHv4oZUxwVPXXbzzOzBFGG
TzWQPEJFcj0in9TJycf/QbyRW/tHgrTdwKBKqpjMrrefUPIRFsGg2JohIN/a1GxO
1yxPfG9U1ZD8e2HoCfj6jrG10H1dEhpGJURyB/pOgSt7VU73CMmUTSTB/hl7Tikn
yCRVvXm9ol6Z4lU0ji+HQ/6irtH9sBK9yydMQBc0FwsLl0lJo/Lsyeg2VbOQNZzq
qWFm/sAb9M7eoMjzLnpw0YPNEasrfYnl2GEnO0iXav3laiqK7L/bSlDqWqIHidYd
6R81P7icuM0J5yLAHoLFBt3xx3/9FLlv69HQbAWSHOLns6ne0341rDrGUdWvIsHc
jXYVNVBvDszIGZUT2VAUbBjv7nC+kQbphcVZjn1ySjGFzRJBd0mealPK+fGbelhb
VHRlaclgY/DP5NSXBK1tZzXOJM8IyDiBGn2Alszl9byTX7Q2/Bna4SMRd6mzwQFy
pWLp+yc4VU4+qaHcIzsw+8Vj4dRMXm5ZGEEIi6EPJ0QJTyW0rANH+i2Iyk4pB/gp
XnPUwIvkFYTeDfZg+Xtbq5U43jQUS+tN1hzzIC7N6rPCtByY//LGu9lKmOE5Yop+
AxZisqoLTEdOSBVI0UkVI68SSU8EnZOoEeIrpdFyVobfYaUHql7bx5Iv/k/1LVc0
1VJhAWYC42SE5zpXSlxN8JzoPDtXPm++XRi+gPbuGX9VKUQx+sqcTfcne+s4YTbl
8f8+c0HaJTsGI6MT/Cxc+DIUToSRAM6/zW+BzEwulFfmr6/9mKL7iyNd3yKU3ooq
GT5dHjipVBNxCam4gz7PbpuBSNGXSQMRE5GKdTBlrOKCfU31V+aNJUiaKlFDpTlu
qqlSwQcMdexmN7633ui8rczg2Zp6do3OhuWEJHxmYBQEdCYXTPVqI62b8djZf0O6
tkXH3PlLezYM52gTAANsEmKl3dsncxRLE/w5UJV/9ojh8GPlTzp+T+a8xnavOs7+
/RWmi8gWhtAvUetYZ6+BUGNEk87n6+4f2Ia9Kr+ibBNPMgATIHAc7G1GMZbtImZD
P1IqgAZ7pDnBGo6L9kNnUOv+XQgQYXYzmoj5ciwl4MDAafO7IvxsXY1cXFTMLFEg
lpHYNBWdhw76776+I2GxdNx6P+O9uvrU7tS7GXcA6TVwD2XX8HWp+W9FJ0a6apg6
/9YqHDlu1rTDcto/zwT+YQxH7JtajIeJpKl8z1V1PN/hD4UCAM0Nl0YWdJe7t0Dc
mtXDnDgcV+tJoSw/x36Kv9wDGyRpllr2lgzxOeQKnslETedGo/mBh68XPeE0hPOE
/Tbah+KH6Gqd3REwDsygv5kp0rnac99u/g4kjDNC5nahEVsyni/WkRAuF73vOPqY
Uf+UL8lTPiAe+MkWEVY+8oezIK25BkIULCjYknVIrAWwpuTpJuKOZ7uUd/XrZPyO
F69wMOU2Bs45wcZtKgSk6ftFZe2pT3tInx0kPz3spURsM1xhKHJSmMFyZ8fYZcrR
POuKBdyjHlw7leF/RO+R24tCKd2xaaJbG1FdLkpCTLnGUQxHQlLOzuuxJNRjqPQv
MIp09AEMBVbYi/otOX+Kujc02WZ24m793PXACAAgyj23Iwuvr3QJcYuIqpz6mghK
7z93k9Qr5oYQWQAzWdyoRg9y2msoziY7nqtCpMLVWljlsxAvrNKzlVSyT3j+kLlC
WRkO0jgaVWMHZ0pxotftUWEeWnX0wmQbiTwhj9JrDIevAwwfCWQYlkgAvGMbQlXX
Yx5E9xQRYz0kePwIUp3lQJrlLFwL8oacyG8LFTPGXNLcQikfStXu+gftrq+9pgup
TnbtlJ1MFbzBXjA8cV995TyYD0g8tMR34J9duwteP/LXgubhi91FY8NSlMb4ouNp
vi3h4XDiyFhWPsNoPVpgIUnwlix6V0Y2z5P59M5ILETn0c5D8PqdFst35+OYYpiO
z4mU3RSNjAw7b84znaCXsmmmoX/TlgMHXw7WhCzK2SNRbk/Qb3xnGffxO5BSH3dV
zQDRELRzpmUKwzhoHFyoOARL70d1XZNs1LxkgMH1jmPf5lmlmA2P05c8T+Qgjcq2
ihiIXVH/6IV/f3u1ytG3P1oTRSgspmrqvSzYeeMXmYGmRmrGEHwwZYQjQ0XkYbSs
qGsMr/WCq3nkYKLsn+o8zvjnSIO2WgEmpxowYighMppvzrLU43AiiC7IKUR1JmCU
6nU9TalV7lp1Zq4s3HNLIBfkk7XFDfrZ8d4yPB1eXIouNWTqmZwRLxIUqzefEzaF
+jJvCmzlo6Zv/ejt7OsgJBrr0uaQXzFh8ye1cBcRcgWNFIDknMKEhlkebhYW8Zdf
wBs/Gx7BCRQjd2Qqae5gL/Dap8alPEHnYSK1npWJNMrpryEj6kMpJ3G1mrfsyNpG
BD87lSvy+rteCY/XMqEFEfMSTuNsirr1rJMSwILlM7fh416GZbGXQipOoK7LbTVK
RPwYPNq3vdu5uH6uSfRvWX7zteueLnkagfBp07XRXmbhQ+URSD5307lO/Q5NlF26
bx/9nJH91Z8EM7XySpTNzWcyzmtPt6TbnwgVea7D8xOao/V8VcvkvCzBslVNS+e5
yc2tWMZZWZ9ch5RWOKrh+QTGABCSZK9UvcWkmXUTA2BylQOG0cvEYB+nSvYyRZVy
d8Ml5sBdctXtriw+lHwf/h4jvXcx0rUXnr7gyiQ6GuBpZ4jUL/Je5y5diApdQ3v4
oOuS5l2P6Z7sFfCDbqZx7nEEPIdb9rQh7Ks2Y5klREID9qjQ7vkpZ3uAS+vbst+b
rfpmvXZfa1BoIjCBSAAU54ddZ6XpE++yVGFtNObSQy7MejIzURK5Hd7N8CTEGDj6
K/qR+12s7Z2DKNDNkyZ9c+vhOALjtVgEN8lQHvmYsKRAzJfmnWOeUay3+ZMuHrLL
dAunCsjU/R0x3I/kCDctKnM5QPCW8bA0bS9QJFOXYy1eH3WpArHH3H5aMpchOPam
iYzhbD0aEpRgLQSuz9Z7Z5yXNeAr+Lx7dgJrgQWzM68ZbnhPGM9p1s72tmwIyynL
rm9T8QYaVmjjxffsLi9ctd2nQYQWqA5BN0X1gbdEXdimnyUJi/Do4el/HXwDhrHA
0zIV8sv5dRIePUQfrbuUZWk0fvlSBiZe+BCZ2Q3PuWNiyVwzDwRukeQCZdKxfFYN
gjEtJeELq4f4DRMCZsyLm9EZGgt+KM1sKVr7iXmbv5RJU7+ucU5CeqhwS5WyWBEr
oduQ0PHGD+zcQUyg2Rm4o7Df3OM1c9dmCSU3q4zaODNxrdpF4D/kzCJtOhqgh4P+
cxj5NP1t0TvhwzKqQR9BWlBAbBJLuk+ai0nNlcY74yjTbim/fnR2gJ+sKN/h4y7T
/4H9Wk0vgT4726W2p6zL7ExKYOWmO0zZ655aqOTRMdJLswRBT5pIPOWPGCQjP7VU
t83I+nn2Gf9r+W0GNYyOACTIs6Y2FgT31PTKtszzOjuUTJSnkNWL1zLmNuGihS2v
mLlk1T1NhBLQS2GwRbHO/y42uDbzU0ewCUHuuXWVTrTxUuHJRSbHSF0gMKtbfwAy
Y/THnsWjBsKHkWq89KT9Yn1AHqk++aTLTvaSWMyj/gz/1kX3mhFDOdhujtlxs/Cb
3oYpqNz7I/1J9IxZ8zE9Hq4dXHhSA0a5ONiUbhkuV5lMBxlCDlyuEAbX4pGCVVYp
Hv3MHDLO041ugM8YIjSFM2jbgSlmAN+ahyLzdIRstL/kRAzEPkC3QeEBEpV11J2X
p46t46EsyaS/Kr/dgzyF1VZ5oswlORa2xZ3mTVkbvvjmBI7V491siL2JWQHk1nfs
vqxYoOwNAkvVW8RTENwimPehGqMCxq2jL+aBRfBUmPd+a2/UuXffPEbcLYcL0hKS
Sk0HyswAhnYjOONafUENiqP9qh6mBRsLbbNsVT7O1EQZ87JOyg9v/fAGPeFpDlfy
o0AezGVH2cEiuyrNe3qaqSdlXU9T5UdmSYN+6VLI/k1TXa+8Pv5sc+Xn7VRWz585
2amVLxst3DcqGgDYJjt2rl/Bji4Gu8L0fwcER/YiHQ+SxX6T23lxT+gVb5jFivbw
EtuQ33aY8kulPumNBu3Ye4I/UOHtTVATi3ERHmsv+MMQh4H9iRDgvUmtRNX9hRWU
g0oXjpEWkHg/FSa46HcDZl0ZsBSqB/IYSnbbqHMvScJUsOPoQ06/eUyWeFIVbmX6
ssiuU0ltQMlR+d27OqRqcoWJwuBygPkKQaPdYC8YceUizbnIP9BYS8/GBT4weI4P
LMIj3gjb4WrBnpJ9cWpacu+hPG+SvA96yYSQb10fEQCif+/F38iTokfCHZRT62Qo
s+gTMibA8LFSB7xopvlJFBC2xObb37yzCikOy+kBkriB9oGm9/NY+IqSnIrd3H1O
gCmCNrwTu/KmyXzkqTukzL1CpLweD2vyboqb7H4XrC35iEkwX2ZVeIqJjkw9R6JB
KWZInIYz5abvZ6+Dg4fq/t6o0G/cX8XKnb4ycyDIGRjTz5YEqmryGEaNQa+dGa7k
AUj7N6lXUoBWAB9Ngt9KEpkd28G88SFOzVbCkyRbRxhiaeFcK8h2Oat0yHl5cJ/y
rFQijaDIn38v3bp4l26Lef6lVAKNQqsuvmpLdsNyO5azYK94rxfJoDmstAw/SJDd
bp2yZkRxt8IWNhvnJVQGkCqSU5/K6Gd6NnXty0SeMXwG9CvRPSKXxZJlzDcoeN1T
yB400vceqJQiVimz5O+FaG/NXX23UQPhXoIYqjWwAdTAvYeNIAkEWvM/qMc02ibu
snciWmTPBfR7zr62DP27ygEWL6VhqSYNGG5DknbHJlmkAkdQiivcpH8/Ge0FAiHt
czjqx+6m6MiuoNmsizx1R5V1kGvMU7qFTTAiJxVniyoG94iJLc9Cbi8+zVJk35OP
Y7rdjoManB0b9ub9GymEaW/Wi9XMqoWQdTeTJ/ul3pkAyqCIZ2j1qv7slyEMeJQ5
UkyhCrbLmFoSHLYxVx3OxhQAcpNgy1Oe4mBLoEQX5lhY5DH5MjLU/8So6fUh/gFK
dpR1yWw1uxcmChefsx6DsUDdTgwH31mfG4qLqMamcgO80LTaYT0Yzo7nwe2LW8B8
xZ26yMooEuayandDOC37bQU7zm4hzRs8gTqVrwMVTBAv1/z9Ik6aN7tbywB+YcG/
Nt4sz87s0Xfdn82GM+CM0i3I7MOdUsg1YM7SK2hJQUg7gUxmvSXQnAQueRyo2zsX
dMy6kYWfcEUe0//F9CnGZ78qi7uwokrNW2kK46myxIrEJireitBzOpmjY6QL2KDy
CiHWtauAQiltanJLdHzN2D+mQmCF5NkLU5PBhDYQmNNkoFIpMp/C9DsM/+GZzfMM
71ZRG49YmcvZdZwWlA1iYd+hIb+ZCUT6IdyT0Dr4MjxDKyJHwHoLV0KY/ayoRbKp
RIfqwJ1iYQJKBZAL/Ge4xJPzrNaKH0i2dmQCQ4KL6Z2xWPrwc8TELq2ZlzXclGiI
6k69/n/UdjUTIvCcZws8/Md/mJ6p0HSOa4XWy8Nyd2uXWcXTj+fI7SO5yTQSuHIo
7xZNFXjoUYPxdihxaR57VbareFcECyJFqF1bLccegdRt78Zg3+wyvKNfwhCHt+vm
LmMGFXXW+mfnWdcj39a/QQrbdWd588vjY0noJiZL0XwDo6YsQ4tzTM5iAU/ewE6d
6SF99N507C1hbuK3v9lAswX5EatDlCVY1Nl2M45PL0eR1oL2QZQNNAwhLclLEtGq
SGekQy6w3ymM1XviA/dlEi8i1JhUv5bYf98zhfyzevDNzFuWUaQlvOnxP/WbdGyq
8t3MhHwhU4kvHRKAv2e4Z8enmBKYjhSratyfSDZkn69nCY0KX6TvrQwbKNnAp6aX
/XGyb57t3CPS4xUQof9EK89REqxhuJnr+YeqY6LfgAKZXUUhdDfDXGz+bHEomDbD
eFfoY9ney010SMOErmrCqQ8NjUK+Sk33gOXMCTPlZJaWOLi80OOWCStR4jspS4XA
p7iLQKKJR+NmTaCguGKtA7A+DCDpAM908RZ7rs+Z6Q0ylNVUXRUWBaEUltj1HuDV
xCiPjGuvd+7SMf3x4kHd7kFoTOLuxBA9fb/dGk6JPGwAxWaGo3AyONDPRJ24DcHk
EN08gMQwvlKX3Yx+lUeEbWxHErJ2c3HrqetPf++TOt29Vpbcp894qaekQMgD4Sz+
varDDiRPnDewPBSzxoCsz6LBEMIf0XO4VPBhiW/4+FjUABFwl78klNL8muWV6QSI
LMI10ONRkrQDktPi7o4aYPiJ5trUV/juCmOKjnp9CURQqgj6JY2vmUM22AI5XMO5
80YqVD4sJWfOfrj8b/VT14Rs3K/PZy6H64f5kPWnaHt4HVM8wy2y9IhYqnxD3Dd1
JZZM9f7fP5knyIPD9qCJe6WX+HO3QJwbxFn3KW3mcszmxu8leQNQegGimhhClZJO
M+YHawzBVssIsKomaUStnKzZo/RVcuHJqRjNqPa855TbGAtN5N48SYckVsqGqUFS
h58rCCDE5mdLeSoVOCqeqk7gSgY5qbrPtlBno57N1szEfwaq+WRG2vQ0VoO+3m66
UWUNiF94exdsbVk7KQETDzc+kBQ0adN8mZDC5Au1coSvdfjLotYAfXJX/bHECU9p
aFHWZ++bd1ckJMj6MPEytDmbF8Je2ZFthg8+9CEjsaC0taztvB5SMmXkN8XgV99L
Zepv+7MIiPT9hu2UzEr9S2fbi7KSExBTfY6HnVT1LAFpC9iaYPSz8fJqodQ81NPc
cHXUc6YeIKZHp1lMEvF++jZhKJZTH9MBRGIvCFgkle5XzTnyw1RvjY35DyMyuvIp
5d0w6TU0O0TzEkX0x7+nw/O19OzcTbIomN7imvaIRdLjr14KWbsOoOOksG3tU/Ku
/xY64LWIAHLyqCfplNj5GtM+jkmAvJkZ273EERm3wRBkU9ExFM1jceBKimD/XFFU
QIw3uOTCS9xa7MN49IPpylBD1k6z8uad4yAvAnbqLjC6zfdp3X2Wd7e3n4JAvPDr
2zbmqpVmvCAV1Q4TKDApSkWee1cFHCuz6DjHhea6fd2NpiXmVZ3j4bxMuZaHtlzv
Kn7wAsI258WoauayfbepadHWCv+9TW2FDkQSRtRZ3WvZbH27hixPKiUQh1w/m2g4
V5TKbQdCv6ttvQHBE1cQG7XmMw9dvbQEB7/a/5913b3W79p4F0rR6Opk6N8MgdAE
x4hs4Ku1GtRUDXifv9TaS0MKbZr0N0p5xXrZXyPcqRo1nf+iyHLbEL5QSCqM/WSm
NxC7TGfnz4RN2d9RAFzDfsw/L/sRiDOUy33nlh1C5UOjka3WbpzWIVrf4AJIq1uY
zybfqLOeHEVtUArv0ce+Ad54zNucWK02JyXZVWS6sf6FTYo0YBewhTUy5u4Mq84C
8UXHlXqGYCdCLZsGKbtcohFKC5edUXf7blQyoGCPfPqJXUzFeGG0OSH76rpqNNNR
zQBY1r/eiI8AYMYsIbZ8rhu2cDJO1cM50O9bYmW5UlT+25p6UaRD3XphPOhAQpuk
B13D0W/qmlEvorKVwnKhRb7uv+TlJdnp5p4vqmGmjMEDJlb43apGL13bMPuST/tJ
TfoH9h1Dm/7rpkcwNYOLdjuRz5y2p0bLl4yTq5d4LicZnm225c5JRaQuqcLqaDcF
55fg8YaeazWjp9s8OfZPkmxAuk6hihfKeV7+4hXgKGxgimYVR09OqsEmOfPk23OM
l9BkX101+tkWMSFLX4jp7ahzajcPYafmt0tZ5uqTAOFe+d/YhZ7VNIEhUp4vedPu
qhkOQW2xyytuvtKZuHG3Maegth0BsMLq2ZP8jsRywoN6LmraTFE3Bbdbn6++2zn5
kBOKk0WiZSI00Ma6AWFjSNWY9mTj+D+2rDlzlEtgMIaaWhNIvFOqA22HGAL0MJiF
PkHQ3Mq5CIAjrfHuilYNqtRrxBDWWpYZT/5BxdcjxWNiRRuWTCtfItiwJdqOKoSN
YPAoDAsGVx3XBa5hdHdutBNoQXqdfL2Y+sEtdUgKUo1H6NwOV6yj9GH/xWeJN83A
JXRC/4XlsdMVckDgktmO1M3Cz0mlbpJY75JCxHWMEJ06ztU+vVNhFCTC00kptZ9i
cWapdJUhT2SWh0uoc7k6VnDKGIfO9LHHS8BJaV66SHrieJn6z7M07gpgWTnhupW5
y1U4NeAbldBUckdKu4n9uoysBM6gN1WcPnJuWwlndVGMtY3N/YDgf7Cvt1iIMrkh
WBMqqJkx9Ch+cs8VsllzixeBTfkdnUFCGBqfNAckJ+K+bIqDwoTFU1AMsjcfF4Kv
Hpsk1GX+dXeyi0VUu3sccv5inEp+a1UoCE1TltW3wnjA/GSSHHv0BcJFdCRrZ0vg
Ixxyte0Z3dn1SWy8iroHvn2o6yGd6eGZ1jWKjJeXqk2A/i0Rve8sCrKdGTesBh0R
8zGu9pzceYZdRb+eJlAAjG/i7ACE/1VXlylxAa01vZSCVdoncKwCpQFuPDUKKf4p
paVdXpvIa8Xp9bMaP4P2gMHPqNN6FVeAYScInhBqEqAKViegReywgZFAE0tF/cW3
ZW/NizNTIGsDvDfvMqe9uQ0aoUTwjQeZZnMdubATm+QIHfe4nP+MUqe/1ryXyPCt
i8hiYnC4PPbapwqQDNknXmL/7UwPUVddWDXjUzK81qtUcNFwduMFgPwMBmPe9Rnd
jgv7PahWzPuoFLgsOCa8X5LJE3YsumUpWCRSOZDcvp5xmaND+1cVKOuGBjvmzdqG
IbSXrdeIkh5XKw8ZXCxqjnh06gajUX00DQuWqTYwXxH7B9gQlIls5op3FqyDFlm6
cT6ajUgLELsHv1/I/CsIXVGq7bWAQsItinxMi7cReGLIcq5IGGHo7HdgQHHWwn1J
OwTDCwnFCwF56DBw7jUtO9Cty8BZidyNF+FgFtm++wcGptPWTyiHN34+ud7O9rcX
qQTtG+V1vM1kNGgQommEZ5B0BT0Cs7YAV4F05qnr0iHnm8374SN9i84c1lI+ARam
aITMGM+vI+9ti0G/X8xr42dwm0WazbCof1jCpEvlbYYjZw5+saGaeBQMKgviqweS
JG5x5VNGEYw73JKHbDcVYtM5avgBCKtkJIUxzht3qqw+ZgJ5pPdtNOQKsRbfan2I
p8MKaqbQ0UOpDsRcGClnt5BgjxNCvGhsCTchTW2+F5FQ+ueFfbJiyOGl7lbAjCSl
VG8/8mJuE3jz14aFbTnjnmBeqJgMs+Iyi4BrFhLP5S2F9g4s3ziVE2s/pFbETBV6
kt1WTDv02w3+kgtFnWWFiesLNo5I9iPfbseQLZXAX44GWkZfq2XGNn1yBl/jgdRK
T7JXpdLuJURlvKZun/IWR3q8t1R0VgEenk5TMPoQUXJHRS71A8fm+EZFRjoeQkWs
k5xetlE+yuIdEw+se+Vj9ku+Xd8JpNkEWZVZecNEbcMrwOgyqv1nA8jB7uqLrrUb
EHrWe/NX0+Hiy4M3/P0v7xepZXTROPI/alDXtW4aUjxe+ogsf/Ofr+ljSfZUO//D
NpWYOmSo9pPbwwo5K0/thgyP9IrVMd+yJRbUq7VaiaUQg7Pe8nD6UJjApb26HZNj
xNt5IJrnG37pSZyemXgTQZBUbC+vusj1BISP73EPSShdIaXH83Z4RuxrXMtbh72L
oMTKVGKKyLT1ZEDiNauCv65UEBEuZgiNLg7ZqFUjqMQbXi0UuCUo9Q+nNoVvRqH6
0D0jFKuMv6+TjMr0wucrSh2Nvm2+fyl4sIRAvgiQql03Ru5Y0z0E2i1bkdkTHFh9
gaFWCChWf9DRKzXvPF5plMT5oDq74cyddeUCOn+u7V/D7M5jPiRfzqcL/v3h9iWa
anypyXIyWAjqLlyY+yCwnLn3tp7YrVMK0wXPvvVpuaQREeVNd/S3c6mLo+O2yR0R
YVEXjjW2aKmuWBoOSIP6CnGMW/UlDllGhHMsG5nIfMDNHBpk5mCuCPWKjsrq+Vps
tdHseKfHPgahkFnMYFfNsXWF6BGMQg7r3K5gmWY2bQTmV1qXA3cKHEpRxkW4fl/v
PjRBJVziLcTJnTw8xGc7HJCKrPrHi5K5n/CIcBIrgu5GiCrNPut+Yr4FgdAXEqAM
l8oGZPlOjPg0bQJw2mxAaRMH7NcnPD7RGs1zk2bOhCYmUCPFyv5HRnp3GPrQJr3T
YC98dH3NZMlOyEx//Y7LeNgTt69OiTVHIzKzNy+ADprTUn69CDY5roifmdigi/Vh
Snj77inMjdkwJAaHyQQEaZ4lAxP+C4lcSpXcIFcyJ0kfGnFpRv3FIb2AjFbJPzTr
PdkPOWYROUL7GrXJn9+gQNs2yc/N4+UNMmwraJJxBbveZ+4CsrdSKlRL0/fP5uGM
tHdim3MTaCkoQnUl8q8BMJMrnd/8rlKuksGReLXgaZE9fkqoZOi/EVN/woIs3Luv
oSzXxqLkBJABhwrNVIL1LLAERqqCkIIkGhYcHHqO6uUFZtAcZsD6e6G+4XMnbRzv
eNpcB02rhszbVC/5X267svgbi7ERvkRLzBdab5ieBKZvEY9AyaI2oxnPcE5jIzDm
/Pmv1dgsck24KIufC6NxoPw571v38F8Sn6DPcV07dzQKm0hwNzmw7+ks57DixK11
ffPbZNNScRCGuWvBxOQSpROuONhxHzeWeXnUxmlzTvar1LcM8p0Bbe28CT4ue08J
YX1rxNxGXbfyvH16/yvOoLRlVRHKYhoaPHz5cjuy53ynfZhqRD6IfVNtg2xg6BjW
HrhcfwThb+kw9ka+ikajD44dvs3wvEgokSO7MZD9/GpA17OEB5mbIK9zX0Vpuha/
HpE0PmLwZBQZUxNCyMpgUfk/mpNkQYNR2M1Xu1pPcEezxsBu3FyI10L/iy25ulTF
B4bmNtxo/sFm8w3x2Z6x2kkZz+tU+Q2OX9dgTTOy0Y1hUmH8sWTuwd8CJpIP3J23
InOYlqu0yvXFAhmVJat+A8JhzDkrYDN01SaXEQL1NScsM3HWbDpxYuV+MM5mVA5V
7kf5aittB4guWJG5wdtjjH971YAers1JCGi5oBN6PWnnUaDfGJiuxjS+qGq4+twp
zzrEpFqQhTfGMiAgzyvLoC80Buz7av5kIJZsq1Qros8iRWDJ1tkNkJWYV0hs9E7B
N5MiR44cMbUBXXuKbGR00qhisswIxpGhz7s7U33C7sJxbe7CoDp+ruOY/7wSq+tV
+e0p/dK/vwZSHChNSExw+y8qKNYf4dvrYFXySiBpVPZffG2qgITL5Olr/ie48oJQ
uQV8EE0kuUQTYrZkz6ZpXtcHKtywoeMerzrMz83tiaJzeR4kBsuhinmQ+zF/MLZu
S0aTdAN+rSW7V0Js4Q/5xC11O889PCpeatz9COqdMcuHEXuyXncEZLs17hlSFN5z
++sS98Ms5sC13N7/8lcBrOufRqA8D5O2aoV0GzBpsSgMvWhJGLcX3EJk7fF/PoBM
sthOe/c/gvqorcD7kkA5LSP6PKtWeX6QKo3dffhvwyt58QIkwXCf9yl3eVm3ucCa
2ACRqwsWmjGkSw6qUDdkoDHR6aT5ok5rHPF8ZlTD4H6WPxN6WSWzKK3UyY1z1jvO
Wu6CcEy2r/9c/1chhnq080Wk+lmNQwlQZExKq/KCAtniGrq9MGW2ShDnGGJMbD+g
LD1D7Tgcxg/4e+bNnkKbLY7tEFAH8fKGPqkWdPgiz5DuFY/A1Nj2IsRTeARhdB3V
Y/DKqDAeswTymAR1qNiGv962vPwpZM4Zuwm3tfCpGiIiSgg5o9tmp+OsS2p0iXgD
wEq3sG8z3xWJUkARcuQKaFUJvyL5Fp8C+xdYZvxM79FIBZKV+SeYHNEj9IYbyvu+
m9x8N/Qs7ymUynCsBKy9NNAgUDy3CHJbCEEJTNrICPif3f4VSJZ0e8jLOIA1mIoe
gCxaExxAGM9yLudSN3BDzO0QnX7P/LZjZFt04AEM1hvFqSy5u2EHWtz76Mrm28hc
9fYE9ot4MqkdJRK8ZAJoH7Yeuoa2hnEiZky0IBKNx+toJzLFK8i1r1wfXRwF2vNI
ZvYrT+ESlH3W1SdNcQ5xKrDp2jRTqDY0Rnw/HXhE1K/cNlDQoicYhWCPdMP96Atm
ZxW+dOroKQzVESqooT2BxNqoiN2Hljh2EpwtdfHdRD0HtNm/594690sFL4ljd0up
vDcmIwRWS0S80EHBL1L7E6aO1WC8Rg4mhSa6Xcafx8uw5otSC0mvaG2p2zeOK/B4
cSVh7vkLwi5XfpXMr48qpD8mdwxNfJPJWmFbKmOeiQFheNdfF+1ituGtb5tkm0K8
dljJMXsF6TKJ+m8zWBlczEK/A9T7ltxwyuURsNUTuy2LugQt49Ynk8Q6QpOoW6Jg
it0fDVw5Zrak0FMro5uu+0gpdiQ5WT5aHdTapq6u4a92Jd9qKcSAL0D7kWUltuTi
QRArTscBkKnzPKEbRDrZXKn+NMgN32MgkC2ySMv+NF90zjR88SX2dApsYxxF51Yu
KnHGjVU9SkarFxpzyAgi+RlVmQUBy7jQRaP2cBcYwrAYEkwbmBO/Xi03FP6ZQQak
UncJDBUrpvwhsAxJ+geRDEDVY5ZZnA7sq2RkUMuf6NA5Pba2nf+E7IyQr61v2EiA
hWAaE8qYAzxUgS+g+l/SCEu1aEhdeRX9CvkbCVArDyebr62BPF+QWxaQ8M0HFhup
A96PQ9pCxdm5/HbEVhI19tAwiMp6dtj4bNA8WyyXaE9+ZdYNKQeEWPs6fG8l8YO/
OwXllteI2V87nDJjvSfBSc2HIK5r6c7MGzufeI2mlLDmueilLP3n1O3rH/L7h2VJ
WTO3ojb9fquoQjIm+Ifi4pvzXePE98nz+20mkk8Gm5JOvpb+nbCKFH/XZS4EPMYg
pqh094dVnHp5mcX4w9LyeK3iEKxdnvVYo8mhPm9/r6Kx3Y++vKqyJk0p58iL2bSg
p3b8fBBnqUmpLAIlq26YyTS88bsYMM//WOrd8J+XY6gdBc8/Jl986mDsWoKuSBUz
mLVB7gBBeRYl0WPpsW4mXqx/sc3otHezMMMl4G/0pzQKOYWYppVnNrQxdSH+fQzL
qVoiLNhIWIm0Pxm0HmgVC3mINnIsS4ZvPZSTiaZNs+l5xZs/l5rmkl6xN/SiWzld
xxHg6OcSc/I1y7Jqg3P+lgiBiSTk3aZ/hRnZmmmMiDw6iJeV93/lLv3K/hvf0dVl
NH4sv0+WST1nHx2IoRbfnUyx0UuSWbJmSSpnKImUbBrfpv5DDnkTK4m0YSjX0WCd
UeY76aNK44C31KvQcSwuFuH/nuBJQ6aL/h5IZ1mQ1GM2KnX7ONCErNUVxich2c3d
m1nFY+9a/GjB6FtPtaZYDIh5FICd+QlcGIXhXXwe5Va4Na3eGLAiYHa52Rq+O0qf
s2IqFHJRY7WmLN0P/rxT0ugBIFEzQ7OLgOa8j6lFt4cxq8vhxAxI5YmOPDtO79od
Hki8fsNJPOtH9CqG125CqKrzeZvB/FMe688JhEcfs5QIKA//c/tdq8PI9zFgsPEW
j2n6ppQV6FbnSCvTBtqvkCgGD2ShS19UVXxh774xs+n0pjno8mB1f3GqMBF83+TW
itut0h9H1VHCt2Jr0TpfR1KpUS6AFLXcwtpHgkSuvtSH/cWb1B5u4mtWK2cY1CAj
12TBsCejKezw1tr9aeSaMXH/23a+Q+vl6+HLo1+tzmWcl4B8kWyzeUoj6K0blj5K
nRCtYZOoOIZhbJAxZX5BApqhvfv45z6f9Dz8NNm+MifwcdDxMGcRVEygjruxxy1t
QsYl+NMSj86tYzRqUnvk2LA6G6Q524C9h7bd29UGonfo9ywps55/waRS8KH91/zX
n2ZEJpuPAaOTLG6wT/qo3sO7HWJF3bnVoRTLzeFQuiOYVhiZtzp59Utoy8TeFiWD
RmtNVYNXujlqaqQs4TiXPOVZprle3PLbgCU+uzWjS3tHOq6HHNWVpKuByVz1YNc3
H9qLrhDEd9YTnCew+/z1K7SsodVRNYlX9505DpBzlR0Ozqr9B9hPeU7x4zWdvQ+L
lxyMxYUzxkJYdxC2l0joh/WmyVXInGTxpUDTlscbvsEac8qPf6Stukp3tUn8rf5A
vVPrwYTcngsD8quJoXy3L3y6KcODw7BhzJTPGLm23zbBYILvpbtjhh+NRvjoMlZ0
WkrAXg7Zry04v3m8jloN1sBA9JuifV0p1WqI7IgOzSSl/NE1o5yiKxUIfa/xlnrm
LC3xcMUdH1K5KqiY7kwg6K7tAMSm07Yfp1LnOU6LMYDyj9a1uVB1sjCSQD/zPxoj
F2fAuFXMVeHSeKwXatnI3eo5MEeeUR39dqxJNhvlJqmL6nIDLTQ18TsyDck6Re8C
ZEsQESGpCXTBTX3QMS6QmPC7n+irTRkBH2Vc1jrIYH4so5Zk11S+bEe/rgG9DmvQ
byMtPDvqogvR7FrM+8wQAoon7SBs75HDUcON0+8qUVrS+ckDxTYeAJp0zNjK09nQ
gIOMF+0RnZAGjTuUiw7MPgbsNzUM6GvCpWP84pn25vJnJ+IM/FfTAG3UzcebYSyw
q9eLxBnfXsya2A+KSD22adSxfYu5VeX62uRukrk/xHdosTdgyghzXE4aaT3IvDN/
OBh41aWIjmqVSLTyJmWoKaQkCI/8n5aSKmULks4OHXTWYD/ecXOqQdr42hTEa+qs
pyqJmSguTaGPerbmL70GwpdS4W7JHzov5FSTgOFzWM8Z2GtwZoy8oTtQWZXcAQUp
+j1+00mLfiioFiiTecUCV8y4etanDWKK+Ixvn3KgNKR7DcYtq2QEd98lZVqQ6uSV
5b72Eo65uftHwj1Xq2u6zLsX8jgeWpupLdLaiEuz/+q6W+FdSpkVg1wrrV6I3mRK
zCDB+xlIgzqi2bvawgnPO3AMp4WDp9sG8UMZvOD5pPtvNnJv+EjuYb34U66sisqU
aLEq1F9yR8uaK1W+i1dvtsfhDojlzFHDFhnNPLTbCsneOvlmik0J5srt9/0rTzII
FpX2cVwzd2NNkDBPe0m7GYzVL/XILcTH7cr12QDPusV714SEGBFneObPT7SAmUJ/
zcP6ocZewrdVW12hegcLs0mANiGZxLriivvkJ4/OczITWAJtZo2iPgpnrUcnozNG
jmX1bQIKpcXink1WDJFqjjm5VYwspY4TasDktZ22YFGbdZDYjs5AlZPcWul11q/1
jEylIFmNfSRPF/BKQO3zc+NE+isRd7vNWmczSGavZffM+krYHYCPcpI/OHmcdKun
3lq4cTas7PPKe+TvrboLcM+dfDzDrbrJgVpaq21SkzGBlyo46yNO6ZzZSVatO0tN
iNCWoQ+OF71MYoTQzMRqmQqpO3RJ1t7fpsfiYDkxoa50fKWU0yR0tRq0KgILX4Fv
PWOFp0kXGWfnqOLRvKtS9ZQR+t3tRtCjdaWpy26J0n+l/H7RPTD1b33hwIu3JACF
x73c33eejOvMZEGvdKwEuhT32EGwR4XGEq4cSL3wBA68e0tHpqO+YgT4fPc+bD7U
X6pj45drBsEurKe2E1CXMAsOfpZlewgMJOBL1EeW4ZK6k2DDFSHjZBCzJBiMHlr8
yZ7hL2dtS7On4cuxHIVpM6WD36szBZDIP8Tj8jPMUWqvE4VAQee1K8Q02vMR4ant
VuQVE8K95vECuuiTbLlvLcWjFgZ/Pfvyj9khII22bUeSCfTnHyAuB6dscyTjJ/YF
fkqJ8Tw/74GBBWfcZg4evgN0cLlB4E/Cl8bg9wkvz19yX/RCBEVooUV3UvFXIkaL
veoTQR/MAgBQJpcwIsyRY2hOYg7+aPpC3NFsIV62QzlpzfvFSUa8DQuL12d1BJse
ugc+Ni19vBtZm0JE5qoSKklSv1/HbWM0gOWTLAtJzIuZu6RIhWLR59EIMWUl3Nkw
T3fKhHyAq9x55qJxBi90vbxeEzjewToupmXm68t9d+dqWZRUlbfmC4ykQo/DJdfY
VQZVU01YIJhzwCA05xGiEDala7+3msPwfLfZPk3tCNN+GacuODPWhAy+s/wPzQue
TKeLAFfPzU411cDBHs0ZHmsezMboxkr/gpN2o7XRvRnexTAlrJ6JYFBu1MazfdF7
lLnRTSOQs66LnF9igEmw66caaDucDTe1EW4esn1ruqDQ4+dcyQlb2HjGmrPYgGLA
ke84Wd/HQaVFbKJ+GApFSgDAyQIo7SnTNXHbgXc7pj5ikk22yoOk7jkUHhmnEC0j
aDjWoe+I/Y5ei5zOJI1P2K03Pl2rXOm5KPQ9BRY2grmbSXzsqHDRI3yqzOgVQyG7
A4h4ThOqDoXCK4c449ZUTntTp68dMX/AZcXIO1PSUkAjFDg8Yx22JO2mEQQdOywc
aMh810kyD9xYNACBFN65f9lmiSJVmutxozoz86swfDWEMUTtEfiCZKJWirdGHsey
BL/K0G6LdZ66xIWPYsB/IYZaKzqsE2Bdcd39yOh86CmRJ8og6ra7HwD0UzB+uxzs
X3kIvFyXxgDuvveDaCA53FTYSlnEY6TDVyTIYXc9kLNSo8LedDG6OxhhUyo5qXAY
8m9K8TfI3ZG/PIFkmhHwVRFC0jLZKxQ4TL0hlwJ0eUj3dDf1XQqNLN3MME2ChmJl
c5i3YytmbJgEyQWInEStOmA6LZpd1o1spZPtWnONeVszeAUB/tpOjYws7mm/D2bk
u/z/b6iSV78lllmDhigF1NpRMuuweCYseWXvoAjDbSltQOpzys3zDXx3k8yNIblo
cXCDTbZQCelLxCsmR73eYG5GJP+m9QY3jjTEr1V7k9A+93Wo42TPa8iSuIe5PgiS
ZCgBXe42z0AIUwuv5KS6oBf/Cd9NMclK/668/WbizYGSPAeq1IoJlSVt1YTuP5rj
Jgwv63piUg2URkrQzwURQGbxBgjK2PiaYtUlR82S+x/AFtBAX6AABvG/GrjERNhg
zz1eaJCklH3FWucSK9/3whAbGh+MYKj4y3xgxDwsBK1A2/WbR6EhAaKYpZ9OyBK+
xwy30JFI23RSgt2CuLoVpWH6r3of29SzdZtKIj4mp1ch54bOBHrPCAnQArDM8aBM
cP2qBtofyQZR7ogwC4+cxi8hoAZV0oa9W9VW/ix8PZsd7i1BEj/Tz/ss6NOWc1Qt
IGFdI3/m2qp+TGlgZ7nYXgox2uMOJBMRBeo7Xz+DtmrDAJS5sexo7zCMvDOlsr01
hcpprdysdnmUhkcjNPeVFUYKxsVZkinAlQT2g1sjqYc9J0CwWPLuR7TO8VY4k+0Z
0d4x4jtmIA5r2t9GMttTF2uADQ4vHJ0E53KgAymQz2Dpg1R2wePPvrE7QYbe4AGL
dezfnw6vuVQnFBqY1oezdnkEKCTgOpObLVQ7UIk0FFrUX1W/KGIoy/FMp6OFO8tG
gtsCoamnUbxzjFpoxKA6vN0Q3596ZhcNmois/KW6tvxRr+8qhApulxpdsxmwNQEE
64T9QX8fuM4MnZRNfU53e+5msD1xc/oxxtsdEl0fOePyXoqFLHSB/Y1XC9T2AAfs
z4Q/Y0NrEb530w65Ns0AZoA762QvbiusKoQLXaolirSOJcjbrIXD1D8AFGwfDZvt
RH46mpJTs/ch5DSDXfmYgxvTJ8nF4afdsv9rVOsmKl5zzCs234RkvWID0yraSzb5
Fg/PR2sRVVXcqvPvHDUk2WcOMDH9E+FTUGYWjizOhwuceImIsu0cQ8VF14qkTBk2
hPKDTRpSdgtw2j4PLgJUMNOxCFwBkFGnyztPNnkmM2+oO9xm7Z8b05vd6i+oGlmG
sJP1i6udIpe4Ln29km2jIshiZ4+gmhXoMMjav2z3sKDKrQPfAxMTYlKJT5Mkuzp3
gtolRlKV/5bnUWUDNBsNnroRTk6iziNpO9uRdoEtmABH/C8eu3nXPSFuM9oJMlnb
9E0A1lIHxZEES6TWMH0F82o5+4mEW09qfgon0/MsX+P++8nl7uHfgACJE4oi2FNT
EVoUx91FgrEXctaso4KuaOUDDppjkgzjjEm4psS70kolGdQGxa8an1Vo3UDH0ZJQ
435V6pYUVtM/WRZs0KtioZbeUb8Xx6AC6v3Fvd+iX7Vrlf4knV6ipTc1HOt6eEYQ
xVDdXmflhh5vJ0aV9qKHU1ItF3rqnd2gkQJyfy+8kdOrQJlN/fGMbA9K/oBsvltW
O5h1DzCE8Hx2+5etJrtnU7X7Y+cZdORzs/aZfyhKymIMQvoOMUmoPiO/oIypRq+L
RpqbQJiKcFlt5GmFAsSfsJY+Cu1DORJm4koCX7JhKNcWAuURRr0i8NMGHwNTcAKV
tjwgzq/egTO0a1H4Vz93Q0t0YpSkVdiN+fV9ySrKFfDoV4aeFCd6Ncbvhdg4JFxa
zrwCzgQ9ZIffE54VTUufK+tzPouNESiNyg8Dbazh+mcMUUJ3yIsl/p7Ia76psacg
kTYO9J5IkPomKy7U8qnPZ4lcetlFAGVdKbeCQc2CxiTdzcv2eGB6EtdgTiulEjlO
JIwiEyXPrTyEi3fLh/Nts070M19guFmK1zMFFMvvkMYXJ+TUMXzodDmmMAe9nxFF
tfqn3i3/Cjq+C9ge7H7awwmDWONlCWhMotKL6YckNZmCfFFfhbVRUJSokafK/LZh
fy35tNNwk9N1EAWQestceINAuNq+eT93lNtmomSNPg/orLsyLb02pCxbldgmj1sZ
K4GRm3dUMR/Bj6d3zKta3wPaaIv3ciXJXG/c5reYmI1+Sz3yDW9LdQ1t2qOdcYlj
oEhBX0GTI0BIDE1UCdHAWxVpQVRtoPrOmjIzyf9UJ8U5k+cfoo32n6RTxIab0nVp
5dadJhBdRhBcsQPq6f1hNEubpwud488BIVUK8g6Q88AR09pCf6ZxRmJ3OADFbG4s
DEX8ZhXf0aTdcggoH+7ltdKDUGndOu0XswzTq4lNnWyVLS60pxpHgCcdxbq0x+82
AoR2pn250xpg8QTjndjG+y4g2/GbWINtHRz+FlK+HKmebdzBsyVyaCOaIMXD9epZ
u9X+fO2Y9eh/nx1WpEs1RE++pBS3NBN8qILbiFgvOat8p9Q6XZEiQk6okk1pl1KL
CL6UKQ4t+xz/esufCXvvUm/fulePfz60nm2if/n2K/76kUTY63O5rI6IoX2ngsK4
5LsYz4ymax7C/zs0G6ze0H4zFT+n1Z05qPn6hic4Z7b0yieaj44VLGPKkCsxyylm
NqXPSqWgQiPCbdsNcWr37x1V+vlbXI0jgElEf8R+V2D/9xaoD23WH2IyhX0vg4c3
aUYYbEa8wxpRvXtaDYfx/F9g+3MpEwC9fmbap/PPkKpX/hUkpFGKJef2dSC9Ga9S
kjnUDquLYUY7eS18x6k2i8ufbj8JARihu3D9+PADMcGw/oUe4dAa32sQLjdwVhbm
tzMP7fJq2VJAKXLVINyHJt+LMZ+4Xyir5XIL4jSB0+MRYq71cNiiLYpqvz3z19t4
7yDCVNzJfuHXzHWHmsShr8wxB6JuoRU98zmY0LS1M0LOpm/sEciSJsefPV3eSLc/
sEU9EKtYOQmWwAbxOzJMav6dvz91C6YeIJHqpLX2rXtSUj0h2MAwkQOsViZvb2KJ
NIJ0ykfVsv/JLYv2xYKtsmeTyCEOb7hIYDKZLXw80F2byLm9oLctqq2Vs9TX6FL2
5skZC9CkcPf91q9daPv09L7Uvy6Z+v97CcYsPKwoWmHbZcOvj6HhB7R5bOUylPkY
+rDZgGWdwou9FElzsAEd182TZFh0f4gFAUiEHz27Zr0CcZRgwUVzvEJ3UmhGxUkG
6P5O7W+l8Uz/vKdlk+0UWN/LZ7llYZvkDk4yHgGGCxFVSde2Vp1BLGURlU8MbArX
Yn1dKI3RmgRXI4RY0eQ6t9K6Ts7h1vNl/3w140wHJtd9XagP8FFqxGrsEu+6kXp2
EHK/iHLY9vACzrCZEzX+VNK8P4bWWdX4H/wK9fiFDzMAD0DZosl67h74WwU8Mh18
24rwZ3csClf3lHuoO4wmptUN8ZTsi5NCezCo9F9UOSr1KLU6HHI/k7yKzAY9aTeF
81wQglTLFHcvW7cV3CN77PstgfP1l7cR0ggjM4PJBOGLdZAwSYSYZSK4FPcYYY2W
fVuGqOX2eJ1+GHUGVBaNnCQ4hw+IVA4dhJZ4709bpwRG9bY/6jF2siQ+MuFo8dl1
tdNgmxQM/GAYcL+oreyJ1vI8mjw0CwTSfx73XL/2hwbM5EEyBMyqfhRD8pIChsrH
zgJFpHJVruoE3y2VNziiVK60Ky9GyhxAG0ga8mM0c7SadYxzQJGM34bMeOJv1egq
QltVA/6X+ncPn+40IiwyajE8ClM0n+F6dy650R66tDT/ymH2QvAPpf14/m7gInnq
QEk037pgKYEw9EJNYRSV1T6PasHZTwjSdwryjWXBzkWmHJzjSWiYvK8rlkeEGJ0s
lCGV/HyZK5BtO2030ixDIvRUgwN4JO4cA6mnFuBg9rKj4j1wU/dFkSg9vJLSpUFm
mQJyCj/uBL0/BU6YBts0s6sp44jU+k9canW/z8ax3gsQeYWeSUeL6GBaE9QmGgQy
HLcnFkvT3PfX8QjPdsTDK4rxCi/TxbtHpigR+pqNnf5tHZoemfh6IdNJLVM5/AFq
1+8bl0H4PjzsyXps3gGMM8Ify8kQb5NCPAUQuyapwWMrpfmwbVBRyt+8dAkzLSqp
SEqa1KWdj1ZlX91tqIOHop6AnavfSVu0y9uCue8XdRhbR3S035bx12Q1PueK1CQl
aiVSLt42Rfv8kzN1NexqYH8kiVar7VlwxLgEpJykFA3NcsSi0kcxlNP0YR6aDA4Q
N4HzEspnOAkfszFoD879/oiW/pDzd+K/0PuXmEv0TzeNNzIIzuhaY4wNbivSBMdK
hEB3pPphtvxdwumMDAJwlV4WAvduvLz9rfqc+H0D8lxZRvXyhBv0l9kWcbqWVAgI
mKds4nkmM8fhJL21AqsKeKJzmTCgBzOp0kQZM1Ed0T2rhAE/N8JLZ8tEAIGrDMvO
Fr5/sStSaDBv93WBq+FcTDrYAOPnjCNYGgqiU1rrA1bN7GwYPlCPmajGDxkKi6jI
EFQTdcxYpMnlAPEdqTzV7uWkDak3xn7bSwOlHyb70Ddep4UEEzIbXN13tIWEAe1l
K9uoAzDwcj1zTIVDEYo4dYCzoBE2QBan7L3rO1Zzqy+6cyDF+JCi0YNzlPUk+gBq
IFqAX8DY7yuujFUx4SA0uP9qN/96kkn+o8tzLg1vlBfYsi7j6EfUsZgJS7eVMSnu
SFCA9YN+PYFFnKejQpZI18CazuK9SyjfmMoC60UA00fFgB5Fm88E2cRekHqbn06e
MgPb94Yk8gQLBqABllgoxqEVzw2aIkxeLvsSPwHbmNK3oOIvSpWbTgl2jUBCJwSN
st7LLhwFntyCqEPzJpmaIn074s/n90WG/aY4YJZnfe/xRLjiN9knLEIAJGmf9jY0
RPznTgodSBBbl8L0lEE646L3JLYlH0fhBfAoV8A5S09g9NvPK+h8hmXtH2lF/oZf
pug0RiIkS8Eb5xxr2mTt/2BuzgGsRfCcFvmG2sR4g1titrVLNz22w07k9aOMJ0v3
I0wvg3G9n62b9z/Vg3XOEXL/zHei+deaQHEnDKRdoxkC3E1KgKqJHTU0GNLBmY4Y
7jrSg22VIQBXXy/7lsgTHfyMyVUZE6zzwN3GeJNl4kCaVntftiHjJPfP7PLcAxAN
HlEuteigtstIfeQs7/9U4KJSRY/bmqVBlbtOA5uQQ7Oavb8P/BT3ag9RTgjLZ+Fa
qcPCqpYsxxoc9WnF2V44qdUKlNMmmMpZ9uSBbqyzyARExLKNkGzfEDp5XzHbNLqo
3zjakoC2gSRlxWrvXXi3f8vgbfi07t5rL5xZJM4oJOwzHk/Q2EJjXRYk2B2pmCzE
xdevG7fJ3fBk+2rpHkWKPV3W1hZQT/6kxj0tUaYuBA4pKpl3py7myQfOopmK85FC
jqFQSoZA5x0OSNLURNc9tmDALRlIg03lK3FY3wnw2p23HUiTXrawWK8togI9rxL+
fUKlYqtN5lXcNAXZ5KveYyF1OR1C3HW62H+c7Oz5yBqKqjHojg2PJPmOrd/6lr4i
Fg9c5ATO0ajzgD59R7zzm/gP1W3/ofv0jmJkVVfVgvtxJqWgT8V5X+nrrCGYAB3v
ojuklaalhxbHheA3U/aNwGLHUC3o+8h91WcAQgcnLZbrPku2F8Gl1gkn24CJf6q3
etCin48yr+ocOQ0X54qae7nFWYqiVtXpnVmtCXW85IoDtF16IAWzj2PNpso9BomX
mHaO3HcujYfhNfXy/gYrfhVWyZfJKkUNPm6r7TRqhSxhQtMIlipUMtT/Z4Jzn6zD
ymJNRKWmcj7G4ChE18cplOz6HW+bCjMDbKCAScHbA0Lp9e1C1nJa2NgRyJxawy2s
NScsT2CZ9NFopcCBGQl9JcKDppfFK0z1jbM/yHPJ4aEyjmaruM8SAqdXZn/0bRL9
OxVPYFogNpqdrfQ9cu7GMGkQvX8Pik54/Sf1RbbNMjt2Ips3VqiuoRqCuIYBIlOp
grV4jTEkxfl89yHa2HzyCnhmNi8LVhxIlk2OyJxrGm4J55pUZesOh0CGygk4GUa2
6ajUtgLUgs2w/LpJqSsX6ixmY8e4y3h/Mim0kboCf1Di25wpImMXtxD0saR325S4
g0oMl7dN3PSo4tG9NaUeNe62r70tFSInq+pQjlSxX3g4gBaZ1267Ou4R+D/Fz6jk
BqOB10cGxVcLFOiSmRGxjZhQAUYEQvd+tKA08OxuvP1Zr2sh2iEMhxRxmS70kkae
9BDz9Cn6OuII9Nmtt1nqoZ16jl7ZiJ7cjsTQ2YgbHRWiZAEKwP0M6wsOtCCxAFdG
NLs7eyl/Hjo/LCu3XsAYATEFEtFCzeYvTdnxL9Smwd0wV//S6N7HZ+9xuWYmGjsx
hv2gf8rx5XhU80hRVXPhWeCk4L7c2RoYUbGFfbf5uSDJ5jw+PW9BeTiJV7+jBLGJ
t3S8FBHZIMr7QV1XsCGSSfO8j6XbwavRwx3W3cyMfo7p13b6+URs4ckrWoNAeuvh
XF/w9qZPP80WM61PGvy5GYiuiMNcg6Wj3IlWjBgUS82wq8w1Thm7laHqeWCr/olh
xJZWuhcVL5s3kRAWc04gxPYzV0cjM8UvBEFjwihRp74sA7sEtpjzN3+b3W8e/8hF
uuI5Mo2c0UwVB55ELTPxzBB4HtBcONGWtUIGAvVzL2mfB7lp1EP1/WBkSnt261qr
6Oyx2TiYjWhZa9EX643CEjfa7r3JpffmuGqZvlnfQliL7uYNbJA8RKdD5BvCQmBR
vUfrgEjaULhnf4LiUK7pG9ZORnpy9BkI/7wQtYXbYqGUWqcNtr0uNDVYbo5cR+B6
OgwbOp2NKyZx3xL3CSqiwYfYT5evFWzTGvPY3KTbKk3QIQArAm4TuJPhSWbm01MH
Yd690HeBluBVUeJZuk+TzL5h06zCOaU5Yp3jBH9y7z5/ze8xPB0HglN+xqwKYKsW
EaQU02FDX5Q2zSPkzx8jvhenjtz8REWmH/wTsJcBhWUW0wK2RK6FqthRE79chfPu
11w8qEExZeiAN0g/k/LxixrRV4EbzA39GgQUQM35NCqGr/W2Ndk7v5xsaaGC8m5G
qWg5Geo8PwlvyfyjPj/6oxPpRI1JxXXfus6/OY3VllIyHU/yFvxjgmeHiWs8e9ys
pCERBITitUIyGPRuhMHl6O9JL6yQAAt2o1ffWd9Y8yVqfQ9pLRfZtcgHHtZ58rcT
VkGGQ3vEQYS055phMVtWXSaKIUQ21ZDiyHxuGjseX8FF2o8VeVOvbq2V0RJp3dgv
s4LPpgT4A4jSXpX5Exb2Zo5+1b6WnrSKVD7IsJ2XonpbYC8aAkpAX+1V++xXIqTq
LKOXSCaKN7lq+UedgcppU0aXASnC8SVSLApSuAM0jM27TZYOWGhrh4BUHs9L7SsX
VunH3xc75SsnduROr7iy0gCHbkKqw8Fqst+KroHq3QqcOYeTDgN24Nx09i0vmXC+
3wiBQdBclKmgL0pTy2p8hhz7J636gTln98U7tocPauxZ/phA1drV/MZ6k/UMWUqQ
VYow/4RE1tnoDr5dzfXLPo9y02SWhVquUEuCFxx/SSnSWr59g2F7eabF1I5Jh0Vr
GpY5oHiz2h6unZqHHVSWfAWBch502IxgMHy9xhxFuqguZGRqNUUNDnkE+DU0t60U
7VMB7aVnGUUhlfay4E4r4WDrY09s/eehoBVJNmSz34dUrF8UH+n7QV3POBbdW7gG
Q6LxKi9ef92TB1aXs23i2dEXCXH9j6FaX6y84GNVRR8K1yWFb8Zsz6sB0hIB+NKh
V9CLNiGpbuW/qxzHrNBj+MA2Zfmref6mutQa70VUlzB6yiwn4kDQB9SviDdaQR86
9mNEH0xe0bCZZm8Rt3J/VD7AISu2+hvfGEw2EJLc7xv11G1Hg8D4OM/XOaJ0saPV
AwU0ElbxfPsYm7E5V8dggUwmVqmrAgfhhuzJvAvYEc5A5hkVeQib78a2xbU5bAe6
zSTdIyatv9FFi05ltsIV902vway2KaIJuJdMEdBrHH8TJlu1yfUB1/M8z0B1hQ7x
YymLEGXvVfPn/FZxDKnKgI+ee6+77BaGALTh+NJ13d2il/dA7LyMjhT/cssqOZZA
tyPy37eCSsKNSU8ALZThILetEUHoN8ri6h+luhn4HgRzGUz8lyapzAiQ4GCtTvXy
dnRFp5FmXwyHdmF76QClywLfHnV4WC94DMquq7ER2HjeNt2Py/LT/Prr7ivY3Wjn
7x4hhxxl8cBPzlR7h7fkfzvOj7C2i6wi9mXdmHIBXl29G4DCTUy5rpyrj1AgZwkh
3z8CJK0mWIo7wEdQRTP69oBwY0La7VHmG2mkZCcLyC3fedYNRvHO1YD0u0eYghqQ
V3VFQoCNx7aacoo89PUjulaSOBLXUAojJhHd9cZp2Yp+JhOoZ00a3sU72R/lVde7
/S18UIqLVJlPcNUjRl6K9oGO0JH5NWcHcqa7gLJqQdtDF5Hnb+81ldfKiblcDxPE
VR/y5A4/5lTR4ZB3srTgzjVd7WDYc97x8a1T8VnTC7kj7tvypZvxeWrFYl/MVFrk
cWi+zn2k9bL9zd2dHo4zlNIAbdJUBKDrZy+pbBioayT9c9kvMHKf7SwtnHLHfAzN
jJQ80cNNF6L/W5zRKQrXL+AggTrx6yNc6GzFdUVY6ybl1pceVvpZOUftaS2E33IM
IIWYExWjeaJMeyFMCSKPM0sI8uOYiwKJ6uzAMgdEhDkUhV/td1eH8JSMD0lbs6vx
83K/pkfWLqiBRf4QZN+m9sQeYpEVXeS0UrImi0FBga6aJC5+7UG4tCBbdAQKa4Qz
gLE7c3VyQk2jl+fWK6ZeUFiAvPXZZuPUNn2Yp+Io8iP7cMGNdex256uOTNlw9rAF
7jizws+9SKmC3wmK5mhGunkWJ+fWEySauTWb4URodotHblLi4eJRPaXenpG7tfTp
aI8zTYTGA4B43L3D0pYM3m/xpJz1hGFf8DbcFBwm+Fh9Eo35IXOv8c8+Bn9IEeB3
doZI2q/HB7sG3AvEJWidRKddxWh3rlJm2DTV+H4pBF8d+CN0muWSLhC/EDUDDi3W
G9+2RoqIkH8kbxHHeV0GkIKg8sgRYpJ6HY52SWwy0fz5Z2Ysp2rgksRFaUe8xdrW
dSz2MeVd9CUp98auFmspgz5T01nCOI0UXwVqPnvFE3rjsntP4qsxILEw88PVRmh5
/pqafYDL+ocSNiAp4pkxw63jmGkU9ao9kalw77lfGueaTIciwW3KIHUkNU8+O27M
NqiMzH471Zxcb6+YQVjJmYbtIcrpwkofBiUskeKAtB/bELjULUwi4uO2/CJJ+MUU
9MsAqkFsNCIt6n1/s3W7vsHw2UKZGlIsgvyYibNxL20FbzGm27ZWiwhPVsFmYtnR
493cgfoQx1S95nHyciuGgbzMpYyPkOaEcrA7bmvLaiIuJear78Yg193h/vlpSO6l
7PhSKl7lER2v5L7/fnuRwI3d2EskOwLxUuVfnkIs/+gx1VRpXQjvlzyOeClqHsHP
MYbggc7XO/35eMr6LsHgyZ1gJHIYswrMATO131wnJUXaK8WDVXzyKQOvSs9N+on7
MhMHbsGaayQY3ieu4ygotUiyUTDZwCYTbuq/LBiIsbqCqof11FOtnLgWLNAGDJVg
yNCB1BukLg1kiqsLlwdegovU8lKKXJY/U06N9C4hnVYXGcOVifoCIt8UtRZdBV8T
fpnYz1bccBV4wfFLv0Gky7RgSn17wUxHP9xonfcv/zHlQyY6ZNKO9Hc/4s+H24v/
S2MfthXFKdcWGlYj90feKNse1CjHT914wCxV517En0dz9DliTge9Ci9NTq84mjwf
5SC6BW+CIN5w2ES4Puq3AMHUClLTCqNLUZ6UJG3ZCivsc3Nd41WrJh83nqBH1Eb/
FGUro6ccfKYLlc2J1BPybPudqEZL4saW80poZFhweKxU9LTaQS7Ri00GObx5LZMc
1dYZhXgt9mOh6SPB74Qgqp7eTWj5EpSKhExHKoe4l8H4IpNG8bQQF1cm+3psggOp
2gzL7b5Gk3B1XGTKSgdtr/tOor6gThwTT5Eri9Jbm4rp2eEEj+HbT4+Sr8d8oB6u
ZL+aMlfKQd34YRK6vduOXDbmCEgxD3jGxzUDrVxGAeselCipj3pWNH9NbzYI5e7s
3G41nENwaYk+wpzC2+ejoElisa3zA4ttrTKUFHWh7t69UJS7uKBczm3Lpqu+qtrO
TyjogUeo9Pn6V32/FXxnkeVGy9EBv77s99Uxb+f5+Tau6VGkATeF2l5d22tmvklr
UJhayPzvGUIQxrm/PNKKc9Yi0iTXyrOFTG1lXS+Bc1IXmfxyhEc5oHwO32dmCllr
zsFf73rz1o24Ig2GesSld81xKP7ROsHlUOjlfR2cbyqzTNJvWZBTf8ShRwjxRp9C
Mfd4tz+r6dvCG0lR4jHb54/a+RtLboYEZOvukCqsSx/HABNiS9dejFzflPJ2+Jxc
M9BfJXkccS6LTz5omfSfn38E3SHySMLremmQeMaRfjgKNfC+PhyI5Te5rVofY6qB
Y1Xw2ua9N6B2uTlANY+Ua/N/HB70RFepsenMMbjk6YGOmysnwAD/pS/H0g6eUSfD
rG7kjUuiJeu7VCiBuIcyxwb72Y18LnCllX4yDGy6bew+h6Aim4Em4iwk+2H27wmF
PJ6c6kUapvTP27HU4hnt2Atl+hDgPeqeyceiQm4SdxsnBR0uDx9UfAjErwq2Tcjq
8w9yIcvazT+Mu3APkGvA7BS04Yr4yc3f+Q1e35dQXZM+n/WG6uEzG8w6rXUV2UGu
VpnlI78O59ekW3LCXY7YGbue43eTtfq0i7wJMpiqRM20zcdWaXvwkwGEV8rcuioQ
kvykqn6KaODs7UOHionNiMCxcj8kx59yFJoqi0xVl/PXdK6BrDiwsFBAK12pu1g3
ixyCMcMzy3QuLneO67CDHIGd8Ndw+KVtTHec+jPfPl34CC4oRwsg6K1FmG4ycNxB
uCcYvP1BkmAKFFoi3dzRuy3+fs9n56mRJ+amdeyRi6ersQpywq1EXPlEmU+PknDJ
3k8HhK1ssWGOf1V5tGlXLpxtiTQw7d4OH/Xngf0f/PMvpld/svWYoE26xDUjbTbe
hJxhsineNZIVeGJvJyHm1fWeC3AxcF+wv9+3iW2jQjGRhHbe1WWx0XAKPTMBT0QG
nFQvDfT8NsqFup8Kvp/jXbzbfY2z3sneY6hwNzsGN9mgS+83ICV+zpCWtMVhUHX2
S2nvqLbOQgGsS8ufnNNcF6IR1CdVzRR5xBj8kOJch/C2FV5Sq8fTP+iwh3Igq9qP
GL4IPmgeNwFJKwbvzQg+TxLHtvPUmSWLHrMBHFryqFFczxM9NykOxp9eYY7/KXxZ
DF6ur8rqUySsojLYLTXgBKieqhzKVy21K57KGHutccxnRIpGgAaQ5BfAA7QszJ2R
V4cIwbYu2u+29HVV+nf7a8m9z+H5aHS9S7DhuO8AMzOLdRCWxAl0h4CgSf0P14b3
pT3mnhnS5G3Dl1wPYz1Sk2raT68N7n2X+eZvq55wNNbYueuUxvKu6XYLdniWvNW7
XLNeZIshM4ptqvOU0uXIT2yRAs1RKsQakitaj8IE8T6YkUSSyrzBoZ5quy/WZVvr
evv5578U1SyT7Q46nnHTj98mVayJvfPKh7reA6hbDLYyG/d5NjyG/2dvC46bMGEI
MVw9qsqeRV3r0anqoHHksDRR0TuFziiRJ6aV/DKabvYkIawhnypT5jEIpPWHRemg
yP+akeoogdUEICuTOXE783wH1OdQDLwO3nZd0b2q9vJOXoC6XbsxEu1Vc8aYFef5
F0LgoyKQcXqXy8sZGA0KYBF4OlJK7Xf38KPEETUz0BxEDpfm9bIIKR3V+Td+OkUu
R42kPkS914rdhSrIGIXouGlU4OUvaoRlpiDu0jYm2Z8q/zTTOXFAedG2wiQ6lM3e
8j8SdomIppH6tUBQsmWJ+a1I3qCvmmqAGL3SYt9H+XqcnKPPUGCXRCwE8WoVg1R0
Cm9li3aobPbUIvw8onH5F/MaHxzcHzF/Jb0OEzGs2dyoS6FgzELLpDjayC4eDYKU
RfV3yqgoe8MTa/6ahNCVz1g+8Teb4UotbdZp5ebZa/X+Sd0dYzMpQram6mjzE7I+
uiqAdDi4wFxwp7CA8bjKRsNPoE0TP7VwzCmRc+vNcftGtfbU3UY1HG3MjOVIr+fY
1AXE678nnsKbhoaQQnmkkfdgPJn9FX/0W1dhf1LzyS9KbSBs1NbS65+3EZiT3yIZ
RLGLkF0bNb+k9nZnkahUkUNAOIkd98cHakytVtNRs89s1uUQcaqMvQxvYWgMFbqy
VMFD/IoIf4hpfzwVkQS7k5hnIxP6L8xzeoBVYN0GkciI7BwM1C2dqD40q4DvsB6Z
Hec/2HP9F6Pk8VMTjxHiPDcdFfFuTKWaIOKW7tRxIEMJ262ouOdWfLOkq1XjYiXY
TPDQdI/lvRgt+DUspG/5LX1hvGy9eRwDR65Myjpuh88WpgvqH/Ih0cvHAytGDeG+
r7u2yMIJAlakPgHICzwp0vqEEHn6X8SJDSbtlxKuyJODxMBjWIQaQ+WSaIcvwGCR
IHHHjKWEZ8XWifm3uhAqV3Iko5JmFuMHocphWCES6ZktMHO7+Xo90/gRP7p6YB/S
AKNRyK36AsdMTRqe0lK8Gkogbm4k/3TUlqhNUesiyt5CON+OrO+HJmlHqs/sqrfZ
nzGDgUk704TUHqv+opyAGL49xyhaTJFDMsPaaK3JmeQ/J6GH3otTOgcIlw9ckXFs
ojGYfytTz/L05c/p0krHbC5tLzzB84FUu7d4gygpVeX4u0jU/sp+TbfsxGEaBZ4e
j3bfEQ8KgHkePF/Lq121boj2pEP4UI+YbFjOVHrEvwzU55JI/qI3ZRh0Ulug6h0i
oGz34BeXMCSDo5Ht3dX66x4+wJcLO7G0why8z6ZdbsJ9ZSdL6HYtGm3MkTzhZr62
hc9omykjgbFWbtDstzFLZOXJJLRaN6tNddCjBEKvPEEVD99joiNum05kCJ+QY91v
3Qi9To3GqLa70ljoybh9UtJJ0ppc98/LN7DTwBj/rxxZ0lBPdGG/zGA2cLBgoV5F
OiNMddO1jhwN1oC5Q7Vj7ikD1S3uWt++awm8fBwzYk4LhM1zIvzJn3oq3qYSuEOt
qDs7Xwb8KXxw6vY8p5hKia0/RgGs8ntgqxvRN5TyVHnwo2DrEAkSGvu7tHicNOon
uGBXzwPTBexQNHCf92VR9OxdKCGOOXWVhIXnz5zssMm4EBtMaostWOqC/MCd1zEo
vZya+ILfZxnnoolNVlpxp38Z5f3qN4CH6v0ExKnaDm6Pu95eeGnkv8cE0FE7L2Xe
5fQJwEDt7PkNoWcULWZBJwnEl6YJ49ReqzCI+2tGAdd4fvxdb79RVUL9vwNwnZYT
5e+1IBqtxLx36vK9j1d+0hOni4BlrSIWcJ0ohB74lriYkr/Jaqz3ES18ORZ7vvaD
3np40F1pL2A5CKXMixuRdu7E6mNWnZjacO77Va35hg14FDTieYFtF1UlCBjBY67O
IT2OH7n9ZmD+exkIBRWUrvz37aUJoYMitqwFYbzqN9OdwKxmcj/Ld80uKtswFB0p
jCTLqrDyjUaB+VODjgECRdhGz5bec53D6ztECz6NHWN7ob3VDn1RY6v1xfIoRaoS
zmXp4gbaK6dhJkz2Hv3+OGm723DtE0Ehc8BYkmIb6XjXNj9dVE5CBLx2mRkjsCnb
3iqie+C4b1fjVnwz36hbq7Aczys65gLAXPkUQut+9zVEJvc9RBkGbwB9RN8hLBCa
YVFQoiourQP0ZglBAbrhbuJ/PHynSu0UGglwvNkGJuM+7lty/3frXusnJd1MeOFk
CNtMHkswW0ytNkhq5/XuH3LeimvV5eKNk73nO1hQ25pHEeu0kleYH6qcDPiPT2bl
UvbyosWz4oG3adYshk36mg+vAEyfFCvJQPlPk4mx2zDTL5hVjg3HZ/14OFPXH5Np
i+JjH7Rkf2saTTJb4WtUe02UN3UxDGQo7SvHdntmsnS4Z0T5GSV8+EF2/6qllimc
PdUZMF0+2YGiuaoWxBIYeqokW0KRdmN8u23rrfQnMv/J7SobKproFDPbMpGnnAAw
M2cJ0PjbjU5sOEZL+xbhm8wz4nd6fkoAvSapn998ua6kyL8cRsOzN1l7NsaRoTXn
G56MqX3wwXLFpT+BrNEk83hA+alulnWN+JBTCQdbLNEfAkq+/RquGqRg268X32mj
46mltondeBs6m3+9ENZPa94tfEDztwWsazdt+00FoAXCVQxJvatlp5i/XJG11Bye
WZdmxeqs5kIVrcybr+Irjir/9vIoROR/aqNWnXzx5of26eV92G1r/YSW0zNzFR+s
DTYVuTtxjQ2Jxss1B24uHaNCbX1cXqByB8gKdYkqhhWZy+7h/aEG9INr8qW8ib6s
Ngx/44i2VD8xvP+7JN2CwhCNiTqitDWxzFTqf8INJn49HKQeCFvDxZgAGRuI1fJF
bNB78zsW2VF3yTnpolmuHhEoFdXlyFOmRBfhTqwDJ6m6QUXUV64uFXk68/xppCff
eUwDHFGZp9Ssqjn2oebcpjHUxpOV49GCAFFG4Esc7p36qB0S2te4GyG/UvSUBzek
OC6WIeve5LEzGXxLn+EcYXkLzgFxK0ODcmCjgfvnreSDJqIRC6U+FF5b/AAM/IjR
DipJI1pG5F67sBoNHwud6kAqLNDdWIjzohRTB1mI5uOgZXQt/zN2GcU7EAW5DhJh
P+XcIqjcuYY0hKhqnjpoLaTxC4vDjt+UDyk7dgPRk1iCNVzeVbZEpAQCb5AoAFO+
pQ35UMmnsm5rKSSAjzVQj8SECusyE/VFvEmCCJQ6vb0knTbe5lsQYRCQqMYBSMmK
M/ERVMYaCnxjSj2TrsjRKFpOKgqW7B0RcuTuxjQEo+dVYPkp3K2Yek9YEa0/SLaf
EiJ8reYqodzYTWGn9le/S7gvsDj+uvtnUCZfAiMHnUY5ngVCfPZ9wFrgfPTnkUGy
KwTv7U+anqDPZ/MA6HkCeEtXD6INHxBv1xodiXu+IARswInHYp/7KgRd9Fva0QOw
IPgMnN4lfPzr8ovajGcbOlZVDMm0SqNSMZW6Je8lxq0ci1hccrV/RirrAEfPnM8n
Z1DAFUXcuRBeyGuS3MpR0do0EY289vi6a+TLMmzHV7of3UvkhY+kaj50SWN/X3Jk
KrzoqyQzxvAfUHbWeqyOHS7mM0eJQKY2mR/6zH+5DflRTuPOl1Zb6SsBp92n03P0
3Zaq4Wm2k5q/jV94kAaQW18msYTeEIGn8fnsVsbWsaD/MccSGK2nWU1oUj0881Mg
ol6G4ma4qTSi6L4+i3KW8KtbTpTh+w5xcmLaR9p8ZSiu9lW/9cIX2aTqW1H5dt6t
ki0dt3iXflsefcBBHhqm01qUgXgWuq6Qdc/nZ/eo82VAc9395Frouy49elE7oc+w
bwxjVXSjR+xNPzGPlMYCy5K+Tnpv6LyAz/LTJCtoOwJBEqpXeQUKV1pBHUYtyQ8D
b3IsCH2UFoRsLDd9ueEZTlKBx0R+oQ+GpjFzyoaSy4vr612q5xvfkCmLzQqtCos1
8+pePBsFqTzahqVR19BJuNbyYc5RHZz9qcio0GxM6J2MnxC34kipNNtvh2VvREcK
6OQH+ENC0PDQEY6BMcFXen54Oq+ee8nxZc+eays452KTgZSQARGn0CVLO2vjtrkQ
pQEo1eycWhJOTABMsxeUIxIyn2SMivfNW9wuLPqDmzu5iF6d2oTruohpny3to9Ln
5BXKew9nh287fcdn46t+Yd6fqnNjSNeEoOHwl9J36PJwKnVdesCd1ELoABsSdTd5
V7CN6dNrwXjdNLOaoqNEdcZzLNr++mx9zWIiWqP5Q0cea3UbYkjhguZRBJMQSI4A
jfH9PcsLAIzcDiNOSPfrSXFM1m6rbcrjXpY+d+Ybydut1rw50bYbazSSfXueAqAV
lly21WOZe0aQPmHTAhIIkf14l8BSRUxqeWNYVEGY8XvzKoh6sqyDvz+sHzZfYxMc
rzl6mPDcfKKyTSvn6JBXIk9HHRmO1jYGsdxfzmDg/FXFzkm3PwZhrLWOFV5clKSN
q31pDcubl0eTV/lbVRfSiWWgVO17Hthq4Z5+CKbKtHoaGZLmgMx9KZtBg6z8C48S
PpzWWuVZxkrQZijMxZSSljGpviaxzFy1Wd9Sbr8q+k3PJW5CiwvV9WvDNBbrc+w3
yRSK/4AWiA3+Rzjxaj7rJLUSNGYKzIn1VNsqA48mfiJ3NlLqw6O8/cfaWmn50vu+
9PH+Dp4YLp0U15Z5tvycqp1WTl8qqkO0AB5EmtiHdqUXuvkiU1u+VQgw4dGFiDx6
TQst0mDYD2wZAhhJF/Djf0Yk63rhMbgpEsoDrRGrv/xC+okEBE3hdnjoYGbJg9a9
6O3LXHsU6RDqtOl3cU6fTgR8JesyKqPuuFn8o3QlZfDqx5GvlH6fcl/82AS8+Px/
HZSZeZYiKxIbjsn6vBcZzVCZwarQFsBm4J1R0aSrc7WIMXwpC5u86kMCYjPUrJ27
TR8tAE58lZ/hkEMFp3LVLH7s5aWXLFsk5G1GI1FbL7PmCR0GlqNljm66LPAu0TJI
bo8ocneAze6B0Ftlwtzauj4Op7zBazueOBseVqpFO4RnfhHV32L//VR/tFryvqFB
svl/FgSSArUCFZeUN5DSGZcUBktBS89czNSKCkA5kBmZeL89MQFD5BYMQClyOL/L
Dz2iACQ6NLkiCN6/ZjMmhy3s+78rx1OAaqeZuUz99oqkwDkuTx5IhcrFIsD2pDIy
7hDkE3EbWIqSzMjIiiaZGraPuDGdKdGRCMZUtBIpvAJMXckbfMa9rAcnpxgKB1MC
wxkKQ4qrdSpYlpE5TY6mX3ziDlljuDRZFHdlSlRNxvo2zmDGGjAup2dg/Xeqc7Hs
tmiTjFu0vFMMXq95bVRMVM3FuAzEm91fsC8HJUIwHelEvsT4Celw1rCm+/jW7noP
4zH6IOcwyyfR5OtfVXVgnuEKKThsM7B5qTig6D0Ksx0lKjFk5Gqdkj3bfsJci3D3
Qb2wUns1fGFMVMfiXix6L60lHGPWqtOda38KMy0UoNRWnLcZWPuQnnKIvphxGsNP
Yg2UufCjfkg/spxXXkytcWr7fcoMv+yBXkNYlUxDoB8xoZiCmEQgaxqsZmmTD9cl
YWJdaboi7t5ZV23K9iGZfmxic3sgRLLNGcvCUeC6GFgtus09SdQaurM0wjnyXS5O
FCMPaXBxCPcLgyJwJtP8X/2/f+G9PcCkvJcqy/EqqoF0dL/dzYNsWsPQeJDO1kto
mpVWKHYD6kVEkDAJQnWgUIKZ8d8WqjRHmu18NeMmfCBPXD/BL90KI310PKiLibYG
pv0QNarwOpji/3KakQbnGVy43NuC/O8JmKudCdio3eBggk+Q/5Wy1iliAfeX3mHl
NnrNaxTUNCkrEOtsbjEPUXbws9Ij4k0PpzGcdwvjW5UKZUKD1al+Lk/B/+MgN6KL
HXLBwJL7yRGw3qzzS/plTrAjW+Z6rp9ovUWmEnvi4WM2yoJLUpStudcJBz/JuMNq
6WFd5zj9YX6MIvyEGdlV9MIgJYdjz7z3zH3NoZq6ewDBGWAJCKegpC3t3bRLziU9
lM/T1Vr05tsGgRRbIX+2dmJ044J/uceLjHPHEzwMg8bpvDriPB+FmK8BpKInr/r/
D8wZx4UqYmP7KQBpZgQ/l7c6+HAmfUhe9Or//iJ2Qg0VJlS7IfUgxp6MUmPmmYCr
S7iafPtCUIahJa2JSXlAeiKKdqMv3y6fayscM8FRBr8KSoOkcE42BuDLA6vXHwto
vfG7UdFlfVmTO1lcGE0LQRHzdbt5p/paa5aQkQQpMrvySMDIhvvacmr7HEJqDFQa
qPa6N2sAWICj9LAcandWyYmwDNETVpfD6M7xMOtVsVIn3bfjavS1LDGoYlkNTigg
uGPD/aHieyHBkeR4tM28ERoy0cF7e1znR93BNdyOEadd4/ms9HRPLvJLYVBUkGHd
tOYzjoOawC9LePOtKrTF5EJewzgThy5oV7NTZUHDjFe5YikLkxH/AHkFfUOYtbdM
gGKYHG5qit8iIAR2l6CiUw6ac+/EIRdgsNUvGl0xK6PvYjslkMt2su8p91rH2/g6
DWc9TgfaBbVfCp/HaYLjNq0p66hRcGDBvo7ldTvwRysptBZALhJTz99DCJPgTnb8
D6Sd3EH9e6EdjcXcNVojso+QrrGQCO/FgufObTMgVco1IeIndk1ikzzs4qXfroLO
Xwqmik8W7jaNzVE6r1RJZkpirKwMpy1O0zmILjzHuUT/rfxrcqgKwQgBQd189Aaz
12NKkvwnHeejFFDnnPTkYhyn4LGag/Jeo+fO4dJxTbB1WqxemOtyCWVtFu39DNkX
xXf3EI2yzhFW0S15PiwxV6Wf9by+ARc29+0lWRheBLY+8GdFpDQFel0VyItN//I7
GKMhHbIrbVTMo3if9Q53aKWsqOtdBMdKH8eUlJPCuoiDBLuouRBCxIKBTZB79Izc
tUUPHU/kA3kGmABZLkTl2AXVvsyWFzSAsitSKgx4T32QksgBoQWAKuYNuKnzxw6C
dm7/E7VJpS94f//phymB5wmRxLRXGEzY/0Cr1YlFxTvd8mgm1CR/ThDXaPJA7ruN
BNxonzhf8sE2r26AEknAkfcBLlUMPSzKJSXkpwmogGuOsa8bW24ezmT5KhSxc05X
InXDv6dHuR/p3RKGCwL26qqlsch6qbAdgwc4hdD3LV6nrO/pJOKcTl28nB18tO3H
4juAEyGl+fq4OLWl/J/9Bl3zv04vaQijAOZDXqgUhV3BEkOJh3qHyYoRbDKzq5gS
1I5aT9ENJl+EKyyLo7CzuR+3oJSby/w+OrxkwNxYzLAEYL18SBx9ubTIdn0VVVKV
Wz15d8dG54gGeuHYvGhMNXqern2luaDNcJ3YSagIqgCQy/1L1rjvOckjGx6lDbkD
eUMiG0o/4Amtwcb77awfFZL1chNAPoRds+qGAEprWpoEaSC31tOQqjb0jkvRjPFK
b6GrbIsLgFLBGc5EItItNHIwNiRaWKJI6XEgRsZHC3kY1Mt+KtohXY6FPg4QonRx
HMGY653sKlfmHhLos4FM1Vecx9zg3/hiBXSngHv2J00F2GBFyPirFDXNA374dIwD
GbQF/k51D0HukmnV8VfODFmqfzLhEHsuseo+S9Bjx++I5Xp1glm5c2wSKbGKLW+d
/i4l2kvvnGDHF3gvwoovsu9omL+MKmvg8n1J2DQgJIbxQdFLRPJjtgt6hTXGYqqV
sa+2peBEXrh4YPHYgnLQ8s/XdtG/sunyU/+Bqon6evW9vBHB1IY+unP/lHTrK6lv
5m9R1+hOC1N/eTvoIVK9wvI0IJSa5l+a+5hHhwYa29tZNFJhh4Ssrl7gtrNbAtZO
8NZNCFnYo++qDiZUdtcEup5NPR3lARYgPRkunCXm//TlKnYChYxOhzhygMhtW5Rb
Va45QSESR2uf1q8VsrYnZnUibkkK5+BtqDvQuB3THqef7Zb9B/4/KEuiCvZfBs/9
E7Xhl7gSjfcYBRB4aO4KQud7VwRkFB4HOBRZDL2GQkyJtDfKg8Mm5bItrQl5B+FD
C4n7j0TcVyyzd3/u8UcjuhzeILaflmmMtxebpRb1JFUp4qT5sg9cAs9+ffzpKepk
m/gOdpKLexrlRTOWoAnMpA/Lg3kTImNuxrq9brt+/MKFlqkz34RCaO9Kg6i7MdS7
HOa/hn66Ks3pMKUbsVIthbfTy/K9NksB0fDtCosM3ZNELPbC/O1qbN2d4VacQ1N/
sziUErU1ai/jDVBMiXbs1vFAvhtVcG+Qkir49xC79hVniv771bc7zBCy5p+MI+6b
Njch1yZXeEOy8izqdeiB9279qScOK7fFX0B+klo3FbYouFPCJxzNRPfcmSszCHwD
9i8xPcIdbJndA3ohhxoAzNHVjTY3G9A+UhboJkk3MkxGPEzgfKjuzMm7IWmm2VAK
p6MF09KWmjv2OSiwgSaFcqkdjYqQU61tuMMPPpKcPNneGhsj4A6MWLGCwv/M6yyV
JqKA/X54NFphr3CHmpgeW465jygw7r/TwC7V2tAmtNo006c2OmNtNhS8fwMUVxOp
7siiEIdkd04LjF2BklCsyBToN7GGGKJ7HcHbJ9AM8xk6bKOQLwtfgIJEhixqaTpj
YvjMboi4L+HVg3pJHlpKdvEYOHtCntkL6wK5KkqpKHq0VAMqoio6Rf4vonxN07RT
tqSVB4XkJ4xu11+Rb2pKLP0WMr+TbTbjxhDjDse795IcG/JtK6fo7Bq2oENY/qbM
gtoyB764Lp64PvnbzQ5DD2xOASYti0g4PQ4YW4RyC4CCPFaeI8WFeQ1ea0YPgTh0
7S/+vtuLrlzULIanegJ6HKOgkgNFW7HIVn6NK/aUXgte6QtWQ2LZ12j1d9gniK1o
ZjKMsWHOaE9yr5CSq66BWvgzUzuO3FCaKurnK4CtBTNO0IQDvxcHvwd/prVISVWg
G6WP8RLG0JkCEJfF1ANu0YKBxcdnutiu56sjlT5Phz5beuv+ns2/AwHIzQ5HTg3F
9UCvxZMWydwMhZyzvkVRFTh2a+l5rdvelu6kb9XnlDTTaVTSUeMGOojHsxmPwNrX
GUh8LbMwAyD/AFMoWE6wCljV55Z/Ma9P/60chCfEShzb81CDZpCmqKiAX0GNwNU9
QVl8SWd4sjDCG7tLqZ4/T5K3z+KSWNRUDw8JKoMVkX7CfWQmGCe10Cwy8AdxD2EB
oltfQfl7NQbS6cU9Tb6j7QhJhuyHFG+yO4/V1l0/40EuBkbuVMmKSL3lro4N7qqN
GEcLc7VEBu6cnCBprcBvi1PmS7t8yjchNCNRTQVka5KjC+QGlfcz108H/S3he+NX
2qkqjmCU+xlj3nBKipz9T9Pny703h/d6A+zGAFyGvP5Kg+Y7qqDNkFVibHzozKut
wYfz17Fm5HqS1FHBa5Monvv5ZP4u03DlX8rKbI6X/K37yO5sUujhPgqXKFtBKm9+
BauD/b/LTV0baeohfAFf1/ONbSlQTLZDulrT36nefoKWYf43I2TQVixvB3LOMeU9
TMN6Pzurgc4nMCyFP22T/3/c0uQ4B8JK8Re1jMcJpm9Vl1rymnIHGLHN1+xtVqk4
eYty4cHwGE85NwnOd0htjM7j6LAkm0rGKC8enz9TfX3qtI7+Tjl6IKVLJxOC4nCs
/FVhjiQruxuODMmwxS34lDO2C15ZyNDtwLIXlHUiMOOCSNBV3oofAXzwje5SACj3
EJ61hppO0TybA/2bY/h9MgCWXB9qcNE1nxapRUAKVwqpA0g2NLj661NHy45gANmb
i0HEIpPSDrAn9Jg5DbPYV/EAf/tMESphPsToXxVitNGv0vqBRIIbwHzLnegzrXvk
slH0wXaxGfJBR7Kw0ihc99tImRfAeMebmKFgPiO/0KGiDPbO6RPe3LvIZVus5xLW
zI4Jb0IjxnDbOXVu0ne3HEtEbzb7kxwEgIca6AWXPG75ksbEIJoD2l8pEqfr3B06
cSsvjpTmoO7KJqDYP0GSQnDgzs1fsTbm+0+0zYtPLYcmWhLiiA2mR7zz1BvhleVL
btmyAE842+FwC1MGKbx6xF9vPFdIRU0OW+QnyHXj/MD/cCK2YgtlwZRWTc6ZJJvR
Gfi6iS6dM9pLK7UqbmfA0WC6orPgU99cbuFMEatbvki1fQTidU4pbjsvcKRSpwax
saSsFFbwEPvPqHVIjApzznygL2qAWj9HjMMQulWfXQNQCAbYo8fSrlhgqIKXqUp+
PIaV+a5d0LQdujF06g2PNPiqSzoJQPVztEeuPZU9Fd6i4whX7dSDf+W1+E07gDi2
zO/3m97BBqSUxty/Ct51A6/Mf1DAWweOHudDRDh1ed5XPTIqMlxh8UGyIYImk5Vj
vdSRzQGKr/t2ZD8VH4AKLqPqRK6PhNg6wGyLUyvvG6WAfJFqsOIDyTLh0rzCZraL
N0VT5D38EyYWjG1KHfqiS0uybSNgnH2RQkkecGWt+kb1owU0+Xe2ocMCdQIfQobf
oP2CoLCs9eIez4a9kfryxwFwSB+El/rO+PQMhXbJEmmZBwHG/J+3Vao9sAmPzfUJ
0/QU6dr+6VwT/buDGqrp0WSfmieCT/E5xhuJ6XpGeDXf/vRN7LpBu83ImfZ5+1e6
qnL9CcKYrIIcWZGt1ovoVyEncc7a5MmOxhGnc87E6j4BUsqwBUJ/ZViSVUIgorHF
5VQGAFG4MxBwOE9fmytb5aofrjTxnQnIR2C8e3ZVssfuprnV6fmqIPxgljvS4R3S
y8JF6h4+l6gbKahaBPY2PP4hyJZW7MKLX3amh78YXo99eFy6AcEbFxaL64eUTsNp
WYfXwNp4GsVMxh5gnPtHxW2DjrpWv3+qhcMSK5HYtx9xpAZHDp/AZgpr5d/I9x1t
DuDHeva6DuXKFy5FXgnmj6RLwBvHzCGGkRqrTYby2F/YXFqCQEc6vs/7j1ntDtbZ
bmnh5V+QoJR/A7pC0UdqwaTg88hgOlVC7cUt18Ih5B9z3jQHhaJQNF0Q0wQob0BR
bAY1GSKHnlQS/chOLoOPgVZVz+sD+8QFAXFLsRCWm+rmlnYFFfUCaLe5AR54G740
CmzTGSoBawenTLADEj28XdehGKec8YrTjhi/aG8yUi8VKYfAe9QsQoMwkEykMuQm
UJNdn3o2To8FU4H/rCVLm5PYJPShgp9KsEa4MG929xsrsh9vWnT+z7RyH2GNnoPy
VfBICtH0QWMbUEy0xZK1+Q2JGxxIaKMgoQt5kAYb6FJ5yDjjMT+ggZIclZ5xpqz6
qqsVuj5YxLiysnFgU3Fku2H/byHWf8j9ArRf/GVeJ71T2bGsUpyOhMSWO6ZRfXUm
21GhlP7rDKp3ngFjSQe77UE2k55RB80p0oRVuIt0k/zV/sNJtLq3iXwcrYRIU9Nj
YppUc3ByLwhay9Vt1dhA41guHpcwU7ia8ysb9HDyBzfeL9WVqENEn6LG6YCbVf2t
jOOvxipL82ud+rLUFNHOp9tOTpHkclJzk8QNdCEUteQt7gAimCG1oi+w81eYGCy7
Nsh/q3LaeMX38tVKf0BdJC4CiUe1O5kYsBSboJ4lBG26/AixOFcsfdy29aLClP72
OI9F0h26yNVX99dlBBjjzSuKvLtFGFHe5QID7Wfzd1kPsQe3F0njiE43OMlSdrUS
huMySWz6ZMlc7WwPsViPfVncT/L9RLtalRHBPYEkgm573lCxV6DB7DZQpFMUC+CS
Grn9kK6mtT1+XfnvexTw5YtEHGDWiA4hJ0YqhOD5dLFsi6HgQRv/4R2h/6gCB12C
0geRE6BVkj+sKoErb+uby4WTK1f5OZTaeNuhzTuwIzF4Jix3ZN8HnwOXQ1LGD5Zt
enVt6Yo1m4McZrbEqhhLjip7l3ZACqFyya3BqgYUJGEZbW3bHWrVbVuvL+fzhxEH
UrtZTJM1vszEZXmAgU3yXdO7RvmVbMjgNBaDYYrTsA0lgUGIDHrisr45NSaK8ojG
Wp/u2L+y7rDhhZFZACO7YdPWIH8d4MUe9WRBWyG0T1MG803LqzXf0JfDgR0JhXsn
3EafAYuak5/20SkHxUV1nu7nYjJ98LRsdQLWxo05FaXPNNbjLfxgEfZ2EpXOnE/+
QZNS7DTyQM8TwC3YkgmXvqsYvImqgAf34DaXQzKJd2GKZcDSQCHrMOLJgx+Uge/B
Hr71H3GN4wQV4kjkUglU68XPqvZGmKSSdXa28EJDctcT+5nQN0GWgIBuqLrDiP/A
JQB7mAVVp5ykxhKIjohYykiFbERn/HBPt5ldx4gSYS2l46QUISh95N/T0B+u3+kG
LGlF2Puq3y3Lm7qpmzZbxRy7y9p2wSYpOWKQgFXQpcadS0KvqXmZx5aigfvT9OFr
tq/Mhaeh8Bf0deSnuJpnJHtIMfJONOr67iBGOLlJlNe3px04+pByePcxchUuNl3p
cMN1ECu4C4+EdQODbaeooCiz8dnuWNn1aSldpDb7rcW2H3teziaaECjJN8vdeoS8
NVDZJglUIglqubDTVqvgkfqqFRZlHFFOMJf5+0Xb3xLmEaTaYhaIg55q6rVIsjP3
m/jgrQbqTGSuKxV1wKii3Meil9g88BAwRcOLu9RHSh2hymQcYx6dNivuc7ecaiAV
XjjydzUmCGRood7kf3WAqfFRJ/kzv0GLhwtK3D+DocKPHR7+T+iaaOSHBZ0xtRWW
B1GRAYEriBTSuJi6C2lAyR65jqKp/2kcSpLPXuVkGaKpVtauPYlXWDWIPEAwTaGt
E8e+rO2CwEPIsm+hirWNjieXlYFcYHV7eeXh2deY6bRbyVnTrkAyWA7r/1FB0neX
EglcQHXH2Qi/blrjQiSQ5VOtrfb+XyrKOs2xDyJlpHYWZXegsZ547T9FbiyxoSHB
n/IZU1RQ9PRnjgaWPDJVScrVF2MPBNT2uEcnONpYQEGk1a5t7HlHH2p6Tf6qoTno
uwM4GTHL5cTl+2lwHqxWkXgpZ+6GNxlCm7vOjfWAreLKewIbe1Cun521qkdKlJPu
mepzTuvibPr3QiiSQ+tEw8xqZZvs9QMb5gshP+i39a50D5r09E1eTr31dARsrDbd
OaQYCnCbw8n/9/M8vpF0UlJt+86eizBdy29W+ORJxi9dHOkB6XjY782ZczuOglin
FIl97ijXPuMMgJ8hVdFhZWRE4dd+7DTyUigEEhvgATVffzqDqHB8eyokfJy9A6hJ
3CAPW1HqZXi/eQ0CYbLgCE8DG2a1utm1K+ryBJzan6apnDycSDkTADota7CXAjfh
jCon+v6lfMj7ZEE2WCX8mTIrBi5cDQ8gWh+S63jLt82pMhtoU1gVMAx6Xmo5Bnqm
OaaYU2nYOvOP7kPDQ/PRcDhxjp2X7fTurtVzAH15bIbTkYxRPhtr2mMDoHQROlAQ
JZCgtPGSZNyES1lSJ8kl1rjP73ubWcXlKADVOrfyFKgiqcTwTiJcevH9GIgAmPHV
0XTfBRD3ohrlp77/YNHWjGbFAf/2UALFvJVb1o2rxMb/pfUhSHf+5vyH61ezRNCM
Wi2RKt1h7PopJtxroCzfGBjJq+OnHaiDr7GXUelCp/ZPJ1519TINl8atzF+Ry4bw
kVETrDRmflZdMvRl659sr6e+M2hyKE3bCMp2QE0kmEXgPNtyv+WgZAzsXLrlfXzi
cUDt696v7runyCWGW6do3hBbpbEXP8oqOmMA9Iouhzl2DRhDI6JMIHsnuNh6fOZ1
tEYepshAbwB6HIOoKzH/VATBKS50w0PKxIOQMRIfV6ozEC+sgN+d+fiL5je8Kv57
w8r3ZpkXoB46jls6UpkPQJL+yCY+lX5VTfyCkHccOZkS4iGTXc7wu3a1pTVq2Xx0
niUXvSU4Y+NJ0a7FMLJjjBgsLDzA12ueQfER+MTnUgkFp0URxq3bWgLObF8pvq+6
DA2kdgfQi7bJP3uNfcKv3jHDiIGGefCkHTAwHRs54AwRcjuPKd5SqBjDGVvizlmn
n5XReZpOtTJn6bkUtIKEG4K2zRYQ8QgOEz2x6GucRReDFvcD3cvm+x/xvH+6ITfO
jyFSmcj+lqE7E7PpRjwkiIDt/LFz+KdSuWbbpFw7uSuvjt03ZrsfRqer0y0C/onO
cLh9dyf4uCf9j20WEIkcfbu9jGsGAc3GVxIT6qei9KnSSjPTV/XbzXl2xtaNu5P0
qjbnhDdIs53ln6Vs36P4hHhAquEvhYIoC6iA162dccBhaNRa6je5M2GKX70Fp0lm
+s05CazmWk0TCYFCcgz7OXCY3MKHE59D5OctQ41kIvG8ru7gGM2VtPHEWjtSq9vz
mCxndA+LsD3saboQZTEbJkT6NP8MTqgGzumegjXr9pDb+3pY/9mlS+xO2am1uh1+
vulvw8ynlYBCMPl3RNoXlNorrCq/O6UZnFQiUHhwtDoh7QZbT7Sw+XQu8tDW/X5A
MVBpdw6OCMz/nQCacXfevBrPF+YiH6M7sQ3zJX4wB0MxcsLhxb6p2UJev/R/+uKW
95eTvWVrS4ZpNydZFi46Ghy2RmsE0zb9WO6/iKHRtaPLRO28w32STVOraoQWG8mn
AQ0BT1l6YN+L8En62VtRwRkxcRFDTJ13NnW3kbiP6A3VctQKmvoDAXlxgaxXj0rz
WwcwVFQnMqgvbCpFfwSgH+wBWZLacrKDhzFIBlfKUoX4PMH8tsv0hAT/mPp/KIqa
eKSjoFe0s+FhNcBArr0LaYDgF87rAEdtXnn8DLszTh79oCHYVhEXjS9GAuQqCS7+
/mI0N8fV8REBJCTY7SCfegAbD435zLBeTNUMOcGJOWJxrUfXaAi9H8QkjmxbaiG8
xh1wYMdY2SbatcUjLTxtNlz+7R7pKjimMRbUGmcVY7bVDqYQJbzcH2XSRPXgTubw
SmEvJr2YlF3o1nqImf22YE6W1AO/N3dSOoKaKVEXjTq5P0Hlx99PQ1LwdzlhqyxO
4+tiMEE6GuEZwefsY78A/WpSaqaRTeVbwH6LPbVLcoFQz0U16xhiBEc4qVTAtbUY
fpunnVVe4gvREJQ33zRoDg45/ruQmr3Xd+2WpiSge0uuKuuQxCsEYwnWWAjFQyYh
5hvEUI2/KyLFfpyLZno/3ShOF9Rc3QC616hZtxDaJgQJ5jL/QeCE+7YfrbXzUGg8
BdnmUnsoVMrdGAx4FkbX97o9sZHYEJo8SIfY+nOYcS+a4olwJhnpW4e9SKX18/dZ
Z/9jf7Rdc415dOTjcvoK3KM+S15qVMVmP6N53Vli3owibV1iVafF5Zn6OSISsI5F
zupkQK4DMBPyiX+pnmMIMXClERiYsm5Yv68Vm1xhf+nRk68m0h0HZmzVwRhBNhPY
xoaqBAIvgB0HlPMAs05Qt+Afszrcc9wIsWLc0PDqwShmR0enVZMBjdvCDsfU2pGw
zVpazw6yUte7wqrho56SRT4TtduDCUUqvcXY+c6WsJR+tD2j31t15qbUUgC78+bW
XhSFKUR2np96jUU5pGcwwDiHvSwzfM97v9S/j1NCu/lNfw7o3E8LJA8irweJwYMl
jm9tBC84QWnY8F5w4mvnqUOzPDwsfy7HO4qDqBu2wbRT3yzJ508l4/K25j/kjYTf
OcT+00RKGXj7F4TbYyxCBOv7Ki8NRqG8NmgSHxaeH0rHzVidmvb46BxlrOkj8R4B
2P/gGMz/xuskX3PATQovurRs/YlFqbYFD8swZz2oDW4VGuFm4hj7c0n+VPCtX5sr
jUkAgFAqbEzVRPl3DRyoIBAD7fqpVWVt0PyJasRSVCaMI/0qBALtjlWaDwaTH6Di
c7g03YDvTUzfvKm30PWrP7KO2EnysmxA43cj85zBoOCZY4D+wacQ7GaMv7yIqKEf
lDvgwt5lwtLtZ0+DJ2iZxIJkHeWNIXNdWR4NEAJG/KF32eIcFDY0nXC1n/1imKsj
XT/OXOGG1HHiWIIgqAxGesTarAurd5jN9WrhSvkWrH3ySOqAK1qfmhIcHVF8XpO4
5qh3pzOak5uxxt3pzLVVS+x+QqpqPaAQzUGMeAIb0uUHm27j3e1tJsJln3JPh8gr
wTSf/MUjx12AMB4gjHZl8C3MKLfzOhn4MAryCCx+v/KkFOJQy1veIhwhpFVF8ad1
+ANXRtDVT9rZn74aCsBwAui3Z/FoUFCs/CfRonBzaudU6CkQHWL07kCDJQvnVFYj
rEaCEDs5c8kuI9AUCEIt8s6I0wr6LbYTDlb+6y28Bu9S7Glo88T4gLxcQKTQ8xxv
+ICn1v/8kYgz8eCPrs1qcoVxKFyYS1IBjk0lcVxlV/kVuUUoyZ2aZkVP2hzvjPzw
15f81hcjV+duII8Te5PKEL38JDFDVvP01lhZFXKnxQzdchm1EIKuOiuU7NuA2nMv
Ub+Ui7fom+vnqknITmn6c2c6JGldxMItnJFbSA5d5u0gg/oI9fGZUnz2C9O/qRPH
Qyky2ElfkRF6fSs/+2xJZ9HwDdd7Yox101LV6cjPTZmw3HgnVnS9XZloC2Nut6Qo
kas9Xl356BzyP748a3ZljBYQvaxxpbRfrEzOdAWDTE9oKMJSqAgLyOsfUWw5+JRP
fnyhxfxFxFHF4FNqy1BMCc4xj6W1kJQ1QbNMMvxlFIQAvDD4gvr/3KRJnxw7nirL
n2MMC9l+7+yW5pviAhzeI6H/tKaIt75RYJoLG0eI5u3k+rAjoYzILKsFud9YpB8n
c+vEwf8kXFTzadzenLXCUTdxvhkNfpwsRUxLcZYE9Duyn3/9QnMKZQcBM/bdaU+K
dYM9dcj0HX5syMy0MnYLj02CWG6pxtQRRwYVb0JEMdRjamij5RgSveoqxyOO9j+3
kyg+A+lrHfCqvaKomHgSNl+a12fqV3axfovpe9EJVItQ4+ysfPozG9n3j4jk8Vly
9Px3ZMwXmniDNVS39pYG0/28kKWfgrlA18Obs/mRYO8/6D5z7OPqVEnaZQcaKCs2
tZrCv7nxcuiMuQkEEcadF/IHb17BJkoc5Xj6wG66FVPIFsXneIsl4y3ACvaOBwNE
7oIkcwb57tbkVEWhkYPfajoSj/QohCflV9HP8x5Dq4StB9WZnF18sMHECJvVWH4G
oZ0e50r9wJRdOHggsboBRkXgKol3NkUis34M4ex8bbaenruljKXZ5lZuRHiPkCWY
mYy/mtc6dGAJaf7xg6WQQMvfPYlQSzUEhSSDnQH2Nv7FP4dkdtmpg8dzBCJwMORB
HC4isOBHGww7FCge2V6XzGqkId+Q4iGaPGzmru4m3LZqjaNp4MHRX2bGFSRPlTjF
Vo1lMo2wj+QA+KRVB9WNgDQnO8mBUc+OIK+N3bo+gsJAb0vza+f42s6LAPSO7sbs
PvVVMlNeMVL2ZgWjAMMxInmFXw4/5wLDLp5BB2b5ymVDALG9LQCZcAmNqzFf7EER
AQDTWloC4p40EM5ngv1dfy+z1485L4CqX5bKLr4nvI/TAfMSHt6dC5oQW8D1WvBi
PkzO1Tz9uLINLZgMNLeLc864LZy636vaHBTnaNqnmdIckNq2MvqRgrvOUO+zmjAT
t6gMS7VU771kytMu+X2D1T8xCBKF1CFS78du4QygiaBS6YpaNyazKhnb1v97hp0q
uzx7bWpfjsCUL1y+krSpFZXgow/DUYUMjEJRKskMOt3Mz69f7IcYzhdVEkxu/j1t
LUNseo0WeML1YBDYqSbRD940p1mm5JRvU/M1gFm6lihIu3poPFSKYP2sdIvq7HFO
c6o+nrZ42HoODHiZvEzhOSFOxSS4CTOX1n3vdu1N5Jb8knB3DePo74oGkYAZcZEF
Ws5LriYTa6ynlYTPwCG8ENO9ft4N57PTHPexZy7zFl4e7iP6b0Qr6y0TunRS7EGd
tT6Ze/LYH10RGTu+Qp+9fwr8px29oWVt6M1a1h1SnvpNw6WSkl5dNwh6sAX65q2S
1WwSQYXyaoRlBugoM9lYzsyrfqIWOUXba+MJ+dXVvvW9hwIeXOTJGmzmB88R2TJL
jzbgJvH7GqFtpPowR8C560wQHRG9XUimEOczP41riImA/qJRz1lr04BWtdbzuFJ6
oD+nCQx3R3+Xi6EZWwbjrKHKhFoEFVyXuoVSra4xcCouJYe43dAt/5XkhtSXTIFX
gxjSE5DTlH+s13jI1dRqhlFBu1Uq8LGGj6HZ54r6GDKmyr0y4LMhmCdGB/iA6Dzz
etVBcGjgThp+68ph2CXGDT1jIhuyI5cSM26K4X3ipQ9UL4TjEXDw1AZfxUjz4KCz
JRmrt4zfg6vUmpj4B7y7yLqc8A+W52IgrDQ2GEIDdhF3gCD0QqID3giAvLWW0ouJ
6/HVlWVKFPJ1v8rArYuiKY5RUlca1gp6n8wIR3ii1Fx34qqzxp2k37IfLeFNzQ90
DQCA1H/w4S/H4NwOjE9taAIXqJ5GAvVxzuPgSsR4vRx8CSj++kBn3cNddkSVtkMw
aWazQKp1bAGxK/OT5cSRaR1b308rY7yafHRfzy11tSXhR7F5Qv65QQ9RTH8GeJFJ
RcutgH/oxtV2HgwFONZEk8FcEmpYx/HXtgid6mujnwil5IKmS+xNd33pVF2I/SGL
nSwEUdYPKLYr/H7mpnLHEZOV1fKdjy9QGmTup/NE7bRo+1HemYqL6p2wMjTWDs3x
YrtMn5vxETpSsFvIZgY1jgdLQJrhNSD84KucDQj/lf9IeR+jOVsNfJc+7P+zjkTv
JhYnFSUS7Iyran8+JAdth++PjuMmrn9eF6o90wTs7swXcDJMEU/g1onyFmHJ8jku
2mTxAj+D8y3OdoA6twM7XQiPY3fw1RcMyrgtlUtguRwWVBHSXNPtWWaYcAMuVz9K
e/bMCOrMlBxZnpTJtDFceoVq6knuWc8CECj+GINyyw5g+A7roACpL8RIVjY2g9Yx
+JQGacYTrnQ7Q3FLApUtNQNWeffpM7e2vfWRLo2kIgebVaRp+XaLc5C0qW7bPW+G
qvOPgnpt7La40VHPVx/c72UdEZuwZ5KnHFMmjHiI1fCRYzvE4kDVnZ7MvF7Q30Sn
YArYcUodOM89qIQuH8HMW9fNhIMhjVTJ5sHNYd3S/rJMxNO+10hYYMEysvzk1UAV
7oxl3RTxl3JI+z6QpSX8Yza/kzmjqiYEIKZvyHRD1u7BlzKerafiBGOx9D/BdEYB
jQOwHzzPRy7mrzPrgwM92ck6m9tPPjNfU8e/AXJwklhZDsEiFcSlWcaWqxjSS13V
6TeSOcYQAfJrhTcw2GqpXmIEX3G7YkPrYx5G2lB8X/tJVok1Fzj9OQOqgW/WcG5B
5QkYAQ9b/NjDPnvctq+dMgc4qLVqXXVggiMk9jAj9o7jYTueTBJDJzb/Z26PG+pp
ouIqMiHLbZvV3Ld9QNAx8yosgYMeqxAbpwyo0ZCPGIStqgjHPqzSY65WuASQ4wx2
QQqGDDHEBPvHmwfEKKrCCsS5cpm8jouQPJa5KTbGBdlIyywnlTxYvKupaY7j0lhC
rmFVTuAE24aq6vmC9XsilT3s3/b4BhYONiWK6bnU9y1e4iE5VGO9pMwNz/FerTQt
6+c+PmHlnZ8bx7hx02HND7g/yeoeXRaoJlv9QRLGhBQ+txOd/FQpUkJ9KN8AYV4a
hmxJ+zhPX0Io6V+qkV/LRcrp3K5iB3fRtyvyJqSJbN87qrdyJkbOLP4WplQ1lyyb
txADXDFVNtfm2bZG44AIb3duBEUh4PVxuA1GC//5Bnld0srHJyczKD5TU7uUEpoO
QyF4nYMkcPDEoWk1U6ZnUt0oatudeRFkGYmya39Z2BR3xY+Yz+LFuA/FFa5GlGQq
m8vbQkZsabmYi24ng6ucqnX+/Yvxzax/BR3Tr/IY6RVmx1CwA9/vD/67KKTaZ3iX
llGlz6e/z3EvQZmIveBcsp1fVAYzuHZLs+6HyAW6odxL3cu/ibnCK64oz3UbeVDS
7x55qBmZbEZCnvOXeQpIQZkyirCJVDvpQmQ8RSFi/GFmLPW7XQAehNKW8zltZdO/
VR/dytKppOQbv67+NRRpdB2ho1MyhRRyOZnoDKgo6EEeGDJlZfQvr1qrCGg1c61d
TvrgyiDXCEAwBGxwsk5P+OZ9rig4lXmoH/Li4mRSbQlA1xdNGpJSaWTGs9/fLkrj
X0vgVLsmBw3/hBsCAjlEAaAVJCjnJAN53w5Ig5xCnKPSd2HR2mBabDP0GpQ5m6qM
FNOw5BfeWizz1Z+mPoe7EQpeLJ6P9KvtVOFCFb0yO2JyqKIO/91ETwwUmHmjvM5j
9qpuAs9mrUOy32sxgcLivjP1/3SA7Qns0NHT9N9MCcolhYEfeHJMXuzqOXKiiRae
S5Kgm/VZsYQB5ScYwQGcJtfJCCUtWYok5CLephP9TEt4wltlsxfXxNFymn/rVoUO
bQdmxNtn0khLe1HTaHglpLRXuQyn+nKRx1mNNsyYq9I6DNyk3n6u1Lne8TpoMluw
a6JtgBPlQibH2EBHtKravYFUfM8PMo4jkQHxg5OLY85NN+znXmW2XxziUxbhrE5c
R4snESkanGAdekO9ceQKgUBDsquUnGfrPEkUwJux5gqzB1QzMjLpSW2YKUKRiRhB
kSJnZkpFgmF+1Ejbz0TkzxKe3JtrNdnqspwGg/j+Mp3tNZ/ZyEGy2mrNYsNt6l0E
V8wM4BKI2ThcuFdM3Pgx5dYh84V19DqnSJ24oGKZ59usZczlBYc9GPJqUfu0mdjp
WxFZZzktoHihKhPz/LIj7DSI1UzyhPfWUyVmWcWZbaqVz4sufbVb8mKPFyUO7tRh
444jmgvWzvIC8DAc650WDLfXp6mrJJdxOXxbMRmzxIRhTWDy/ZS4byeqt25cn5n7
LVNc34qQdLonMQr5WBdEr9/F7IxbyztwopA5Fvl86nQz1jEz1eFgpqkaxL9ewSps
6RpPcvl9n2YrSQrRdwBm+DbLHbWmNfQdyuKK+pe/Pos8yjSl7d6nv4Z99s1TiVYR
TZPZnMVSQh5UH+Q2Mp1eBu19B/2rGGovnGKvkFQlunlKvCZibkVvIy/EM29G8E41
u28JPuV1ouPnR+GsFgMwp47fkf/abOmRELz5ui6u2mcGS4G2oZT0ALrOek5KjWQ0
HVFkij3FdsgTJ7pxjFweC6Bxu3QZUC5LrXZDMNOVxghwTNpciWSZ+8iuXzNwzp+Q
eoyZ/9GfGy7Uo/C/2fOLVITtglxCMPKDD8OYcCUfD3Qt6aR8QRmgc49Fg4RiA/wI
aubgDO1wM4Y/hNQ00vkAe+r2HNhgEYuCAB2jdMszSQHhXhthFytKq8w+ignPnDGl
FJUOniZSdG672GR3XPX4PVn7+RNqPbVv/w8MnzCma1RxPr6uTM8HDm23A5eSRKlb
GYuOIxtdTHPjiQvCosOQxRe1Sg0SJO8TNQOR6RjAsZxDC0aMcX5dtEo5i/q1mLsf
BifZGUexnxuoSLrb4mskdIohQPJrgt35iGeba90SgSO99NJ+gFPptJOenVMqOcqQ
Ts3qe+ZkbZtgrDTHqegAjCP7K7ukUf49n+GZz5pKUUo/UPEgkiW8UWEXALDMCcxg
9PpAAJvlTcfYCkvdqtfKMquIKRjUNRwzcyT0uQJk67EEJYfNsyt3jHqYNGVHzKNJ
TyVFXYKE6+ix4aUJATZ3j/TIzFj0hLfLYZPZroOBwGXQ3CE2qVcIWpeSoMD4ppnC
vF4zEb5Fjyit8Hs35236a9HRpdeId+7bmaGAqZWbq9EEULR0qLW+Sk/0zzc1vjac
nutFGO4KvyTfQRNjRHhcOSDcvWhjlblVADIdJZWO5quJjSxOidH5dKMqITqyoYLJ
YOcbf15et1+22WBBNPBVHozTNEPIQPEb5xsuTpMq1n1OhcN3MLEj67bRY8RDtfOz
orIprgORh8/JsfHp1RGH1gGW+THDh6jKYhU1EHdraC1dGk/Kvtwxr0xGwI1uXmTt
bUqBuAe6N5A7hHZMVMCXbq/q2IAGcHd1LLNv7u3n+ZvXiME4at+6/cQ4uquBLwsP
UNrPhRUDswoFxYmni+Pp8V84eOVvZLE+F58pvpBG9rVjI3pjbS1ERNJ7k1inqFM7
Q6N3WHNHAdFOn0B99x5KMnRUydyKkoe6ffn1PRnDbHuVxhIxU4x17Fv5ekIHku8v
Hx4cOAm2SSGEPvDOuhKLCH5iwsMhJblWGFKsbQh4VzG/oHH3Sc5GHK80xAHWFb+c
4iJusJEKHnukRBnn6Li5ZUI6EFTPvNrIw2ph10UQg8HfUSCaLs+/vYI8Z0GFy6sQ
+jsMf9HtCqjbNRSEytysL/dsnKYf2C6ngz2NszAqgp8ZAGNoMSbu/oDMIFFchzBi
65QsnEfJpldH/+Jl5qJdB/skwJ7hIapx711EuFhVIMOlytbgiTLrFW4l5TwECnQS
aAfQGIc5laLKeNQhaRAKQgm1sKDfS22z60NkngvXQTBibBJ56laoCxkDshd2Pfe0
/ZCoBuw5lpXQouApo/yfNSOtw+7ZvCtgkEGxpcK/sH7ClikXJFV6BMh93AUgHfNG
tL4RUI6012q/96ATWZE4cx2gjR2rakPTumXkq29P0PCJwNzPEOj45Hb2OBwJtLga
zTNPlg8i+6T2B4NgkRcKHPWrUidhHf7ui5CgUNa0Nq0jht0431oH3tKlpqtCBT/5
+PFHDeQBBg23SDEOEkvz8PiYp4Uw9auTgs0UQyvxUO2rzOeZG+CVvSi42LiqLJDi
FvO1aIwHCyhkZ5LD5zxEScFNV17sQplHWWN05M3AeWZt2nbdJQcU4XPbK7b0or5b
3+fizUY5CGNGsJSB/28PbIouflfbns8rDE8NtvR56gr4gs2yl9ZkoPTr84PZ3VVj
OwHtIF9/2naRHZ7fo+HoXg9xZ9KilwRUbzzvVrnwKIGejei/KbYRwnGsX6mrChK9
27L3xqk+DsMu5fmpSbDUPC9qiXGFHO5r96yFEZFPbAEUx1arfx+y7z8SvQ3sQtJ3
PPwZlmCeDK+AR/pBdd8iC+A9Wmvh+4g2aef71qH7ZW8Gvw2IbmVvmuH65VvoGJEq
HcJGwarO0Te33P4ZM4urwPY4CWSOBN/Fp0K0Mfp3hOUpeg3oGsnXxNZByljeZhlE
RZFMrEAFCSyPT8kkcjWQlglzoanECwh6POzaUmzmb6Qp+SymazQXRKv3qNWWMj7/
TAunIw0ttuWdywbIkJXUaJRpIxrksK1XPE5UZinRL2t9gVpfovgLXHbrBB0JAlUZ
VCkadxLBiY26Ski4ayhSLfPoizoKYmI7VMR9IKLxv3ChVijvpw/Mt/FVUmSk7Rg/
pPqXQ/wkrP/havxhh2Eeq4eLtULIf+0ElCSvECnvD7wms3cD/Z2Asfv3Li7XFsv8
K9a44g2GVLjBSLzqCw91j1/AODMplY1bCJ/okDT6EHfDFB6/kYJUghs1NOZqqTSh
/4Ot+bTzENyqZs3hRg7IkiwzbbGeguwqGRnP28SRQdPPxWr2XlKrBm7t1YKmnssg
3VXo1RUQvkAFMg6qfs8YSB6NxF4JeLGv5bz10TyL/mMNZhl7jNvmE7QILnfsBIfj
zyq/CJGVi90wbL3xSDbcSJYBi+ohGOHS2eNgp+zrPTxAqmnv9ItAMvpBNmD0+WFA
CXFhhZaULm419Br7bl2yNqUQGG/1umYeA5KIS7UVMYflF4tp98Lx2CjO2c4eEjTw
jBxVBN7h5WXns5Z2ed+qMsT8iRknSaf9RCBWyIm9H991Up5HyMoa+nHGRoc1/bpm
sqzYPDFfec0Ai8HLzIUwIQ9t0Faq4xZY/bl6XjgxZuZk+AOiNob4x9ZdjB5/IjvX
WApJUBdTOQ6D971MZ+cWL0Ql7fCYtUZWX7pn6LFD1CAdeLjgAEsd1XDPVIia2jpk
1quz5wy8sD//arCJiuwEcmpHFXVD7bcw8SrG6JMXCEFusFAhqbtQWkulc5sPmURk
z+66v8yhXGG0CDhp1AOrMBf1fWJg4vGBF9FOHyGnlWPyLPtcCZXIZaLAGh9rzu2F
VA+CUEMDao0iCy9YpZmDfYvVCvvE32bJc+o3NIi74WgYtFZUfsQqxAhXatooyPd7
bK7D6yIzMRjw0fTaWjdgyYX2YCnfoBBR678Ncb3WHf9KOIKOysCXSklsZIkz9yqg
MrU3QwrNWOS52gcsmd2WtIn77S6ATblgYYvtgaMajAxUx+gmjYyE5un8ctN40fWm
dJoZxMr5BJsLpLQcAkxh/Kxiu93ie1aGjyBVbRzmMU1HOuSG7FasYEA9hm8qAccN
adL0N3wRQ7ee29qNUfaboTNbEOH50737a1/6EXY2e0y2l9KCWHlcqMQPCCQPak7F
OimUsxdglTmslnSwu4+1HVHUY38WIcT1dbsAK7Obg/64H3BFN175inWCLHrRy/lc
Ji1BhV+l92Sbv5Kr8bSA/Oc6oxPXJGbjawsCXAbGuPvy4cx+otzJSlAgvE43hotY
A7GHTdhKxWnaWLfJekI6bjhexvvlABGGoOpkh7KqkCe0XDFSarp6k54m/1DiHLfh
IYtIAywYz999SVXPNCfKqZpTZwWkUL577w54JUBMOOeD9II0vXe30UzXvTDFXdmG
pUMH4OnhzEeVhIu5RBUf9szPKN6wDJ79vxGSZ7BaWnf1zl7gK7fOC5fifx03EA+6
JKpDlQxDk3B/rdGCYOGv5oU1WZqR4aKCzM5QP9Jd3zJNw5JoRqqxK1toQymLj+fQ
AQ+k4yi2UWo6AszDQNiQFpJfJmZZxxRmheqqZb/pMac9IfJ3uB2eoHo5X1FZV0IE
Lr6DC2XikwYA+vlR9aQzLNoo0ul8QMPSm/tA2JZa6/CTKAFLJQ1DmIgQVVpr0TnM
hQAo41wo8SNHa8D5eA2NCmW/GfQkuzGP6rHWQT/726FsdWtOzxavApzejnZ444b2
xrjUMaZqbsl0UzH9shfH2LVKU45166f0v2upF+Ixz7cwG+cFPIOrblSc8uTpp4ur
KrS38xHtZWNy+c/4CrPfrJ8+PVciCmcpr24dgP+cP6XbNL5z+i63o3DRifa0ujnr
x/5sQM1X1F/R+aMARIo0zcU1ZnRSET6pByFP+tWc8HdmfWeX0U0EPY/EyY9ocA/J
l/Y4LrsHkxObrYEz13pRBxM+wseFd4YuGsYP00Nre34zHc51Dvj9V3UzVv66jUnP
qHhJH3eVlKoWjwKaRVhpQU42n2mc0AN+DSIZKCkKgw2OzHUF4JWybtmFG5ObHFGF
p0JIrUWyRYxTwcTAke/5e2PhOpNQRMhGVtoQ/ZBVAiT+Q+ZGEZRyiX1AQHIorMEU
fTu1W4l+7aFKmM2uysS7yO6U7/mpz0goAO0Y1yOxDgqm0Z7IN3Pvawk2QTsBBNT3
gVxgDrpxhAOX0wNhUBsYSYyzd00TMBArdzRdVS85FvfkbxNt8XMZ1qKfbPoljA6S
cbAjF0/g21Vj0oK/NkmRSUm9h9zD4KujeVcTDXiTUMFB0SB8bldGCa9xmuZZJY5x
/q8EF2KFFiNWvv3ivm1UOsCSTiVThBfSqcHO5z9MIaNstimX+PvWXuSCCsUlQ8Lj
34I1+zBoZnt8OteXLZqPod7mAAUCPo/6gnte6VckVN/xX5isZov8sZTh31OapWDH
pOIQra5DTKBHxkj9Y7Tv1nNmYLMtNylzMfIGnF+neq+tUMP3p6CfXgYRHniMpMq5
DQlVs7JcaWqX8J0DYBJ6Dl7U0HpuWAI/n1jyBt+9OD2y9BqTa2h7J1p551b3fcyM
giCCR6hyx+NqXYciO3Kc3mwT33oUdtLpW2AgXMxXJ4lNbag6DNQpVVHNGxmkaLYO
qehEjmUYixoYOx+4T6YNCVHyPmTfuiSEpRhkmVNpL9VPF0DiEO4XMRL6pVFTceTV
r8Psbbl4NwNWCkI30HfjpKAcgCTQQy8oHWGMOpshK7OYB6ULvNRjAOyZ9NieFfBc
OY9KFXpuYWiq74bixpg+hjc+2GZSkxjzLgqCN2NhB5N0pkcfWe69QDy6HXyAQ/eg
gntI5727ch8KAtqB/04o3vUTIw49ur11Ruo1zVpF7li7/eBVy9UYMB62yrjxoRbe
bIVg1BPPtRHLUdHUuJJKN37H1uzkPwIAD/l4dxC0hnIumvCes64hCoHp/PzbR1ri
D8pou4MXApL+v0INx7gqcVD1Sfvf8gN40Fd/DgJBXC3wtKJCTEgaiGyR4fiYXE2V
0t779nbpPWr8+zlZGPjBqpU1WhsvD4HrY/PZfTZKPM6DuRYlAj69tzduxb1ab4WY
QGsVyR5n3oEPIzS94Mzk1VH7EkhP6yWWHxkd34um7bK4QrDkfquzWxpePFfX4Yje
Hb2cJ1QLDx9MSs2mW1jvjdwEoNnYgBhtmlZwkrZlhsCrWvCe4s1/LCrdaI7aQW3w
iIfSmFo4k6h7vINSPZAfWCxy9lrO8TMHHkreE/4YUgFUCoVT8XRa/+DJI06IyzWx
eeUOcQCWdaH66aynjWwzBKE1Oluw7sspQIjYJZj76sQC+cBMXvLW9nCckYps77UE
zkcvemS33M1PXi0K+LLjAReSX+jJzz6YKu8FIjyqzZ/QxLzD3sxY28alx9eV3isq
AlD25JNheM6xp4o+V43jv7qgS1YKhXYZYi3ZtzKFhyVkvRumgbY8xxLKaa7PHSpZ
PiaOaXM7r/Flt61XrwDrU8M0vDUJ8w+RRFn+YZ9gzrZqZakYNSTcoOPCtxrO6kZq
1p6jreN3FfRUgklhC2GdTYqvfN/O2KukqkyOWuHyOrt0fMtfcldPl7KS+8v/au+a
Gf8a2bgG0B07OoJghg4D5npq4fQPRu4/ij84kwe3ZoXvGwMvXQqSZVlMmv/LKDOo
pv0hlaYUsCag0BF0Mu81XUczyLMBrIRYJ+xDCWZs70n07TMg1CZ1EmJJh+Rxc7Ks
4oK3t3AKinkTAbciqb04+Nj0Lzun/EUGdp+BPxrKo8id7J9NA1kQz1rmou5nrt+7
/tec6TW0qjIV5mIt3YZ+kLCE5Rw0A0NoctACf8Wj/XBezZLuKG3/8laEF1bPoxLo
C3Uif4AjP8oxhumrDI240+YNcmBIyNLhzQRfPZFPBaLSz5l+UhBFa1nuF60Vtpyl
nL83OeGgZ3uthwSTi0bUl4rJZ2OUcUzj8+eAy/Rn/ox5m5F2yxuyfNzGmEwNjXsK
Iuwsmpyqt2bbYgAIjH8kLnEizF332bYE1iIGUEPveRwZLOYNmftGHsD3HIZhXi7q
3KB+b8DgVlXDbY8NccJFyYOVshVBB/isvwRtoYn1EpWi0t5rRJuH28pqYu3jXOoz
962XQh/RE6h8Jec7J6fLNwTEyKOV6q3Eoc5CEJMMC3qHMtRPJxQ/KTCH3qD/b8AR
oqSGTNVdhmNxUVw6R8mabYCKPCda+vgl6joVxPFCli4yiKMKTiVf4YPUoemYNdjj
QpkANNXQqghzZV2dq9I31iaQjGTtxNpBhwggI2ul94vAX0ikfJ2N2L3qo37BhXWa
iyRwSpKxJoCfMfrcVXKJCq1X4353E/4VH0pbgt6ybFmqu6VdaVukoyn9Xat4oN25
QnaygQLeYxr92jzn/4KbBFTiEMNNYGpNq1YJhigkmIXGT+NjHrwcWUnuOCu0syjM
KqekxPGvU7G0TXnnGc4tToWs4Z3kNblFeU7vI1+WNbSnhJpRsUKX8puIsWRY9XWw
R0Hg/Vhny7H2gwOvx5sYm5tKPGP+bFwd2RehK4FUrNxtEmOxzODJ91yFDGkZ0XGf
7DzmU7G+4JEWRAz1tyUxxiiUYmIFMe5G8d050VEh1zVA/Xv8sqKTVfpRR2MsYTnI
S6f/Jgg32LCP/B18TrSnzJCB8Cab3nARBd9HAgFY2TYq8KuG2YYz6o8mhaNgqv72
PzEv+XmYubUr1XO6Q3R4o182Nt68YbZIiOc2TLaHWz8zE/Q8K0cPAybd2408e8Cq
Aag28rChLlhokjVCAATxGug0uiquM6pG9g2YpA1GXmaQ5udOF/qBbDUidez9wbuP
/vjdfofhiEJwxNEJxY229CZmeThftYHqMmroKtiRCq/RQ6rFI6w/jQF/jMmdPs7k
ZS5TbW4PxdbVdr4cXU0rH98/8+tR4tM9jYJS29dD5IiZjMqiEAFYGXg0pZJp2dRC
8Js0MA3MDFc0ClrC3F2I3dfUraG7uzmRlvhs3rICXVyil4Ot147v/VBrd5TdVaJc
hVBYcsPzL/kdBvtUqXfy8NGkFmfr0Bzg7oSM4v0PtWTbfPm44vwXJsCWx6BTYPRO
Bz0H39k2UzWfLmpaTwwmssmbEbFtvJzJ0/iVe5ISXll69CmR78/tyhzGr/D4O6wP
PS74GOw/DN2R8c7LUP9CEKK++1pWIAZeL56EYu+4tmmVT4EZtyagFJG+DhUxI6GV
qnUmgyl4qh4moLuZcC7+2RKrUGnFFbsJd2B6qeqU43d7rqO83ptkP1rzBsEC+zsV
8ZFyqtg2YX2Lzev5h5wJiPWXyYyJ+ExDK/c4ZAYp88euKQfXWxHsrmmrslaegaLF
L5NKKmYGNMIkwKTq4DF6DJXQg5aQzNGuf3MKyrwz7sWEh76bbCia1je3WraJYkvE
hGdw0clqFx5UiqCg70PdRiq3vowqqaN8UtJw+SHEbNTzpRLg1v1ffRUs0t52CsRf
GekRymkj7HoAAunPwlks+RxoAlOi1jAqSC2VnbwfWc30I52EqI7tEEkVvKdf1hGP
7vhIBYOuU0Py3NNA7NYbGVidW8OMRfWGxvkVRuz8WMVDBmx8Hwkpv6U14kwLAm5M
QKRjph9HArILa/QSzd9mHpTwXuZiYwO8Oxrw/loYHU56BV46PIEzXKdPRi621rJ3
mrLz1VWOaP/4IT0TxcDCUpzsdAfuLTbLCWIpGTVGYGzeyGXx+DwAJagHixWobzYj
8zolWy6szmXwZfTpq5ZD3B+8ztNqNAS7kKt9tKZ+Oc7y6F/m64O0Ku+2Z9MKgPri
ggLQ2irOvro8ZSje78WiN1mZiENBPCzSuTGeIocPJHDm46YLSKYURz+UejQ67n+m
HolNZZqdW5+Q4vLkSZpwjIEVXy0pcbnGQvhnlgze35WlfdZnnRUNEDOomHAFkrin
fQmyn5+hebk9f+WXvLtGjwHPUQhNnRicLcHZg0KhqN7BnoEgohzGrFpfi1hBtXBF
vGAjORBH1TBwy3J3E8PgPf4ykUUr3eVk8gAuhHpKml5nf7UfeLLy8zuoGspfz6O+
P2wMj+Hg+iANx26nH9LzRt0k6a6kwqx93KEy4pnAsTz705cK0o61RZcPCmmvIyri
yaZDn8HqNKR3Awsn67cWg90zfkWkAYoa8AGZNmu7tjEotp5wi+VreNSLXIeGcWl2
z7R2NdasJ/UXtNGpby2a/Y+QEACCnWZW/MhxpH7Fjkf8BVsr16mEuTkDqZhZ0pMq
P8IM8EKIO3U62Wx1t0Fu+lKK2cwoUwRMw6TKFs2lLHXnydRMLCvP+L3YMJHPMBTd
PrwIWP4hoCcrBay4YGRO+Fxyh1cEPcCpOlOT+B66+XL4ezCzqwHKqOU8dACshuTO
RJg6GBWlDKH+0v/yYTMLZfVfO/CyEWYWIy81RYEYTP4tAD6JC6Iw5tyg8ZKKush/
Yp95FJAEfqgy3D1vGmYr00sUqnWcTpldjjJUZ+bXVhdAHeVoOKb/WVJMmXPrmZf8
RUWk7pgeHccsPg3D4Ro4E3M2rUSfY4KvQeWA3yqTD43BlhSfnTwTw9P4N5PZPflS
fIFhECWOeuv2Bz1C8PL+LfZSpKHplKH11z5Rj5UGP+VS9JcAFMWEP5WRAg35gcPR
5Ma4q8vQDs2kXmpGVif5fXg6e+gj7r95Eh0Ix8MlTO6w/9Obe7cqVorcddb8tiJY
3UNwRNNCqfsIqw/+78/7NDIdmAQXJFqM+dZ6X/kGcYDiLMG/6t7o1qsHUbdFKyiW
tgk3daKonHHfZBOm4G4DoWZBcVrkqzWXGV5BOxzIgYlZe05atqXpWR14IRxmPSDa
j97VyysStGLIOhsRAEyETPoGCKeYKypCgu+nAp7KI10gWaZ3F5GFxu9/xq0ESyqw
YFLVn4oJhum+VcwVO96dDCrqQMyIpaZEjMuersg77CjuIL9IlEow3nRmzHlINilN
J4e2kQVVD35U6qQAdibt04FihV00jXQlZAsxgS+B9zEbxRf82YxpQhOip9ETeImT
W433E9fEpTy7QqgXixi31LvQM9LlKmD2yjbIgKt7x4lxJtrF91PbQqqZHsbLUY8S
eanhOL7uZxPnpBtIsgdFSjtKbScRMGDxls3E85Mll9X6lZr8QXthr8xokcffQybT
IvIWEc6ryi/j0613+5zQRQdQMhRs1qDGp4zG995xhCmUm+WcIrvBEtlmMbxolpJ2
SQMsCoAK5DblKWHFZ1Wf41O3OlWlgb1ca/Ftu/QTeacDwYMaUEyhMcuUwFVLrfIi
FamXsR6u/w/a0GvEfbc0FH1Y1F4A6fzYsEPOBa+DPtqsGeU7ekn/LObvbl/meF6u
8vBPFRpl424BTh9QaHrUzpzo2fIvTf3dfGCj1IHCYPOtm6lFa8/vFL7YzGlYVDdo
McERMau/2nm4uebKcLuB08wxc7y1KpajvC3anjUF0N5RUzrefZTmMtyiWVJduxL2
ADqZre8ZAeKTdKOKTqBd6L+++VKmXzkApc4an99swuy0he3hh3KgPcYZYEc/7ttN
+/WYyv61RmQSGG2x94yeZaOXGWL3zyzddZH/hOI0ea+skIZXjqimkFjlAbqGwl8K
HoRA9GcSmapFKJKu/7R6KU7ksNOxdkHC2P9jrye/Mme01uAbgJTHXwODI6ebrGVX
hbExErLw7Lt3inzwQfQhXFAYfGpHdJG4wJSVJxMt5jqHYbDTgaho/bZyc8NaWQBK
49WX4rD3FuB9NGKvGeLoQKfHTHFOVb9EQVqHKlTHAKmsVd+OgzdXJyy5Loas8KdI
sFXzftr07x5t2eP3U6Xj2FAcGoafCAZBTXwKFt1mdar4EEOdtLg9vTvZD88sPCJm
LbiWhdYNixn660Q8H5VDw9GX/Whl354eEM+Lck+7g1r3f17Ro4nzugvds6ZDTxCP
BTOQCT8LFPn3ZZFZDaTrGyDKBIQ90IEvdvWhnloUpJpTGsu0IwW4nU1R9ZdM9joM
dqTNkL5xRO6wxYXm25cepe2mWl0/NZi6/ntfZxNdjQ7pvdUuBT1P6cDSH4REo5Gq
/OOaogLqvyOHCiRmww+LjgiXaDKhpgm+Z7tzMPESbX2t5dDUgiZcwAWsiBSUuePs
4/CRYwWdWcuiAZvabSy4Toc1EKNvkai0ZP9AmZKShwJIyeL4y2xU+a5zPwTFYunz
vWlUYRJSCpVCDGLl+C5M5QMOSnvylcM9hbkZEbXZpne9EMRTtIA2JN1IgtdM0q+M
qsDlHQIW88FKe20/Hm6Ret6hWzuMD+xldBgGoxWTg8J2SAoBSf8ucFm8BGRy0Wvv
u+uMZ3eB+7zkULcqYwwhh2JpIH6bpRwhOzcGDoE0CpeVyqk9sLF7G55XshJSfBfK
3ylKkLprHBjACksx9M/78lqdSGIsfkTiFhVCqzWEPuoSf2KKAo9j1YAVIbqWMFv7
CJnYobbIVu/TxO8pwmFA4APvO2SuYPN7MLpgb62A74fr+mQBFifQrSf8G9QF8y0S
5rBHq6CMXfe8PTgsq4AwR02yz7ogNpO2ZAvKDmEz8xqp1eognV9HNR+GbmNHHRqN
0m13jdg7hQyM5zcbLR1acrsWQ2Z5Zn7mU+wswpo7I3cZE8n31UOL2RYpeYlqCk9w
Eh4l3jLm1i78+Tyb/qg5Yx7uMqkJqLfvnwp13pqEDJqROpp7hMjstJ4F9YXc0Huy
V8kEt/6jPu/N8zmZXyy6cZcLQhR3C7tRPs5+y3Svg3oBHKxTAafiyKGLCpapsLbD
Jwli2lVM84GvSf9SVG5LUTT1EygecebqrsQF8Moy4Pi5Y385OvAqr0Bqo9OVOKgu
VMfYu0rOsK5OvzaK4BTPnL0vYK8v5iE1NSVchdK5z7Oq8fl43TeqP8/V+mpWySi5
HYo7m1Er5Fv0qLNnQlWscttUzZqkuVdGJl28J/xtZjERDCHQs2qe4Uea19GjK6Cx
QVKcnztCR28qUQ74h0HPoSJjOEJRkQBBzJasQ5ullmFmJbUAPzEHsOx7qlrwlz+F
jspgte4mzVYKrIZTGssiyxL4iYY35We8l61HQ4tmaI02VutoNN2i2N6l2FHbq6oO
ks6VL9m5Rwkz9dLbJYQ+aS/ZuiNaVbMr5WlYWFAFLTK9FoG+ohS6oajijAmjLVWz
rrVT7fqAqj0LevIFe6SCHS52b+rgEvXgPWPACLnbQd7etfEOdG08wfOS5UjNPXSs
kfzlBqmUgp/beGgWhqXBmbCkXuyCp4eZSf7fnUCJnkN2HzH1iG93SqvhhqulExAT
EsuWh4/2xJpJUsx/Pd4zxnMoDHrwkAx6ty/uBoCkWjqeSePgneNkrwk4zV4P0r+1
XxQL7WADBpWv/eLI8+4MQn4k9sdeJo+/10GP9PgAyleg2muhSP2UmG7POdKvKfPX
S6vNLBPQid5e+9h21iRGZ1MygafiRBVgWhm1I4U4TGs/N3CcS0gQkEWefncyrM9M
hZwtdtqKmQIIh5FMn4rwS2aso/jH9QIkxyF7cw9o8gOdMQuKdKsmOZLiwQ3E64LC
uqp/KF7oBmi5a+Cff+ZMVVocSYsrt4XpbYrvSD24aBxE2ceXYTJ6WvnW3o1x5VeZ
8LxToKDrVm2ioDQcrWOe8gTAWHh+KfRJh0CI69l53Wxm8YcKjyFUNKA0Nzkr5pNv
mLJZSBaTuaCpP0rvL1n0MlB8W0axhmdWvjujyqqjbosO3ZpRv4dAGD9sjpN7zj7R
PL+Sg620fcqkIg1GTU5Vo5XbzFXWkstbDF4KUxe1ov9y7oC+zGZtjzBs50OSJBk1
VolXn2Z7/A1EZoLuBw2kcAiZRwfG2kEb1mYbuOuO0mrrIZP8zBkTAz6EDE1RPHHD
VONlRl9OLpaaWUUY2bxzmjgkxdscMNYiH3NjiOTxkElIWzyXqDDo6amMqDjjbo2z
k2ZMYvEs1EeA1XTgMtZpIpYQxyxIfjEzb1TgGbLRdzu8nZJQHqj3Vicjksnuwm8d
CA15VTfWzzthgfNHjG2988frp/MGfDaBS47rPpWM0w9P1umeknxQKlXNP/+xN1rp
CAghp6+hsUDD2D30zb79iYJlQWaboBjZ0ZtmJd5CAOK7zwGPBZePnD+xJceaGxpn
g1SwJKoDhqNdXCFL7TQahmN8C6YHVWLfEDeN8MqujqXLZKG9m9O7ANL+fPiV4hXI
1XuKEVWC1784y6OPqDl4qaHQSvoznjr/LEL991ejKcf4g56IgIlbq//ceDsej1x4
P29tBKOnDuM3qWrFA7geMGfPkSW69kMEiPSQ/PnXS3DeVp7DDzUfN//XxfI52Mf4
feHN9qU/bbcrVVSn0rwm1DENVR7S8akOpr5iyR+wDzvnNKrfX2/SAuIfvjpaTGJW
iTB6VkgJVcv9+qo66N7TWXf/YLRzLHiKam/0COZenqtM34uYwQ8BPSwRXgVEQerh
FS9cw5tF4WjMJGfMk/ooT0aqn2e6XPgdHh4FfMyZqRebPadnLyvj85kY3ODsI8NS
e0dFkko+mtxVpUH+REZdt4Tl/R6Rp3mEi0bFZTne2QIWcBhsG+CDX8L15NgLgMfH
ArnZnscjR3hReRdGZ+78x0Y9gtVzzCUM7zmKeLgdmMTcbkD295EcMGeFzOvNCpkj
oXasV1+8AgbWW/X3GGjPagVtvti/g/GehvOl1QR78DDbjTgdWOwdTkV4JasZGdQR
11Ck4qQgVoR42fuiG22NSPkts4loJieAtgvu2TeT4lUUKa5TVFRJSAg+23PFdZrh
k00jpg9iyCjhFDgswZiiZnInw7LUCys35MFWA+h7f/tGxpNKewSgKhKF/WZ6bBC3
DNW0Z3gCj0gG3av/bStk1z9CKhBt9ZJHHHl5XwwYW7JpyiFqTR5vgI9Bgpgllpd7
LFkKGOO/mTXOPiAc7FZFmVLuXEAfj8Nons0uVbUso7BZXUmk1p0CwgtXP9fjrbHh
Et2UmT9WWuAjNSDdSzm04zVJKgd10FuwV/IctTB8u4ipBj4kUjlL1qB9qP/Jzsn+
VLKQZys9miAQOhz3otlp66ixHBWmJy3MtW+9PfksVhEZ1x5V1UgRMZD2Xdnrl37t
/xGadAW5a2d71QnlCde3oKUafkvH8dIIZN+zY2tKE2ToP++xjT8v6IN4wctNs5XA
mEk5hNqN2VZfe4DqRF1FTLOIiXrL1ooovr/idSOdfbU7nFQgAQowLcF3r/i7d9NI
2XezsxNtEZGfOtOJGH4y3JreHPD3f5oqKjj4hgPKgH9WegAI6YdG7ibn0d46NmTU
C48R8MaC2sXXz265SA8XD/ZCclVDzIRd4MtcYQ1X0BCQlTYMblRZEewp18MhaXrN
4axZSuu/kJBdzo0wcdyVTptvr8o2mePR6V4NhbCNbcPDrvzxciCRGwO0J7oVWOhg
6QGSK61bBUrHSk1UXsD9moAJ4eb76qic462Kj+5kxI6ohv3p9jMi4Xb0FwSdpzYl
GGqgYhCt5V+yH996BTfymaTWEIWbwjLCIyrTQiZxVuGM7ey4wVGBM9/2ETKr7m7Y
+cqrX7t3WA4DfbSIloBYAwgDsPGxxIiYbgwBqJ3Csl70gFZod3eEY0Nw0+SXewIh
ErGcXhLWM5aJRnbLpOdcGiTqiVL7thQ59J73Ctzr6xX6LDFBHOxFKdOvv2KwaJ2G
V4olOSl9r36mSIKSiFqLMP6tQv63fg4UsTx88gyulceWKsUrHmYdYYaqOTjPUYRM
4XTBAmq71XiHsbOo3ZkSKgcy13OGkrm3b2i048IBazmxSe0YhHeQNtVm3wHaWgF7
AyRLVltJQkGdEAd/KtDCDnIM4T52dOP4BQnTMEW92oQ1pl/Lxo7dt8+DS2c/kMnk
jRYGVpH7/UogBRM0ukUoOi6LCYrMXdkK9DiDnOpRdXMoZlp0+rTWHQxp4it67K1w
2yoyh3FWjHAbdcKQczeCa/CNGPjt2JTdWsKgq+bxtC/rnNqFmWokm3p6oX3ymCXm
CIRaerpFeJkVaH3xebdu8Kwr9XmqTyCRsqGOER7YWB95bjTQv03Z/4Oj1dWJ6T9z
ht9npuklR/LdewKMcMWbQOHQtp152dhHiloeyvfXwl7fBUVk36BwNTVHlKjTrExO
mXGk02sRbWCl46JLWIhOGrZPS6Fgw10qR/H7WqhgiCsOwNyiZ93fLRjgz1v4dZI+
rMLylPs0k/2Z+cGASCAT5AxTdYC2rEZn/BwqRkAoXonsL2/0PCYj4uB9pfXkyRDY
E19Wmb9QpZMFkVH24NxNmPCy6uYHefOkj6EukGtqRWCskPY5QGIi1/WFo865tqJ7
yGVXgZ8cR2UrBZE4kTIZvsOdSsO+PwFjrAlw2HorVZ3ZWJmljGOQr5RSCWfGOkPU
u44IGo/zTu4cXzHxVXrzJI7FRTtMc5ffAfjq+XQoamc6Je/Ss76fz5RLl9nVp9S+
TPtn0V3q40WvN5y6W4m1vqz+46aFQ+2Ez5mT8IsIImbu/Z43wbTW4u+IfhLAWF70
Gk4YaMdIl7siKmKqf974QS2rJmoiH8Sn+Cx3BQ+4c/gjirUw3B4exfpnpYeu2vVi
cC/gSZ8N3eFnXhGB83M44/5cRYSGX27EnOa33NWnJvxwZzsqaOixTntdkb8VxQWA
9pUyaAfB5gSBZdCjkp8iyI08UbOztCoqdi/Z1YfQrl1TY7TEawhGy4WOJd/Y7IAd
XIFkG6nfiOXo9jWmajj+k4uGp3jqhnoeTNUXkI/e7bn0cyz9rz2crhEOsdheYCrU
jZ34m6Q/Ll94ig9GjwPDb4qBSOOqsAbo5HylbtIJV22+0DJrXIIyJzGHx2XPjacc
T9RzooQBe8+fE+jY3ZdOR7nldaI4GvCbC6pIKCcbLEHksfQa+luMZxmMyzffqAeD
dCsifnpl59pk/ic12iqJs5TfHjHcAL8f9t9pkXLeddvtPFnVuONIF3lVL7eLlY0J
M+/jaB5gVptT9sEbPcLvHPAVY0yjr1ctCcQcKLH7inCm2EtG88deSa7W4is8XYm7
cdgn/AhS0jgW7mluIyGPB97ZtPoeT+mZvBwlKtGxAHqOBadD8S66GEdFQ39SEwbv
d6AjkaKSckzIIIKk1fgr0FuznFFTbH0pR0gm0EYLFMrQ7qQ8TKJZsntt71F+pSNS
5vORISJEWUOf31uV8Y5f8J72HKxK9qEvPO0kX+SZPR2HHCIaNJupAKtrMB1fNa8A
O9lp2K3vBuLy40HxNA6qy4vdqL1RSSgV8FPotPy/NJHCqV9vYEXdQrJ6ZNfbvuZk
YNLzaF2Brm2w8XOX1dEGUJ4xbDX7Wsoo/w8WvidjTKOszXXIINRewQfSrpIPIhUM
DlXkuQi56vo+xkv+XUdRdY046tD7SqJrMBvfdUuceNsAy+yl+oPa09Ez8oqTNzqg
dx4tL0Xs+VR7W7byJzMBhCiAlhx6D9lEGUjEdZWRKQEUr6aoAaubTBC/PQ/yIdIp
paTl+ZgRe+sVVazZFHwRI0LWOIFE0v6/yS7tR+rfK2cn+WghixTlGnOf+sVDJnMe
G07QmmJDccCNDwHpWhPTm/E9r/1Op6oTTuDvY3PO3zm7WDhR6M7l+zA9Gb8K+i5x
RVQV9lJnvo0nIaC5UQSmU9a3xndZ8UXtUc/2Eif9ar19ZFGnODuPbmCqXQcmk6tj
w9yEynnj1x34xwRDvEkkuoG0+8Jfj42kAhfsmpJGV1UaUUwnwlF5nbpUzJB2JNwC
YGKTXfwDiXybgs0gM8xxAhGUDrTvNuFAXlSpIh3S1shVWPt+ZOlwYalSiXCB8tof
+IJyhT3l7umnOE6dWAiWgowCUOM8U17ZW0d2r8ttxiXWT9B4XoHcWjwEhDBiYc7p
DUlGPqimnZMX9AwB2ZUvBxlLhUAI0xn3e00TLPbWvCdaNoB2wFs5NuX2cQpNfSeN
klejjU/VxPfIq54zzLuhETjBr+N+tx8UJujtiLEiX5HWKuBZ4SGfdyU+84wplh48
mn5faljL30t6bVJg2zDwIOy3SFupPH14cG+hdT64eh2UqOLE3LVrvVzKkvwhcIMR
rgVm+p+8Q1QN8Am1kveZRhZ/f/EiGNMXOPO8EeYU9IWg4LlmQJUyJflLTUnKvTV9
HdkrP0DcGFyb75QT/uT487r5UXyENoP9amNkR93ZE6rg0O+P1UEW3LcXkj6vo4Mx
TSbIqMoqk9FaCf4mEGIaHSjQaXukyMFDKdFXgnbdZPKb7+RSCUYlDqdEr20DWDr8
TsVeR5F4D4h2c7Es9AJdccPSfftId5PVJkWG67qfEMFlagFcPWxZ4V0fqiesiH1Y
/QhnTZwIxJIZdDKA7Uuf/4iyTGsT+NlOFzqy/TyvyK173eVgyLBWipottMGKMRZ4
RBTTqU6j0Q1FUCeg0KTcLyEFuGDO/42/SpebHBokyA4HWdF0aZxpguAlcgV6omML
99wLMYKCe7XsMSaXyAGBhkeZW3zXsloBCBZHIqbKDB19wPeSe6AOgFo+8yWWvns8
EpsX1xGPsXvREhZ1/TrLfYhV1Cc6EzmwW0fWvuk5aysORm53RV7/o926cvKJ2Nkn
UyGAIasg0q6fI/2JmLMX1Qt9zReK2NGYhMO5IbuIihCEMjYKTt/eEEjEeDFC9hpc
FxIsK/07QmA284RfX+CgJtnpOTKOIpNwmSxgprHGLAAWxAGFfm5swJfyg+9DP9h0
N8LtkTHtc++JIJ1hh/5U5iys3THOwUUUUUSpwXDRcBUDg6gbaj5lft5CGkOjkv57
04gkbfzxRAeaepJjhd/68SoyKIuITLawmgIEXVrSANNHza+1hxwbTptWWt88Juy/
Oo0xtIVIP3Yvb1FP9d2hGBlRbln1nqeDVrNt/Vf09TIJuBfCUuLpfPD3vbSmXA0q
RqPKOj1bUC7lg+Mag1s7dn5pB5tHnLsF8wpmDaYGO0TIWdNXtBIt0NWQnjrNuigw
ucV+0prbKeJorVSwpKeVsMrDUh/T6x+AjUopYPUcgLJ7Eiu6veY5p0FjzpTuVi6U
1vvLtrTisVKLnuwRDN+GOWlDOuCLHSY2Ex1CLLhdPz7d3T9NKdkebz/6vZkH9/md
dxZXgJK4yADjzwwo6DPj/stUCwHdUzVondElHaGRq/AmdJRwh4JLIUyaeLnENArB
VK+neB338qflzVPwkNm3gzIHRGA2Rbdo9w8nGfU1or1zyVosBxkZZDOmk6qCbYk8
zw3jLxpMCsOe2x3XR5c3iflK+Re0JFEgDy4UqItcXk7bOnvTi0K7Pghc/cJq9Vuw
MLzXdbcmVIRt0R/qQy73Juq+0IXaEmdT78teN0fhX3QYemCb0WOixoc5BKuC7z6A
Roy45ay89jI4ktPMSdM2Z00if+dxGqNmyCH9YdhDaME7wv14vwn7o2yZAsKI7uwI
8JdoGYG2I/gT02wuFerDHDNkSXz0Xgg5Cq3CfPTiLG7gQUE2VMmrjSIGpUxdoPv6
bBzCgpv7d5I3BJ9UIy9YsQ8QZYH6MkV2rUuPfJjdd06UAyAuecy5MvVnu6XVq4qw
6nX0/YnH+LfE8+0cHr7fNdHxeL5VqmQ4o4cVVGjW7/8bEPgXrWUYPGHeF7e0e62O
TqMEPF57OHGpnKD2X3RAi2pgfHTfG6u0XzLwyKwP0KCtgfebdt1HfF2syFjs4Hgh
px/tB7ZHgbdQlhxM7HZXefFEu1y9Mla9fkF6+WmsGLtx6yQS/LzdrEqROWvmuXTt
JBUO4Wo+kCBMmS9B+xpinfI57Ec5B1TF93t8qbEB4gGj643bgRds7wFxo4YUq6FL
YVvogwnOtjNPM5e0FdScYOvaZqN+6o02BZiQH1XC3eW4/eTSGv0BS0H+0CTo/sWn
uD+IhFOWX7sDeR8TGGWCUrThPUgOTIXJAn+3knsn6D2GG6ojz+t23zLU5PoTpmdO
GqujTRKe7nIbf1k+OklX3shUNGJZHfK+4Vcg/6tx3OXJkTCd809Gj41dJVUymGp7
VnKHBU7lqWcYtbFcEmA5BuEQ4VLRoJP1Iofl/N6dEUlLMykF2fQj+xO3dZYhRcln
RIl2z3jUXzYvOGp9adE1V18woj+KTRqwu+c3bvO2pmQVwUheswSx/kF/6ka7yDXh
AY3EUBqf0c3Ym7GTVSikpMRp5/nEbhKS7qtn+R1JfjgVYKVIEteD7O9KbU8ao9qK
Od5fQJtMGeblteor+Sswe2hND7Mbi2i58emJHZOBLhHfAFNOTPCh43ou0rVivDSv
oSSpS7IzugSdtk2lkT9E+uN1nQy+mIen1rZl4v30v4WGL5q29Y8R9FTta0a7wwIo
H1PdRvdOFttcZwYfGOVKnu9sXKmf3jbJLk2ldBAY42aA0IF9SYZV6GoHH6VJwjOy
BgNhYYTobTvZ7Thv6pHnyObI7/GWt33zGv+vvNVkDOqixVavAVF4NWk4apiNOtJX
PVpxB9U8DpZBzblTjhNVbAlL6BCLRTUMigTSYFTaCG9QJO7qgeLBrzU8UtP2zPDJ
MwuQsrMujtCIz8jySFHz36gXdUGYcLGunD2G8gft+6qJxWVJHe6/JDz4RWSBNnD2
jZjtQt3Bj/0GsmVD/NlpK5oifmLUcgxs7/iKaci9tMshHnX9aUOsYjHg25xzIDRZ
VfU5t9sHXqcq/ufXBTM/I7FDZdOwnpumulfYFhebPXOAkcSsl2WjmM1nnWBNw4Sd
EIqlJK19TbK6+I2FrWqWQ31PXKqumuCe/zRwjIpL2Hr7VvN7wTJ7STjsSsXHnYoQ
+1HMSfDk0UoVIuRVO9owz85yuv+j8dKid8ycuEsh6HhDRBptXr6hNSayLmNydm2d
DbHhYxIKo9lWuELAsa0MrG3dl9g2jOVVf8wUkShTxqhZRPlobvHgU35CgIfZiD6U
8Qx0GeRDgdPlNbouJRgKdZRRYeUPpF6OdV/nvt+BmdIXYX3vzsNKm8hxdiGRbOko
Zbjqs0lQvdGEl87/yJrWgizTMgiFxSIeqlkR7WqRrn8Cy6a8OajQj4LEBIocKRm1
IWkPVewj9w7ilR19b+wJPXK0OJRAmJsCzNL/s+zqEGYkYqruAMEPfdrZn4egB6s8
EkvkR17I3QkTyq6m0YrocCq8dPE15gvjhvIgg7CojOrnVer1bykFptJGy5Jf1GYJ
RZWv+BClEx2NBQXT6baz6AItQhaAIEb1xJsOSG/09cYtm8Fa0+vKY6rEGLhqy4a9
v5g2dLheGSYydHoY3oQNe/PUXpnbEWzydGDXXs1YVAZSDqZ+WdraySq2i6K/7xrM
LJeOmC+apxUjpqHCxU5h/jub0CKaPrXv7vh2FzGe6n0vE32AzOxdEaPWiS/auiuO
CMqCmWZx0SN0uBl9QhyThSyoBCf8XyFz866miHq1K+dGHNi7iJquuvdbgNO2uKn/
HbtHvmZOeX78Pls6H4k1KXTEuJ5dAvPiT2W0DcCuXg8FqZKVfm/wD8kDfQY+6g/k
+6hvYwc4qJebqzSG5jtj6kH8q4K5SNEEj9SWmjF6XCrmLFeOUZS1uSTxSvpgASFo
aSM3KTHR4Ez+HrB3Fgv77ijcEClMV/moKWG2vFoiuEGGEy9vODHDLfS6ioRRoi7U
IZa3ohKUken2qxKl/oW+33g5pQcMQwFIsMDpkMjB2HDPPULl/hUWwzEu2b5CAkmV
YEPRKRELghoQ7YUSkNR3lpAWkc80mTm/ztEOrhMiSHZoBY50O6jZKVdkYxcNDXaT
/G0IyQx6cBhDuJZxSe8SkwvnEJnghCoFcVdHhbNV9pfgRnHhBrDyPmVpss1N8nJk
PrPIQTXD+CW6YHfdNy+xc24ziMRfwDzXhe/RRhOYpTcckZD68OJOhyo20I+mrinO
5RXLpcGzMAwmUj4MGaMtNuGPEFkaJVCS7xJop3cuLd+RfmtF2warMox5KlcASkOR
BiuJ8PDvTAflpahcVVoQbIZ9sXVuCtxpUShcWGmHnQscATrP445gD9ov768RlQbT
MlST2i38LH+eELlMC2uCybbNvf+2xVleMQ7Z42TgxViGLXZl+DcEiT0HgAtbM4zv
2V4qI2rEyXPF00GtsvgKiGE4lvFyikgfRanjlnvL4BsLBijEADimkinUE1Jn3qTG
2Jmuf2ta5l+/PFEGwVMiUNfuP+gSoTYzmD5V0E8Rjfbu/5RrhcUQFMXOIg3WIart
Z6quG8E4/l2zCXfndfZDrlNxaXYssBhoYQTHI1BCdW0GigAvBPFdCeKUVmVsqjJj
xOj7bPNshLbpjYr93IqWYHDsUWxG7w1CVJ3bLBBX2MvnC94sE54Hz9p98z3c4Eze
45dWEWss9FMr5Cr0pbERVDKHjks53n47hgJoB5tiBh3YjIhiTTdlCERYfmdCAis9
tkgjM1FF2KTYyT7tFUfuqOinxvok4E7BpUula8OfySo14SOBEeyOVHIJdvkrdPxZ
MUyZVnk7cpy4k3XuAZv2KuPANTZsXx2ZERcF17KEDeA7bTRm0WrvcvK3FgFgGnBz
gb9Cj2l1pSlGw4227yZgStCrAxv5PZAQfHYGUI9uwPEnp4ezfZllYAr117Ms+3Tj
HWBH65qxw3AnQsjaGhi0eHwsByODtLx5pXA/+uQ0KuN2QsGhukiPVbFqmiRT3PYu
12t2If32XO68mUk8hSUODBsDEpOxzrgfgA/QWRTIHL51ohz1zmhEUuxKCmJNMXjX
74xw+LiHaC3Q5ILIVcQ+LRIa+0rIaAvxlZGk8HLWVD5yzasMocNcY6RjUv0zdiTM
NMX3Z/gZQXEATHBio2RLgkePYf3Z7YdvfDXmZY9+0zdTKdk9QjL73G5XVJ2g1Aob
Lq44tyPQ0xRTfkTfGX9Xbp7JhZO/sN1lT1AFWIFkUE7X7bupJ/d3tkYC+PDNKANO
yFNmqeIg34jXINAsgsIoQQ3+hvRhblqLtD8Oo0AUidWDW9OQxQEy6szhBsaezEQn
ooNTHuJTaFwGQq2g33YXzIWt4NMdaXaf3wMwxouN/bWjCKNlW6Va97ETzLKHnCv7
QRjua6g6w1YIENGOhFWwbnIeeTtBM5ohR7Ru3S0J5xMIRiQxxV8F6fpZKmw059ak
PRGdoVx1QYi+NJX168L27JTd8/Y8aYhDX/u6BRFoT+MEIaQX63k1C0vR4Kl46F43
NeDt21dcWIsSKuy/FrpJRWW4cFHxkphuKIZ/HObeP6Bw1lWSnDrSipgbPtVoDLfI
ENjM/8zFelBd6CBtl3flvdI7FgMgTRdqcrzEMzPP70LEvhpjG323FUKVfenk/JvW
texAf8GreLFg+Fco0fCvhp/BP2Qa2IryDjebwXiwbBvUVrMMjKd1PRdz02+0hUsJ
pW8wQvfWBqKbfOiBXyV9QUmxez5jBSV1XKa3iYDztd/+IOAyclsB9/5+R7zWjkw6
39yljnwCJgVH36ctFfca9raaf4Ko/qSEiYVAeRKzlETYBMad8h9V+Njk139P3/Yt
NJEo2tDODaBKar8+xdk/jjEkeSw9VQKyp89dqLZJfW9REa2WrqNL9jMWp8sMJ1+5
aQccgB269NnkguZogoCM2UwpCQ2YUCE/t6oB5Dm2zjIXF8tNyVEOfElyCf3MkOtd
VgJgIO/DwrKPsyTc6iGzkDVb53DjFN99YK+2sdHBZmjjMVFYQOKUjR332hlhopbp
5FEM+MIrt8ALU8BjuMBf78xqgIAY2hEkdya3z4ko1E+vF1jx0BYlkLBqSrVkc061
y1cmTEM7esnHXVqOcgifT0y0ip5X862kmCs70hqG8ggzTgj3OwX9r7xgtnKbeYua
aBeBY5dwUnRjp2kwmIi+/cbf4vLL9M8XNuLStWFDp2pUhWD4zaZyfLYH9kxpqhhx
BJSdVVNi4dD3limA/nlQGtb4oAhiUn7d6tWIJAwW/saoNr+B13k3ye6kl2xzTZ5E
F5AGzlZCNy/Dao9IPdEtmqv/jrtW4KZ6hvv00pOr6BQNh3LuG4S+pAUPw8zvhtyL
3j7ANx8WMP3H7dHq3ijX8jpEL2c7vttV4DOK/vsutYgGYG4JNZoMo8blWl1IiYVJ
qDV37DHip0p1WHL/3sEIi07ung2o1on/UznY1NYiRUpMa3ZoKHlonpwgzxgkDxn/
YqqVWHrrk9g7a4666EkdOiAXkH4nruCHyzUj4YnZO8jWCxPYW4RVKVo2Oy/ik8QU
/9aEpO89OkTg8CnXFhzO0d+l5gl4NyBRcPb+CucUa7dqAZTvdhUzqGurzE8t4Sq4
zgOgLKt763k8zJHPk6haDUWLq0mvw9a96IWCZ/WUQWsxqDOM/LcIciX+LNhaINOx
UCd6ucik+aDHe6x4gFsW9mjjNSSL2ADePOxeNOQTbpVC4nA31PWvhd80eh9EdYYE
5X4k+JEx+OeDyYdILx0HvbJ4FN1NHv4sJSyqMLZsQ677EIo+aXryI4p3UaKWJvPG
Iie63WojGHKMsbdslgeDB/NUqDUcfvPez/7R3HlO1WqYzQhdjPcT/R/NSP7m+iRn
xc07oq1uAEk5HYHZgGl4IrWSMOx0DdeuufZHtfyrFa63MdtULcBK8Kliu8qINyqD
SqDBhnPbkxL+JXA5/kKTGocF4fuae/zkvJVGk9nAk7vuzipvdJZk18RKd1sQ9w/+
A9yBvtwbp6Gt7HlzbR/jaVgVHwUwMpEULS1U5G1I3UsZl7b9bzoi3FuiXwS1eD2t
vCJfpkt7cZ6Hxy85rxzVx+KFi1sdx0hEGafwjw/hzClAftLiXFGjUzeLCUFGhpaY
yOSXcSpFgxyIiSuQ1aKSS0as+2WHxrxyb1C2v1oKX2VnVlg5u2dpZrHpIb1AcsL2
AvkwpfW8c0rysW75MEoFR16fEeJWdQ+6/gW57EpMFUBJ3vHAtpa2V7e/kZhlKdmM
7HvUPTJgoXL9hTZAnsGK0kfIa+nhoG4ZkiNP4S2rfK7arH4IUuSMmTXz4D4iEXlV
Jy5+gDL82GX5UlBfxkwOE6UePZimX59Z5gHuNojC77xNyAmKQ9FXGnqrH8vwY6xo
d8jetnzosZRCyi8QoP4SfvIL2MyJKAgJsK8iCG/oEGC197e6syOpA493G0xKAFx6
rKpOzoX/SqNJyo9zhkWFAn8B6SP6Flqjf23AAdXnRT5GjOnnRS6wBSYhbbv9fxEB
LK3UluK3cSpxTDDJOQEd7EmFpATxlT6gdBkaQuqly3z+o2ZdARj2pijGxc4/T6K/
bXjDnwYYNoZlUt9No3+sBGwiEma82tr62wz5nQNGt2AYOGnghhw8V9JXS4hqSjIB
HE8ctLfIpv6Sn3m59Zvz1RwYHcr8lcSJUQrIhxcdRF4ShmlvkV3tpgFBzGB6ugA1
uZxDm4pfxzT45ZO7jMQo+vFwSJs1YHIWyv3r+og1ck4+R93Vg2HFYGjkCSZARk0/
wDJJa2ZWa+/iw7ogFHnRmKxgNE3udqG7Azq8uoPig07ks5DM35tUwrpi0NE15ve0
NST450o9LOXQcUThrKSnTXfWcI4IAv4dya7TK0jVojjnDgCf8OaiXs8kXaPajDHn
01Q3rPevZd4y8ZZOeWPjSalOBP40LMMxT25YnBmC17Gl+ZXmm4eXGnGQT8dtIaSl
UUkw5EkQOzp8n0aiTuOD0vOkYybiPsbBrfgsKcN/EKty3zxnNxql6uUXcljOE/0E
uF5hl8Q4+WxwKWZHqr5mfAYbRkTRqZ4qUGHdbmouHi1dLMcLgLUSZzgN8Rvlvift
A3HsgMg+x8ptTlVjqXHUrn409AF09CnNgUyPZ6JaWzmLrQ4YOZ2+TF/binWzuILT
0JGOmFL5i6MOGBDiGXnIPPMGm+E4BE9iDajBso3ImNetrQs5XkvsSOms/U0IS2kf
1df+tiJKKDUgSNPyLXp0Tbi/FYQcUIMc/29iijFyBemoWdyE5of2q2dwBljve3SJ
0ZAIc+nBl8K01i5Orb1uwapq1dyXGg+b/t1y/SSMa1Pvi6Ds4Mb56iRaobtfOknp
MAddEkHGeQLIAoU5QnZCQF5OCXA4b/51ZovBh/ygAUfc+lewHQVvc6kPJ+0WgYKi
izlfWaWYmpBrfqHO8KLwbNKZuYusZ62a0QGWY3kxFaDQZie8JNpYdqlJ6/9W6bw/
SF0TZ/7ee0BkaqlbwaThJzgcTQrdIxnIhqJngtDKz+OIXTEhbAaapyl2SeCIL0b5
R/WwP/O57ViCMstS5JDf9I5Mw6m8CWwZW7/OYGZNt2/uMXlI1VnCTVxYcUXbMUAI
1ORxut78c9nXMbEb23pLBXLvBtGgIZyqVJDYaXl1aUKTdjb1pCO2FQWGiuvbmWg8
DVUG4T6utP7CJvXow6KpVAuaZwj0zceRWltL+F9fObWSR33PCbolVRHLC8gHFTzp
5wMun/eCvpECdXQzCrIl7EUxjVPBelkYkaMG0MeVKnw2wingglZe7abSJOnMrZnj
ad2FiL9cW/QgjtTj15HuwssinuHkToHUwDqieGcF+LVsyLwWA3HmA2vK/NU4cNVD
/7Ivpx/VatSfbsXpEgo/aXttlWcvSSnLP9d2xH6xROIaccpAEy0PFLywCaTZkw2f
S5Z0kOAfqVtf5Bena14m4pTXsG4MJeypIdvzHFn6NFkZwYlAFM35NRvY9Gz9jcFj
yQRt6aAVsakDO3NCu4ukwArt2GtQoFUvlkfnBUxLou/LaO1hAybnCV3AUGnfnRQy
V6/HTSuRbw4intM4TXthYUtdXaflvrljMCmz7oNO6N2B3HpoAl9D5gVXZ1ruOq6j
xjtn5VDplly1ILd+LBvMbH/CzJ5qQf+SB4luJ++KhHNGSUyCD/0FdbF2Wwa4dT1T
WhDL+N7D1RKQ7GIbSga64Edwe8jPnsP0HG1qc/dOZZ4Y/7Dq47uLt0RAAuJmi5g2
Nzf2JYyOLwcnXdQUkSSFNbjgRv7AGGTIFcrEKzuI0Pwp1xNchoLNDDMTyZaIQ5aY
8RFPOe/bbg9olfa9npYTir5mOoKt+tQDt4pSl65nbKSFsNYxs9hgABMc1kQZAJaD
YDJFzgyuQgUKNs1ueDiBJfBuTDUMSc5YWTbBiN3kf4tR46LmballMj5+i7BYFPKI
AITfs7+6VTcdwm5PgZWuGzwNithCZQlMpuSiYXrxxhPhwUASj0n1erjCnkJyQrFO
5eSNs/Klm5UI8BvyI2kxhr4vVyga24YGWMCLq/YbT5pnCkcEfZVaL40oqSO+tn/6
2wxjTjARhFexff+MNVxJ9E3vSBjM6RC5OfB+Ykqn9LFums6/sFxGRCO/yxhMsVEM
NueuAheqPHXKl/6db3hIEQJkmkgO2Mi/3RBdE3qpgp/yKeGfOdS/H8s4Nx2a/579
H0BpdWpdh4LYA78iWcdSY8Qc1XgAADayizE2gXPQEhuqJYluQJsB+QQ6AAXDmGRC
LzkIcYGDK4kjBa6KUU5104pm/K4A02aUjpGO92riFbY72l+w0vX2K8fby1Bnc11w
SoBp245iQI4K07LuiblB165SEA7dCan4zBXglaW5RHEft9gxoYwxhh4ovMD10TF4
UF8AS9zCb/i665A5ZVMPUT7hXoFcP3aj+dk82BTFIwlPyv9dpiI7sVIkHY1X5QYC
q3OQMOdfoSFw032HfVPKIJDC+j7NHMoOsW85VUlf0ACTjyz1p2OR1qAb8m3po8Xx
YoCmcTiZ6DFjbaMt09D2fCq82dmeT3Dg0MiFkOISJQ5eqWAAlo/h8T4O0gKazOUW
L+/7HIee0cJdktjQnaPOvN9xTcFnsQOBdB+ImvUCyGl/LAsWGxkMXoNrrRGHcdw2
1VEiXK/X+V7thV9HHbpfjm2Vuk6fvQ72+Yc+P0FEPFgIvASnJwgd+flkNXX/diYq
YH4/p18+arYV/f9SdOD7IlgiDPArKL8UKfctNRSWV+cr0hWeM0qBajm6llq8nW1p
XuA1TApvv51kPwEE26+JuPp2PfWVmv9PXZYCkRyXzps4G3CwddOBZTYCtpWll9VG
0sLIjXIsMf1JqJ+1VbaMelasGGxJWtoNtznSW4HOidezGPKMwFVQN7ndlorjgP8p
2XmO5aaeOhUjwO7TXGFgtpassimd5/dcE75eBizB3k2EvpQI9p30slURrTlkCfHa
Yqmeoolxwnm1JeH7RauQ3fvCrcrP1GuJKPqmqCSMX7+CQ0fDdZ7ykuAE+v6Ypz4V
jGu8Qf0Rzra3+tSbiDSwhLmGJRVdXZXLQFDSaE08eKCDzy1LdmHmd90ERwuaKM1l
FvghuMwsUcHnqvAgLeOUR7Q2IjY3yldd0TQ4vFa5CVZ/cN1A6IqzAvW7ylNTBecZ
P5qpj9DOzIy4LTtUgCa1znV2uBNo5+POlT7Eq2M6uPCf4+5pCvmaopgKAmpCpZM+
BqzdPczA/nThbtBzpoYDp83lFd4iedRS/5ibcXMAdTVLXjUWDX4WxzNZB20ghlSW
AQwQ5k/HNjBoEoiiBux+6vFOY710ITMSuV+EPsBF+T1rnXYHodiTCv0+UBJCIMTK
hbGIu20kUvd9w3kMoc7OHuf9dNzSO4noRnoDN+qsMbavQbCUmr8W4YMMioRaNpUq
u3oT1FSePE3GSz2/6D+Su67HYLhlqMHnd1egj0PyYfWHy2dbTg66r/KlSTjd4Jny
EZ6S1Wg5NizbNCzmi+vkz9iUXV62XCjhxb2x1ekx9NX0P3Ie/QhUD+fW46HgljlP
c2R+ZA8UrPJj3HH3MYfbfcT63zRuyuK59G7Rxey2459cmISa9NkaOriSdvH1kELF
x6zCchUMkoGVu5qc7G/YqU0VY2NKmM8WQBgZatWZHwRUZw6RR6rJ1n2/KwjZV5Vh
e3ItxWtux0FpvOiR71g/N1MjaoJvpcgzpwBEfYOlBvfezZVgFuBnpM53yG64a0ic
+qCBcRmZ7dj4vjQ2gJpsM8cDnWLDTw7Nb9Y3SzJMmg3sN3i5EzzgJz20Ncf0KmAC
wYvqad7K+WP6lLJ6RI4xzW3C926SvtMyMMSxihrxOJRgF0nmMMkFCTII875KxvWJ
LQdWWrXbaJXhEnN2RFoMQVkcbiGextQTF4cnUo5+nml36+019mijVBSAQkcEbSls
W9zBE16UnOVkf/e7Se/BkCQckfCvaLMc6H7P4y2I/IAD91hmp1qtsaWZjmeGrj16
qrFMOaAOKDODe1xNJADy3b6WK2vnWCik5/f3sFq3ixGsLReDtJygnJ/6YOkQZ9Eg
IgJ4clcGf+H4RTGRe0ab150PKILxo9/zBqCY6Txy2IMohiHOEmglUT+t3k+YfQLy
PXjtk1X0uodNdSpUtM0u3opEzt8YKz3jhto7bQXPWN7GWLSApbbjlCMo3LyCsfQ9
pMiY7HNOOAR84FbODu9vKWRQFgopdrG/xR016GQdo4zOUhx09i4ib+VG5Xi21/d1
gTRgJeYIuiAAhrdDoqtDUvNK5kTdV/o1G1wwSm+3koQPhGowlbMO8nydPL9zYzN6
eU8oCv/Ti/TNr5sK+5yYDPBYrTmPdmN6A5BpB3SI+XA258+n2KTBPJNDrU4VMrHk
QP5+6wHraOQslr8BS5yHB1OhEgefy1bpiBuMw81NzQKUVdpzvYlLcE65uRnmMioR
p4KsyRXII3FUdFV6wR18HmuXgiaEhuks0eQ/+qzfFc/M8/KrpE835CdyHIvVjGaR
k4CkwaAAcRwNy7sDuTmy5arWCKGFcZU79CqxWwk+9XCJOF/jzV0yiluVlsc/gXxG
MuXUd7ohcFp+lSoLswQvqUVeLw4ZfXL1hYgatTj69Mk+S9ri3AZgFezyuRJnvtrY
/EyPgXdqJUySl3lNEBVdF2b1L8sSPX2I3eZ15X/BW83ZykePBAdLLwu+QmSs15ST
nOnrETqUSc8FXj+b8fajZJnTJe2Ie2yU99X5C++UvRijpn7D4AuPhHxYb5WM5Jk9
BDX546kYVdXbrba9eHxLKLL5IkdnhsfWl+qmHQEd3yF9S71g1+QeIm3vWvuAY0XN
6xPNFVAdwIQZWmCfPnG824cjCYA8iqGmW5Yc9owujafmaOXG7Ta+MQge5grHBc3h
GcCkfM9tAlHLkwShPJBt5e7aTFQTMG2DLGYjVwvGn1RrpBJr/BaVMEz/UcfUnk4M
bUS1maJ5OKSUvey1eR/OGR/+bndp8PG+OUAM9wCaZYXg2LlTKqPMaTu7dq1LQyYA
JcsY4zwrC/CNGJhlDwfQg+dFRNpNB2p5MyE3iyExiJGJI/LiwkCHNDdJwkgk77sV
gDTQRfGjf4fiFC/LE11PtKodcqpYCZmDsl0U7OKQQyrg2NbWc+y4t0aoQs8bCjvV
LkctVcQcyD0f8yMgdXqF/mkBar1N90no//xvYxeSAReHGjvxQmMjXCeNMKRWf863
gvL2aMjPH9GbGFEi8lI2/hE3gdSP4uMFLMa9WmkQ4xitwJer5w837b9LDWD2KNTA
3Pyo/oXU35FmgPbieMICNcxR/nUz5j49izk2tn8mIMWvSe1bu37I2WuB+nylqGAE
qvmBHKBpJlWX2W7QKxm0mCZhuDWIJ+HzR4N1fzFYX9dBLRJUkLZtg2xi3NmOoqvV
ljSKeeT/09aGBojeWzuq9Z7q2aIHMs80PkFBX7RlTsd3GfmchDgD4hkZPmeBkkGV
DX2fC56DbkSFVr8bRH/rlslqnHVpPJ3ew55gGc9FrkmyZdFkX2V9SSZjn14DHWbm
ZAFds6qSFK+Ba8rV5GyrouOuB0NDcGWnLNXktNt7BNhxLaLrsTRBpen5FFIXaRxl
5lBR7q3EfLn+2JiNk6hKTjXMNXltm80yGFae9/A9NHdO4derquWM43V5KXaMATN5
7kNGbIBmBLgJBl6ih36ik5/NypdVal5ZF7thm32TSauDZLNdT/U+h5+LV1LlPP10
m5zd35rznXCK+ObaNoPtfr3TQMkalcOjCA5ce9+GrVAlyNxAGeWccsZgU8WH3fXT
VpG97kUP8FmBUrhWsHb1kshlYf56QjJJEcLAYmIFtojWPEkGJH/N4y59yVl+BWVq
07VmbyN2YPo8fAq60BM48GfJCEOCn+11Ja4TbcbuX+0YThbs5WERE507dF4E5ToA
ptkerh7/baAcgdJ59zncjttOx10FA7kvBDOnsDraLgrtGFkHeKbYai9Dl4NnQGP5
Yp1qucSxGnh7sMcilgWT6WLYYGQ3eflLoUqUAzsN//ujh4dBZSlzR8sqdXDFtyjx
kwyMAzq3aiaFbb0VRn0JBdipKLLd7+7RETAGCWEV8E42oGhP1pRaEUNLL8lrMtBI
IgrVgrF9+avWm5Dy7fbL7EsR5kkJvvraGRON7AcVQeHJNxZqv/fN/UUlBx6yfbE8
Osv/kU941x9M65RuFNdiotv5/JA5rabFchAs9tWLLEKmcq4KkXFw/WeTWjtu00Nd
AoXelb5nJ++rYoP3L+XX9l/x4EIIFQa3LP0a2Peurq0xCqV/UCdQWe4yf8LeGKcz
egtEoYuhsUd7A6nKWhImCRvdBPk05E4J5zjVtSUdwTn1n2cgH70SzEAMnTpejY/r
ujNTdLMDUzJr2PVFgzU8JH12X/bCmEkTPGR44VPC9EhjPFSV6w7/ev+1jIAnXK/m
i0KAlcf4PHWKNwPjHnayTOK6/NbeRRMrhbdTCJ3oZQlhX6dP5SXD/HM8bZTjfqqh
qs5KkYOs+C9xNJ0w1kJl0/PrYRtVxacJszFJ3qGgHqCc1IV2rkIAYHbQw4iQ6H95
yEsy0r3jU2zaMfi/cw8uf1cWfn30udlBwjQR/5/yh6BMWWDWCCNDzQ+dP5G0soPu
97Htwy8QjSZFqfUFRoNiUVE7l4c3mWkkUP2PFRQt+70E50ybUNDJKyrBgOIt06tV
dQ7TeWTUsrSS/m9fFCaeiCNJQR6wKeKjDDyFhDup+2AajoXUatr1ptfZaadr2Wok
632iWmDsTYo2buXcc0rT84u6yN/OIplL7yWdMxrqzcth0p0dpVHq55zo3UAD4uk5
9Eer1BF/8lSGGl075RHLurn9a+mAdU2p2VWodv5IRWitQ8wUEv3cifodsh4VyEI+
2z9T1tYXudecbmWGhDe7zoMRJEwTKMpGExR6veM3wHEVr+O1ANGdXi1XF31vWUYH
U8NpLCx44yZ43NB46I4fyT6HA8KPV8JbFLcJWviZhK0ObhBILhQvjTG9+wqSEFos
cWsm4AXyb4VoZtXwF6W0HRZ6v/uwxQb38iWzWPpu5RDkSroDrB7Y+NVAeaiLfd+d
mH6Xj7JbaLX9eD8r95jrsYo2mVWZwEMA3yckYY+y+P7Of5uTSpSiyzufxv6DonZG
09eYeYCS6vVLS5CopkZ1Uze3Of+j+7pMxWk5YZkDDOpEreZ/HCSwH2tQf9iowC2l
UnmeydX0Qn1gdqsaCWb+UNH4q0VyYgfje5TfPK2HVBcf+Dufcw/iX5y3HbpuBuTl
3VgB1seoYtKbfWB4CzNvHAs6ZfbPLMh9GkPRrSQl6/1wJHdAZyQZ5Bv7Y/HP4vpP
naRVMr1ae4R3v6JYeubkYRkbkTXhAhgi5L3wTWXEFXHqU+TRrZmlAbEyglFrq/sp
ppaMdw9B8GCnc78Fl/7FyLdXv5CSUiooYxbLOPMxqd7aQ/XL+PviKwIHnCbA0VYx
vfCdaIewSfTMe9Dt4Wx2H/dUGJjv4tByOBzzVPvkq0SxHh8gQ5l6X8IuSFVbxUWf
RKip+Y1KYa6W5nNZgYz2rXYTjyissF1e8xJIUlZNPWHi0vsQOwaO1J6zcMP4+Sg+
ACGISnZI1o+D8fbSFQRLkPVpSvOzhnFsc13FdTDaW78fd7NfgL8oWMx+cOYDyioy
3Y5HekquTh1U9EQXDqwyhOsHd+6NHKebx342wxMLWnWgKpfvdIhtumgiEsA8jmRG
LN7YNUESj78KV7S/QhrmY+J8GWQRRf+bSJ+5DAykwi1dul6aIGgjT0/sX1uCZL1r
vJsV3RS8fmqGfV5qmIkCQv8SGY3b7Bq59x4704nhW2TrOD0joYu+fFM7L+UYkcLF
o8/awobwd9PXxbv27M9Ja/5Nq7OJWguye6l7d2KSSOXSs7SE0wP/d1iE0OwfhDgg
Fs1C7/r+6KvJsdnLjim4CITc85a3Yexb8QnCWzbqo7nRWajRLxjjGcNx6+QK82Jf
O9OxBwyXdQNVvGZ0OdOn82Pjckq/isQjYIoqrddZiCW0sMGiuhtHvbU3dfE2+/Zf
jzwILj62SRAqTMaAdJNfb47kum+gEC9oMTp4S781hC00SPgunuLMFRd9Hyn/plWV
jhFSDyDdN0nx9yVGGZWwDDYaSqfylAnYpTYdbu/2cWXsuGzv9oWd42Ey9AoXYpp4
h7bTgHIgkgWF2SCmt7l9jZvJ0boBLJIbIa7oEELDUhDLVbBHidFBeZONBLdDAgfV
khbA7jfiMEckwFDovtTTCzEUDawhqsANPoGarfTJfHR5jAQ2fzem91rJpzlQqtVt
jzDcbA44bd6+0G/X0v4NAjmT6vJOaC+ConPNwJUADzupFx1RtASbYNqYf+UTdUqZ
YbWwqQjzEJWUF551Bmy23sq+I1j1vvyJRgD1h4i+eiSpUxWfnox4/q9XYCT79lfZ
ucePz00lG5ikETP2QK+n7X+sCMUaHkP68Tg1soCW3Y0WT5cYHecWRXcJbDW+ITjF
zn3SKYYPwpU0kr0TIctcFf1pwjO+Ia0z1owDJJm1kEOtoF3QtuuH7MX17BJ+GvBP
TxvUMuib2OShF++8jbSz/BZ2ogbpp1/V9mh98eXVpiYH++Y6O/z2raD4M9EDjzZi
UWWYitk0yuwhgTrDehoFZrShm8Vuv+ZAQ+P7Q04LXd837RXfvhZspILBiJEzy8nG
C0d9diWgFFWIev269tjhuNyTyQ0PDngKntTMPuiQ6K1Ovn41sviS+daLKN++WEN7
9am1cw4pav6+SQhTBi3qEuYbX3DHIoMpuvPu0ESHOJdvPzH87xm9aNsQ0T+zv28a
yMXtNLewneN7fqYLmF/JTHzn/IsFWxdrS7ZJfzOBb4lYi3zAI3AvxdZaz+A+J5Sh
WuZL6lWsejmBs6986bsLw3BIEEvKP5kQkDkTCxUF9kJJkrjADUx9BdzMmbt4sm1m
7lUg7o3n/jp5sjVy7EsOC+Egg02uU1NMKJNqA/JuARSkFm1pLIEEVzn8vStVSMOe
rCZkBUCIQSmP3nIoBIVjiFO0BPCGMnKOyEcalzog4FLVlyRsqhdhG0lG0ogMaMNs
5kstOYPkPv1iw3Y1O+UwZ8dy7OUsEfaWSn5pckhyhgvilPyVM0tBfN4oeY/nLjUo
QMxJDJgd8vvy/bgXhhQJx1BNBwgUj1FCOkD9XyfG6OshUHl42qiec28dr6SUwzjm
ptw0/axkshtLWvzT86Z8HAz5TU4AlRr6AhRWN78GPkfX9spwhFzr8kJjZVIgC7d2
Oc7OJ9FtUbsWkAaDVSnlD9HeOQwc9rXzO7U0MTKfNe6ufv6y+jjQi+1KZIlKNkYf
1sz9PfBLseJtnOSh3QC9I3OuIzBntauMboDG2tNg/Arb9kgMS5VsXl49qMlKAa3D
0+0qllJWYnyW7L2Aqlsw4aWihMqhvGAA5fM5irsQFkuZmKsNRSzAbABqSLOMv+mn
2lE45YB428qG0a+lNwuPpB+1vED/e058YsX7G9B9pmetJgNcDxx/DeOkhY8jWAYJ
Q1YhHJ67JRIgyDJePowAYEcL5mfTLKYSRUDePIg+FcCyuGPnchP1xC6AZqIGYnS1
NWr7ZBiY6jOHKbSU5KMBVaY1jbZXrjuD5lG/FePBMXHQIfy+26y3QlCx3EZYh9nb
nVHrEPfKzwtI8VyRt22YRJ9HNP+cecxo8oSfRmfaVHKOcsu0DUE/gW4seAq6WmgW
T+q6lbnqOxSpiB35HrMg6wepAnAhUkTWUasA+5D8u+YpqOHo9HsfuJbaBkobRrXG
taRQYOBFxsU9teVUZiTmekXxBw1FKDQXoJTuKhL4IOeQkL1P4HK/aBoksDF/u7RD
9kUGMVRAcOV+/aOe5qiGojADG35LTflELXoR98q7K9QcIL3kyAxNQ5r9PkkHBvIt
tyzyXVQy2Wt33vK7ETvI+a2S5BhdWPiz4LNrG7nICbA2R5hThfhGJlDDvBLGQvmP
lykBSipQXr9oPqH9rUg5c2SYZHzdsy7ewRpfEKGf5c9LFyyoaOKrs/sK/s+nXlcC
xSZD0U2vdwcHP5cqlCVNADjno6dCgo+LJqIcTa/A155GZzPl2J0gQkuAfGqRXLc0
mp4w9kCzWMZN/mAOxA+jUer4KaGPAHs0aRYXMZW9VPpEZ2Jd2kkxHCZZwFRkVD14
x/IKW6ko73aGdMcR8tf/aJ6Bhn5rAiBFkHXJr4beyx4fyuEXhb+xuzKvB+R3mKlH
qaKotw48JYBUa3RDe8gkPFesLYOgW8irSqzf7dhFIP0VhryFGrPJIOtg1E/0+1Hg
+0IbiWIxh5zyqfjyQ5bVdFdUBZjQnrhyup6hZKcqLipYSTVhfgsA535leDjYeCal
yvQqDiOHEgs9yZ9hyPLVVGRYBuTN1uyw1VTs2fdguArZBwTyxVThJtIPvnKUii1f
yqC5VaZoW9gHOCwW6VOqP2YOF9qY9GGkygX8T+JnrsPXuhO5dTtnlPJ7/ElrHZqO
iWiy6ctKg0+sd4sB/XFJMPvLmsjnBzDbzS5VBqdZPQZoPi+sfQUwQ8xqSin5ap4v
EwxHP6DYsZ40CKRV7X1p5heOkABl42QLwgh5qfNx6VAICXh1yPIvYwPtqOK7m7RO
qwmMkQoNnlJQ6m7VI9sh0EKXez8c1n6MpbuOL1BRPi9Vw3sfDjhUx1IliFsCz3yX
+/RGCGCrk7xn/gBVc6Mj7pXPFzWXWWPFSDHval6BtQKZ23cg5mA1+5p/OAjavCCR
bUB2E5GszBvTT+aY81BLZwQMc/wUmp9KhHlHWpwhHCLSpYMWxEhZqnIpgfTfmcVK
/h2mpE5K7e+uFMPm0DGLQz/jDJZGmpGe9sPivdNNy7KAIzgpW441/3nnq6+08Hb8
dKZ+VqlCxv9359RsDkM1K8rmnSyaF6FHhIV8PN2lXrZpQ4rA/Y/L3HW1/dr9wC+o
1eVpJFBQ9h/aQvJQNOd9jITc2a15BLE4MO8cVIKJCzZ0aFbtIeWJaE/JqAsmWfdW
78avWzB5dtiN2J/7gLipdAm1mNE212HnOMxWMvCDutBTCNkloVZPSNONC8Ry4h3J
RiM5/r9Uu/s6vYqx/SvZgk0Ma8Sc8rbVnwQVfMoAZMrx0lxoGTSbFClipfHDDmmm
xR4vkIzYdCaXIqQOnb46lNBlt3JGR52/+vkgHxynN2Avo5tQLaHhvIhWJ/V6okog
epFLP15sZU5PWoWG+eP7d5FoPL/hy64WPuLuTTok5pdyc1V5W3AiDWsF2kUWrZTN
LpqfzwfMU+4DPSW7xWRDCB+VTTWg1EkjCSslsR8tVl9aFZEBnETOV1PtUZSD2KRf
xFAeH6ZLTLn9yRsqeW0VgTvr4yVX/ZUGyLURekQThwSuJlK5LX4mWTCG9hddo0de
mJslmPARZIemIDY0I51OKL4vT6GxO0ZZKq+Ltp/68A3HWOer8HI+XxqVAhJUHgQ9
tUICWpucVBiPKDIynS05kMvoBf5mDL5lqbBK6ABvAtQ+L9BG675dHjqlSMlLHf4G
4F7WM3r152hEzoavGnhDkrgiOtvngLQyVkyxUvfMozCqcZ6MWQ1Tg4B6dtMxZFe5
VScEVmwfgZy/iGQAmDEiaNDw9DQGPJIv+gYtg5aQyhJOJsoKi6usROueBiPgwtdF
0KBTSuckgpYOvehuI1z3GAvsZQXuAJV8h3HeXEm3/5NZ80JDZEsS9M55DzfqpXqY
WVrMwDK7PbgkSwiGOuaoiCfRFR1TKZeqE+zBP+5lnzZaFlUaplu0ykJdx2MLSbFA
HXswLZ4wOtAOPsPeMNFKCRXnh/RKwcimBgWtqR2E9RMFwbBS/jgXFefWXgzCJZ+h
ss7gdNzfsKOSHVlX6h5G8/Wr7S65Hh4IVq3g239u7gfkoenjQCA1T6zm91JTpZW8
MWeKX1YNbWBQ0Izb1u+NvYkvYGmz477TDI94Di6I8/FDxXkGE/apeoPV13G2k3IP
01iZG9WVs5EOZHLq8kXicsCJOfkdaKIwCo6kETzT3puPbNTgBYpXYMcdy4lE4XB7
lw87xQ36HliZsacHd/z6uAD59J8aqjEQ3rhPzeloNWV7W30zSnXrVZGATCL3H0Uf
wd2jwok3ehHAw3lISdylI0V7kGLf73R3oegfmmS4eFO4Q3yIaShgJrmmaqUyK7Ls
eToFDvtu6zfJqIH7i6e6/d5VVSLUYDM9hzUmkN6739SykXe00q5sh1tF1IuqQE3R
05U+1RZnUSn1i0Y20D77E9MvP/LiCFExzPZg1uKhCKSPl2CmS0oYUEPxBWVkl9C5
uHgfP/T+YBiH6TX26nSGnYtoumM6kStCN5csngmX5/S0YFzPV3PSMfE42pirBQ+y
uCtkPtXPyKDEwFI8cc/G05O5IvriAMTij3YUpL0H0YOQDb5tU3knI4BlqIwH0Vr7
oMqG+KyAdC7knEs7xrgJNixnidAwLeNwJukEkyiMS8zy3kUj25AJRp7JIGNZ1LXG
icMI1C31ABDr6RslifMtMyzpG4SMe6f0+bY4Phh7TbN5etFL6j+v8AOGuJ+H2GB4
Gv/IN2gG7Ke4r80oHasn+AS5QiOawM2NlxRT1/e0KsKtjPOWWhHtjZ0jY4bTxzDY
x/O/T+tFznCSIZhQPQQp4xp5VJ+pHicJpglzW1w8WWjWX6G7d+X9aMgBjPJCihQj
Rn8RC3v4+QUq+NBiLE0zKbuSutU8jFGn2AxACJ/jPDGMhVaTchqhQG862Njj5Gjv
Q5kCBbdlLhD8XhsJPZ26lhZ0pvrPAxdYeFu4Bk+RnaHcw/x1UCc1u1QcQJLCXgJ7
VFVntjnYsdX8aMygbLaHpRALjyBhbfUi6+bqLgZ4h/T5f0HVptRfoAiWtMnHp/Iz
GLiy2fehgTp/y7OxemRha7a+hg0jbZhSuw8/Di3DO5gaXHiAG70zC77c6zAXC38a
RTGuMJvy6M2gEMdzYONY5ZbWHIEdrjtHKOsC2CUaF8W4bWknsCfsV3jB0ZY3tLj2
JtgTq44rDJm6MEzLSDC8lJtAvTETj00kutnKJtP/OA+nW5+Cqdra46A7w9blNlVT
BVS+iRHXfjKTS62BRKIWzLdLVey5f/vmgWgSXKELyjFFOw5eYqHfUlUvjmG/a/k0
2Uj1xxH/T3WXgYB9T+LAJEaxkp+4wfAhfZ3qXgNHrG8ISUSDAGWBCMJiPOqTT1/W
Zlyxs3SDvo3gM9AzS57uN3fk3hg/NzU7FAkaCHYMFn95y2KS/o07kUHKKGl+9Qrv
qUfXskyRhzDUGdgVqbaT8ObrIbpqTCxDGnWW15tPmqMWh+K2k7Seepm/juQCzZHg
zL2ZbMKsZIaS4RuyFsN/0wzz1OWYEVX9Kmt8RzW8Pu2l7ve0+vKkxiYK7kprQzXQ
fTnS+fPKYGmPrEgC4cuUUz4vJA6LyH9pnjD2Jt+coX+dUKTVLgI5bJ/DVQEFS6Zv
vCvgkVtncK0i7O/i2fe2od7tDQIqb9D2rOrPhejyxQ2jvmILESC1i9qEN/u0h+pv
myKdVs9vPk8b+jDzckgwcfdhiSFMFZpzxvQmZURagwZbCuwEfMGHNM8HGbrIAjRE
r23MLkkSHDMK/cbEUVrncGgXLd/cqADqdT5VA9dsy10SDMzJkcwn9W1/2VUa8J0U
GCJTlDMUK2qmz+xWJWiRrRBGnvq++hKnZrgKjMBjXTy6kZihBui+I4vuIf1viXtp
yGH6QfzsORfx3VdKfvTQG5SY196d/PGLBal5RCjZn1bfrUPeTn/Qe26rVxqYAMlB
Vgn2OR/mZdaNA8xVNdpfxMUmIGV0a9xHKvLwhFxowOHvgMQGrVOaNwXbHiqZUkfC
QU9Dy/mTR3Vs8eGmWlwYrVFE6mh307JTILBkMh0RK8P3PNcq7uB5YXgKGtWFD9N0
y5NdHn/GAnHFPWcKwyBImf9IRXz4nvjl7ThMafugWsBF9e5JX++RFKzJp4l+Bur5
97UMj00eJzqK0gGEPIza/gPIs2uFDFDh7Py8zMWFFx/ur9D4fiH+uBF3TyyppJfK
71WHiE5zyunlYDCWRPZ7QE5dFTa4j+jKmJxDQhcYhnZEzOFHwyvXxrAQetU2nA8m
pm0YJpjaXRVTW2nf5CIonOnDMtNhA4pblIzF5uUGgEPjRK2xZLhBSViutrIAXwS9
8b1K8pGpCoo8oHfNSG9w/pFtLXj75h05BSDUS+qX24xGDkMGfVVv/DkT5bdOFwUt
TOEMN37GsA8GCFeOhePT7FXQad2PWCRe1KjYD4qo0pkB9l6VmcEa2PT18UbSoeZc
dHk0KUs2jgJrgKZxCd2MAE1/Dxwjbj6KD2i5WF0G5C8wyrmFz8+umic+RVasiQRY
ZGbFMlcUMgGICkJ1Ms57EvL+mh49ioa0O5ywzNcdBkhkTAUdWVFU4KzHTo3xUX9K
biHzWi+6Sm1FHxtCs8BANXp366XkBms8vBvUKSB6W7Hw9/Z0NVJvu1XsUFTke6jR
jjMH+gC9OfVzREQtnOapt876B90RN0we8WilUuP4/TqGxE3LSfo3EvzY3txDu5Cg
tZ0GfVhic50Xgb/Ry3AWVFqX7Eyqr/YwnsNmt1LAtdqTJudnMP3ouF+Q4BBnFe+H
gZP5SGn2YvYDDrAy25zAomw/rUNDAFFXKM/L/TDVllh1zc5yLzHpQPXVxt7r/15A
2l5bkMf8k7F5FYfEeX3bBsozEZwNiSeyjdhvGsmJ1re2sWGdOYZmlWQj/a7jhxAP
+r8SvwOVx7uYrr3WaL9Rijj20Ogj+0NLm9LGHU/nlD/himpPkHUOBCWY9LiAhjHN
eM+oLIuJtHAYJflpv69KYBWqNnnPK1dsPx/rgFP3MXTjE4+Vdw6AViTBigfcKycO
TqAW6DQgwGEzO7HEGMdI69U44oECCufHpZPkbByFm0OWeaVbv7fzdEDhrCTBelgO
2UkOIqVG5pX5oMWdGhuW7Yb480Cgz20kszjxWb+Eq+sGTyE/dGCKs1ICVaQRw8ta
D+VFHE/TGYvQ/+4BSflk7STRewvy01fzepd2ydn9x9H6S7lhqswRUM8TG/Hz5Ti3
gi8wlh2QVYPZbWsFZ/8DzBd32SHIKNaf/2M1cgldmZ8JNokviEVlTd+2u51g2MgV
t4zNxtN4hHKYtWuiB+LfIG2TiC7vi7NQB4TuOmgSl10l/XNV7aWYmagAUIDwYzNv
f+HDy63/h9XDE0FVfWSR4o+ZUEohGOT2Cy3dSfzhpDzCBJtlRWomhEsdtQNzRayn
WRU8bPTbeAW463hqLtW2VGrCtWSbs55gvp6XxjzN/YAAn7xQnEUZQTYtLdDXbqbm
V+qshnOlEn6MeOFoHvId82O93QfM1yhOmz8VLjCsLKAZl0TZOz0Y2uCCBPH2jg3B
tEqKwy3dydpHI7bGHhGJHXUfX0PlOsQLFcdCEzbZSVZQrl0sXFuVu+AyNeBohNUJ
c/T/xYheFj5usmBzKdV3U4OMbRk0zXm1LK/DxKeBdcqXyBvWBr50eMpYt5qiC1Fc
vTI/zIDO6691kT0A3gABHPOtFloSAdotRn8tfKhRQ0yJtHWKSNZUbT/TD0YY7A9i
udcJvTp1IuH/F1/UDYouarOyJEUdl9eYNrpbGFGIJcTsqZ2lIytyHWhKcVEY9LbK
yu+F4In1n7K0Q9K/FZFzPSHEzYltrj2g5QnPulFGwbN4lHiTdxgajEgAA61aNSuQ
cjElEHfLiwXSd3NEuA/ZXjvloEandHIkcQQ+PN2yY3l3TqcocZsprBEY7AzCbek9
1ovFGQue6RTp/owqY4e/PSUGh/gP1IgZLMDOBWTG6bYvLAQ/n0Z1mvkUHpRUtJnI
4yTA0Nzxd5s8dc+HGVySwiZC+ax81kfgXBCJ1c4O39ufwqsTFLIHl9Cz2WFSyJ/Z
73k6V19SkYzcgcElGlOnhOhaKxQQ5BrDg/WV5AMlPpVqnd8r1vpa6IP+XZJqa63e
nhFYFrHG6enqKOcO2BEx9psCPFLHB4+P5hkDdfztbcLC/91vZO8on8FFt7RQNdRK
obCx8xm2TjIXn+F4v0SaFDBmEk37HkGgYogWAdWoAm10Q+/moj1bb5KlgK9THc15
o5Z1FGFm1Ms79YnDymIhQx90r/uE32nfLs/Q7vS+0TVHirkmvbJLcPIGW45tMeHy
7RzuXeYgZbVPXV1TkgC99O3vyGMSowmf3egh0/jZGsGip1DRLFWFAcMyMmJAUUzo
s9KUPeetYL7P7kg1lpWpi8t1bzUzLBrvQezmUihWsfolXz4AGgtoQZ9I2for9NTX
1p0ORqNK0VjcBSlUEc9mPGbIxOioJF3+QI6b9vT9JJZWwlbTIp/vnXsn6Dt4Vbsp
o1tf48FsZg9Kfhv+N3d7ELr7UX2hx02ia5H0JwYmXe4I7f8eo5aGyooLgWz2viwZ
iEmO/CkCtqReUCaHw7F3wohXwR6abUrgEPQGnC4beqlSWWysHNDr9YVtCeqNUCq3
FtOSk803befVa/KEDBhUm6uZaNQhOtJjgClqt59qA2u54l/bFhiWIPVTqIDvczXJ
/PRe0Rtnf/sq4QbJplQmu7MjYrXgAZJ3gWQzS+BnP5HzSGEnx+j8QvhDjOoMNKrU
0zvPS2V3HLzhERV4nf3z4JqwMZoJS8WYOyErQNw4biwJa1F3a5r11SxnCSwHO3VV
SlI8AomGfwRJ/13MgYjJwYY4xxrvcOlYuAYir4jHBzWCHFxjDFuiAtrYo8or1s6u
P9fAaeh52fHAlJdDEwqYti3VPxTnpVDwr7wZsT85dpix19GgbP1yQ6ovf6alLolK
gdyPN9QscWcdNRKZb3ZIzXz9Uklj8xffNGPCBKIGPHPLkXcCziS5i8rk4Gf0N2WO
MDCkyMzZHVUHFT/0Sb/8ZK/PYOquRpows0vZsE+EsvzgTj7V9R5/rTb3Q4z0UXmA
yijcaTdfktPdrzi79RnSkwbUrb9fjGw1pn2dCB7U+5yo7qj3JT+kKhKRrn8TFbON
kHEVGKFrAMz/1rvVa0w9P/pgMJ9783cMVdnA8q5l/40/7rL98kyr3q8z00P76uSs
Cc3bAErLOmcc/KcmGSPtc7HOYSfaPnjqTG8Eo0Mule5G8UUUIhclfMbBFL9mApFn
gt53yja0I+wjTNxTim5uy89FGXTfXZzNlZ9w3+foKTxtAoPviAt1SW5te5y/P2Ez
LMpyNTToQHw3zfkdUWfHiTN4hmrk/1P7SeB0tWK7U+UU8F4ty6uDMB016fupIwJC
B13Phwx+dkgobCGcu4iEQOU2zm3PusJQkRMUGbJn29ra3mnGfvbdx50UsZX5Fre4
9AqNJevq1H1mAjnHEhAAaLc+xS66e+W0xa6qI4ca0as0yUvmyuZZHtmy0rNFnFQC
4k+6ou12FaV3LjM/C1rq+uTYKpb8gNTU7TfZDi6FgxjYGxJCGN91jclbq3CeZrdl
aUk+KT+PtTSgfVNaU+ffGi7X+VdLt8iLeSWxToivtEVNy8hh1wN/BaQZPXao1D3R
CjxPnoaWrfpRuPzZAGcQBxKNBEWIq5CkXAuytBAdQnXoSbmMIKBM62WvlELmq1on
k6MK6dgzwRaWMrPnDBrFR/FP7Yyx7J33cVD8JUj9hadamFg2Rjhj1Lrf5UdUUgV1
jLuI9Is3exDngFkJY58WTNpAkvR4JP9u2/iA4RDA+1EL2705tnikR6wp4MzsUUov
iscilOwRc8rVFK7/RLtrocFbk8rHv+yOF5ptcSkYyUQea67dKtrZ9n2c1WLkYHP+
+QA7tZihx33WzMa+ngIud+4LBmCOsBWa8Ag9hTLZlErDoRtNdCdk5iHJa2aJPXDM
bdTv9pMoYqGHb2B4cxBSizUTqyn0qmCT9aIcbX6vC8C0D4EOgdz5NZm3RKy6aVNx
6A98FxcAXJSM2abTZnjceSuZr2HwiMtuhsZP+rKslr/pmZkv5tsAroW8LUddQ7G0
GNaOc1TCIMD0AGR+cpLQjETua42giqXxCQeU+KM6IkMDLsH9e9HpUBNHwJqpOgrY
T2WHan5x6JC1qo+qgu/Ti5gHJowgV+0bl2dUrZxsqrjuxgwYXK9czzEZ3RXooNj2
P//5BXAyM149KoPNAmBdLEFU40Ame7imD3Q82Kvel3Qngv9ws+YmI9PWAty0xahP
9t0ON91d/hvTReX3NVM2lsXNclI+WeVZLphE/IbOFHughHwHJ/4MWl08WNQqdrFP
LdJ/4S/Tqgp8Yh+jRkQ2Fp74izIPxrlO+ZQXkP6v2KDGohtLmsA7cYEBppNNp/mf
se1RppXnhrEoS7JEL9GbNirRgcHNyz7+kcrWuXDACX1RfgfKjRyvJUEYgABsiJMF
CdxY1dHPsiHsN/elUjsXa7nw/9sJceisQlRGTWoy6HIKWDpnShGVhPac/EzVYgEu
WSnxmPJx6scyW5E0HRF5OCHEN3jRq6LawAQnv66hCycYiZlV9f05huvtwFyIhf2u
ktioOFGgLEU1GKqiLFSPfcUglUIudGeM7wNwHuS288duAdU1bmUoWGzoi/jPR+y+
zHqUJvSOexvVJrP/jrWzd21lRwwHYT74pfnRDS+BbwY0B+eF0zzkw8jo8NmPM80u
DaW0Rx0o3R+ChTgy9kz7rrppA++E294NN0gu2ZlH+Ki6uRBDlCLO8AQouv5sCke5
ruBYYPV25miXZDcx/tTRGDbMMD0mSB1dPns25yI+kXWvT157ZJJhXamjnYxlcy6+
DOkbUMPXq44bZRsTEaN+b4SPhPJezxVuVGC8xMaLrKcrrOIC7HIOABkExowJPd1j
elB9VSkmyw2BcZ3S/2JjHW86Znl8QhSxwpqBPHwSPjYEZvFymqi4UkETSD5iSCSV
dZh+EP+zx+S81h+VPTea+RvFx3bmqx5YGTErpGQRnD0HVpVqzksmkeQjFnaabGgq
irGGl9eOeMubfwJJqpTcPFFPIAe5uLXcKMgTosRbGiAoaum/0GXIGHcoRXR/DkLA
YSCYX1KvjEPgJsizAb+UfjNkAv3J+3kcL5REZEr/wb0/Ks8Yv+SiwoOQoW5SDiFV
B4XscHZYVuJCm3JFDbs+56jBCEIDeSAYLtsCDVXd4CnaWbZBcNXmyvbdKffgGE7f
R0BWYybItGQtJW/E4Uc7u/WOY0CN3kit956SJQzLdQG4Tc41UDMs1I881XzsSmVY
TAuGtco4NSr/tN4jLuHRCixEqNH29zNTTm7cwFLkB209NltVNN3sx7Yyd+PBPU21
sU8cAR7rPQCslICMY4v2ynjHZmLn/xmoG3tx/Bl/+Q8yQwqu3NErfIbrs2s0jzJh
EV0AOvJQYex6mK1PsWZw3kKFuIIo1tDoI2x9UQObmjrOjgyOz89FodcVQwwL+J+J
AzqM1620/W7gXYSjqw3ZvuWYOJlmrXHxnWDng4Y6BMyHkE455VyfTnGYAiNp30aR
7b1xDnyXwSnUIRHQEGpGutKgUgdaGJag3DbvcYzYS4HTaI8Rf2mEUOSr1EAcITta
surqNprQQPny5cU0406Q1MzPHhNa2XPbLf71nfI1wfUYNOB7cHBFb9IL9fSSpXxo
m+hJFAkEGcU9L+GeWa3yBNpZRVUlaTy/GSt3F9FYGNEiqGz93slBnH1fC01p0QrH
TFhpV7e2a8trgvjjYrT8s98Thp5QA6fHxHcFd/SrKJjUQVW/qKxKkgQeb6AygVqL
rbvKoonrY3TZTdw1klVntHz6mzLNk/eWuquP3n7q/xCBnzU7piuVzmj88VTJEbeY
lh3QnwNtZB+Gt8fu4gIuwDv1N6PBKiu3vNLMra7uZ3c2pDEIimeEqMO1RUwX+CVg
SvTDXAcDUoKfsyCUnrWC4zV8n7V5Ts5hRJQRMbYDFXQhjPy9NZFcWJuohzH6/kQJ
4z0RWZOIWWutaP/vFqBRmagjiUS080pVSUKnbg+kyel8Cl6v2Q0V+OXEMVCcd4et
ZxpI73SgIYzETRyraVGde6DesUM9tymIEdOTnDNaMXUPtLHsaTcuthIYoOSMyrU3
z8IjRgCHHcynh5oQ8NkNMkDbnDiht8yOdVwi5K00bBEcNZzQOUnRMgfmoNFrdmld
h/1heb1zxJKuaHgHTpGSdg+Q5wT8XU6QUhLg+WGlSXg86Rze1bX69IDWFx6B4yIq
CM6jnOczLB4YqaBWBwG2v+BLV3/U+8i0GbWpqfGfLOV5ej7hDn4mv1PxTox3GRaJ
Jnp2VfE60aTAdNn7SNF+Cus70Wt6QP2PitMQ0tb5pYWP0xCrX9ZgBF/tV3TddVqP
11glgLddp+e/hAaNIpXYfGsFqHCdh1fOZaAWZS29bj1IhHMxZv3Mhb7ANIX+nTZ8
moTX1MEVLXM53EjhKcUh5zwmzDyvGqEPYGsIoaL6o/6nvltV/WWqS9t5QgVA21JO
q3YRaF12FI51qeLHQy7jAiuB7eE8AdoA3jKHobMoFH3pGO7H178/tUIAsFL8AT6E
MLk6M/vkyGmFOi7zwvGrbGZoqD3XRX8XlqojVbrAINfc6WsWndw1a1nEZkLxLi/b
ndNgxZTlrTjC2fal/AG8ysX/I0QjKXKnz8dZwx9Auct5ko9dWDHpjMGDg+dGS/mU
oSsqZLIc27//YQklDNqS+WSFs7CL0t45wJHVqKGAqdK7raRil2TaRFAsrz0p+9Lx
bAzfBqeZSd93rGd/N3eoKCjrpayIg+H35F+0wk/1oBIaYnJ6zByqxZJHfmqlA9F7
LyEUM6aIJwPfqpa6+rkYiFQIExFPnEetefoRYKr0YEDNplaqsyMokM+dzGebC6Ag
aotpgjf7WxJ/kueu0HdFpLTOh096m7SIFXaKqY2SQxYCmQ/jW2RFafRNiKuXNC/D
XrgRmQvS5Vnvh5YI5vC3/f22ZC3EQjpNTu7zmWi5tRt5z07boTB22QHkjwxt0oYW
x6Bei1m8WDNBmJaYSrnobfa4Lpg3QRJKEvbqa2A7MHbJL2s+kgdg09nB/hv5HlX+
PfSP6wnm+AhZ7Mg9hLZL+SkljIbVTQSpFpr55Vd1hcGiPgNYjdLFtXvE6VYXrnnO
Ltm3E9dxcVHZNECCiBzHrXTG5fcspLMXM8a6jdN9Ak9k9Xk1EktFP8COomJk4IZw
U4eCBSsH3nrvmM+xAa6Yj6rYBzmvU4rXPLyXDLPtjC4SATuTf8VSX87FFuLGOpkk
rt2fnbkEi1Rnr13+hsWqg8jWP0vPiFDQ04c+uQo4aDXVWQYcJFqwv9onltBffJwp
ar9o0a9Eqg4vKExE1WoTV9GoLdWI7hvqmOPz1DBzF/Rv/SO0/8mp2HCYybyWWvTY
Rs6N5IdWQVyywwH3sHmRY7vrdbJcvp7GXT3E0IYxjoVjcxYbYmyI7AoTEo3Fcqlt
Gk1sRJzZxygbw5z5R2tE1nBXzrNwepIpSXkF3n6WOFT7ypK+2g3zDL4M5XpoXy2C
leFN8+MwX4HzCa66th1JyJRZaT1HQREjPeMHn46bu04gEZhGz5y7QKsqhiaIyeds
4a1hwFa3pliM7AdpYjIHjtb6lBEs2t5dVkGmJGgljn2yPEHDOs6o1SFqjKL5CWvE
S93hlYk4Xrq+uCp/6dbLSelal3ykJK8IeAKg5ID1IjWZcz8LnmIH7bvr56BWgBAq
DG4ARKwzkY0dMqSlfsFJeRMporvxcyotPG1NXeI+Ya3u9AWkNRxGPtcklp8dkgum
5RmkXW1L0+UzMt7OeEaGVc8HtSNz3UluJEBTc208fSYvqhbYI7CoPLZjz9wSi50+
fev97ctZyYzb60KaUQRqa2JPzfkne/3Eq7adl3iyf7qFnoHLp4mNZYQpwcerLY/U
OsQIzOA08sf6JJjHyk05K8Rv6bq34l8RjjPRjT4xNMA5HLJa3XFGBceDMBRW0bBV
Cn+1MpXbj+8oVBV2ME2haaSMpF56YWjDs9rUMAPuvhNWOWGAAQAlm8ybAp75l8xr
sDHI5MIsPCkqwWcfN5b9iPqJiQfhhTvdsKvtgpj+lL5GBXjeq8/HE8RFBEwJHZ43
kbwn6KiiBGmFZUVbW4dpDZElZQ4ZxWKxgI/ri2qhZuUMasZLNR7O/TzvvTdC1Gec
3phLabYz70Wexf+1w7ET4E8TrkOoUH35+h/xxGH19Vi0q5U8exdZc16Dv0t/V+fE
Nz8+obSSW31iyHivpsryKXJbPbTV0/pjzgdI9Z99xfT3tQgf4nJuI5t4VkP+xrsG
PbLzFwJHzzRbeR2hS7tBGXHuh/bzVzSwuzbCiTMoCZh9F8d8L5VPNGevL69fekh3
0efstkmKMNeUtY3FiT2xfrgxh9uByAYXbxF2mgydMLLYQr4oPWzcPsWe1+atQHJ8
Uc5p+RsWLvfiRouJJK9it2JMMQ8Srat7YJsT+5tx392Nj0Kr2PPfH8KH80hH68xr
I7hbWFsxT9oD27clXDz5BGiAOSUG77jDCYZ96ee/Ypa6+A/GCXVj3NEHKa7aMTX2
Agp3Xiatzv29PRoaPHJXAopzheisI3y+BuTX+P2P+WIn267uLvILdWnSc3ph+p0z
gQMXHWtG32sQRO+LwkqhvczN2Kc+qOsnSizFCS+jbTNe0IlPr/ixgujD/h+5RLHK
szRJKiYeHrexI4FBlOMsoCk0zyFkZPtyivtwObR9GShDJSxkP9wL/nuY8e4uRY5u
gVEQO7hXiJYb7g9j4P3ytdNHwjtvTbdXucTyFXogjnV42xpisXX8SdFvjU3w7ljE
/KZJadGqk32VYHCTTnbMUjppkcZOMLbIvnB9k8S3jOwhEmUwnW8BckadXFHDiL4i
MCQy3cOG8EQHVRPdeG7Gtc3SCtzMAjHo9iC2dTetWIdqSbaXsMNwdyfiBtb83TfT
Gg31joyNq9p9Gl4pw/AuPJYt8+GhuFu+zeiOPeLN9DjuLKdselbbEVzmL9uAJ1GI
xzLHOtD9O0HP6MuC2Mo7rH9Ypci7wPCzMoKihFSJvz5o/1MU3jPxKTRASIhR/lz3
RGhIaErhqkAoaqQIPJ4Fpx2qZy9AAYxWts3v3JIvFvD1xIfTIqjjcdXcjNmVy7Zg
qCzj1KegjYDLdfvC2qWGhuNrNbdmS+uUk22YYV5sgKiOV44XMnXeZsA4vfaV5mQ9
OpLE5/delsmWfWs2GSRP+HrvEGel1TR+njqhjABFSt6cJ/19VB7EGIaVDQfmlQyA
H1xLMzp+gIH1TVZbZ4M2tU4qCYJxrnqrrgDWlkY/R2iQVGViv1qPj0v4dCcEgTs3
I1zbeOYUOsPLRs91q2ZxeqRJaQm9sfgY5w7yfBLAsNDCCL7Tj3dCyTOWxYn3R31W
wZaiFhDXIyUAeRV1gEF5bB6QZxRzMkwTEY/bNrAVdY1OKeC9Rqd/RHA64sT5Ya0R
xdmJkfM77zhS/aWg2SyWJDdjVJBNS4udJplkx6D6aS8kFYL00SmkM8NJfViG6vfK
a+DGwmja1hQgd8vfwTru8MKlbBTEtUUc3jREtNpFGDz01jYCcDPcggMheE5BIl0t
Vefh9MlJMRDSgmtr7Q/JszpMH/lDo8bKtm96x/H0ufB7hNK/DeuPT9W6Ygp+95o7
wA5BN5D2k0DUibwoDHipcTgGUjWP2R2zHAGfc9TcwSOGdqqL0XyEovTKkISqlz8+
Rd4R1Ns5+5xa8gAgekRnMxfRcazuTuxuncJQcwJUhIM1yNfb/D++Iqxq+m9rALpf
HYoEwpP12uoce5OWlm5XTlr69KJW+Vvex7t/hqK1LlefnIqICkPswuTaA8AEJRLN
wtARbkF+YPU0z5Yl4uIyFgA9gUnW2CewNaMP7uCGDP4OONwqOOLFxTtc04HrIqpr
Kws9IcGW8pOin+h3BY231s/v2shTQK5h02GA1VnhMzgn1ShbLPmsbcxDORIyWXET
VlOTUFrLGSSJtJUW5ItJyaoQptocLTqWMMiv4KIuDBLbjufYQbVZ04IybiXA1Uww
pue1iJFl0hsjXgLoQWHAlovWWsysbW2/OddotyRCOMDAHWb1RVr8SB3tBvZaEz1f
QQRjyVlWdhrNlFCbQdduDEsLzqNMFA5wvLKJXLzoXqYQam2yoJSEZXo9glR+H5jU
zHYt/n0SZgPvouNUcc9m6vgDwgr5SAH+zNfYGNWNAo6FwAd3IwyQIlRq6ltqgbu2
qMYuo+XTDR1qM7jYVGiRD7mLrH7kT2aCOlQTu0zHO3VgzO1S5QPkUPGd8qCK/sSJ
i25iR3YYjvsZI/4aSRGGcgOnG0lCGN5YA1q/Yfa33rzZl+Xcr5pnrbeR3NiYPgjc
VwPQfcYZhgz9Tdgbwr2aZJk+yeFgt85yHzJRM1qvwWBT5UMaphGWgvNCzejo75av
GR0+LctDmyoF6MEpIHgJgrBZiNlzWJJOmF1I1nGiaFPXR+yEDtJPt9LE0q7meYde
DT7ujlGfV7f/Free5w91Ud67XWP0P3iyh+vF5Rap24Rm2g1M3CjrxPzQmSprx4ll
QmTj/UGblbSDFqKubIprdj0harcbNNknZ8tBrHIbEy+dMmAhy558tyKzcyzomSdR
CYYHLduTQ7GFRSeRsUxuVTl73X9KYtC3COl3p1qjb8JW5PAiwfnc576FAObYjLVc
PRkedCXv/tKdxRgNzQiwD2VUkkWaW9k+iYGkWKBkGqDlh527Kb0dQ2Hepp3XdwH1
NfLVEThjgt5KDR+fHpGZqw3At8drpMh7e1g23E82dYZ3k4BQOiVW1jt29wr4lzCn
qoG4wB9b688t/VjBywBvuxyTWhOZCutKvN4gutggOWVyqWVSsnn6xbGCpdVxDMtH
hy85LiWsS8rcN9rmrBwRmcFS4HNt3WswaS2X0VsrOiaIyWcrEbBF3k7Z9K9pp7Dm
JYEkVIJ7ByK0FgPwwpqN/iI82fy7iQ3Kr3QSlWDQ93ZWB8gL1xfKTIi+w2weRVEI
LnfZOyFDoR9JAMesCE2moyfNeBOrtZA2K/e5/F7jZRQ4T3VEmo1FM3OFJg0zhC2Z
KRTrcczTFiXVZeA29Z4uSPI/GixtfkM9FSjFoQZDAq87Qg+k5LKzl3fjoxcWMvt4
uIET2kCVkSJM3Q+IPwJonA5s+11b5S1seYa4jNiGhM04+8E3Xwnss9GD8Eg6kOJw
JxzbJGEOQzx/PPscKudGiUjJnpVNnhRTPUMXMohCD8KGSPYoS9wpzZUSTKqHWZ2k
qvns0c9VrZav5wTnrJOwxKj6JODJr3pfuRKAaM+D0PVGIwmsygklPRM1UdT4lmyC
7eQGa5cnwopO+hxZ5PzlnP8G7Td+gp7GFjpHRwPxx75rChrNAmbD0Mqbadh7DMAR
mHEuCqB2FLtzhYWdHQySJNSPXB1UpdGGvmJJ9V57uLBATxs+Hg9ullf9ZaNn0BxY
85ZHe4N3UieYjql4d+M7GeUHLwTL/UG9Mn47mBHbkg2g6hD/s0rAlfh1IxcoLBGi
Fw/NL9YcYQ/bjgBECSQxcgF+5LKpw6xbRT+rQyfGQWx3OVwhD3ehhdMAfCK4Flpn
s6xWuaqU79P+LIUgPgE2bLLgj58fJoQ8ceiGtj7ldJzeHfMLMRj+VJ51UJgw4ao5
4QAaxaB4yONQv23l0sLT/4GH5RnpSO0L0dg1z6aLr0RHckZM4GaVeHTWhJjhANYx
xcXVMw557I45BSDDrYn69MjzdxPTFMZjyp4OOH/Rq8Sg3+0WP5H1yMj2PjWXq8Y+
+c5etf7KRXZQ2lsCxO6HZbE2vPFYJKsNcqSTzgI0cGPOK7oUXqMZb5bSicGjQbG4
bOFi600trZrSe2qxC+2QJtnS6lIhHxBJODCBLXK+sVLC5y1MV2bZMTTAQ3XA9+qK
CRiNcVD5KEEagMif3gqsChnsjElqmbLzMg1bBrFH2OkAXAqXi2uQnJs9V3xahxQK
RSsC8c52fnpwNGoZPnLtzV7bmqVClOYh0nW3UyNEGA+4l7Zo2Mb6SAAYCwaSTyio
uFMahM4I7HpSMdcjy2vMPqO3RVpB0oWLx7sQOXiVLGLVAoTZqOl61DqRmCoM7nYX
/ULk/v1sRYStNgJZlFR8GtEt2ZO8s88xXRYj6yN9bTp/rpSw6S8eCly8Wg8cRQa3
lYxkdoNwc8dhz5TbF3g2ckiGuOSHLqzpNyTS/ZFxoMB/qliVSKitIsCso2sux0xg
VErqjVM1qPsQOxMXJ4SLL8A4oZN4n/0BK3E/NPOfyS2w60IfMLFAnHqUn2CiwKME
F/OmVOtVDqA6gjTKpAOycM84VS9XsmtuoVX6XeIlcO109q4vdMjkEBGiSOPWPq1X
inhgkRSqrfvU3wtWhAVkdZ5Lqb9liqvSt0GIYNhlrIesJ29jwx6gqdi2Oq3Y3bPE
DyIVixQBy8/NZfww9zX+jd1N171E8XLPuggb31+qYnNOTtJv3oZ5QheFRNaXYWzi
mnnGmwO8ZNiJV3C35biXtlwV/kNNs0A3/Yt2oq6rnePLehTf6dvHhU7TfeiYfeTd
C9kmF9UHv3gofevW9P0M4isDka/fU/osXKwqZ/gAWWGB/BSaAILaL1wdlM93MAIN
s0LX8BZEeggnwa+orrm49o6Ry2nuEXTxxpK6uEa7rHhqlsIwhnf/zQJ5F0dfQ/xJ
se0VxGMxOhq9kJnHT+BDHXGRy74qHLlNsWiK3RRb+ZS9JztOuRyi8x+OVS4Yvypk
NvWVzO8j2eF+aAt0kN5s7qeCM4SRPGabulDyrYfKRlNvQlFTFPfOOTX6/FuyIAfu
niN1nH/z4trllDRJy9397qEdOyYkardGTGE08Jsf8pjzVYIZz+XZoYZw5GOmZ6wa
27EyWFCsVSjvo5djmhjMbtGBCin4P0RgvtmMlI/xy3+/XzIEeuIQCfEKFnGg0Rqc
QDsBvjgXAOvu9UMR623XsHEOwOQEmoTGgsaATsIU113ZfcGHPOVhD/pcA5T7SP4z
lQakME4rmsDtmA7FwOowEjJuQ/FzlrmAIGNxRaJNyN2+IY/QNYmVeegeJ/2N9BM0
Ew92eG82/fE/MxbNTdDRYYXdL1ihVSFZ0RdikTyv+MOu/IuXmrAZbx9MiN4oiuRE
OfZwlny2PMb6YSIe4DJAkHptCQ1nbCFJFOY+FqbFlRjzCrmhUFxjjn20uDU/ttX7
xMOHzw4K2CNG+QYIIAtAHxRdG7bGgAcJ4pNNFJZEZzIUVXm4dlZFoFZGqcB/fSmg
/1AP70czH42TR7UJqzL+cyXY5X3AijnA4a4SevOyfDXpxhAOMmBbRcXBEVhmTqCB
SXdilKNuj3Xh1KlGf7Hj283bsc/5UUvluqsU6Ja8j7m1alGZYlSprZAMevkkXi1H
QE+9jMevYaaAInjE+7hU/Sq69J8Via/Xt3TcKe26OA8qCN928Y9AZ0CLIOwd/Y+K
36PyWUvQL9b/c67vn6093adEsLR3cKH1ZUeKC9sozQwHSVSGCt+V/nQN//hBYgmu
PmeZButJZ05UdLhxTISi+eMPAsnHLwYnrjUHDWr6YxY02ZGBIORIFkL3m3va6H9u
VUKnlr9uY35VFnFI0K5VUtlhj+fJM7W4iWQ+YzAKlYe2CpSpDHlcyuIgSC+8WZiT
sMBvLxrPijbhtz0fFOSowwq3W7O86rp4NB7rBmMbx/WG8ElmaIrOQY9L5XFk/Nwp
QwXrtmIR/P5sLub3EPyGX0n34Fri3KbRqVC+8UOn1FF+9PvS6ajoQnWFpXjgIVVM
aRxde0lu+w/P5boVIf9LnoV0HIxcyvgmZYwUmUVUnCun2S6s+578toqyRzVk1fi5
ub4XcD7zEvt8PLSM/I4MA06wYY/7JjguuIvE7uK0P2VF3sZVevsNSCeSXB4lfhDt
OBObsh2eXMy370LEATNVVS26SGxQZeMlGPuy+BgBce/AIiAkkXNTcczbGjlnfnKF
1pHwUFQp7+L9zZRszGi/6wU9bry50JYURpEewlLV56+ijdgmFE1J4O4ZrD/oWdxf
rosdLRkzKY2JKPVHk6IOIrEJANgHdZKjyMA9Bg5q8BKENOI6H8hiyYDtKH1fh2qK
CJT1zOpjxok5CVChy9CoESVSeldEViyRj/oGnty+TqlR1OxePltyCdhPSjIveg/s
XF0T9tO3Wny3nhTb5jYSLNXBwHgbUvxZd8F00XoztjXryU2Ah/RUFQz4NiRwgLPX
QKwpdLyUj7GcdKJH8uluXBzmcVQPpJJNCLkYQR6np2Zkzu336uQlW7c6d4Fbfp2+
6NTiJKRmSgDOHmrSsKWc/dEhrurRlltKB5yQ87iHoEVgxp8cFVVu2SQUq1RXA/na
xZIgf8B7cR0RAR4NAAFWoo0KCa4WuN0ItShMVVxNKX/0Ni80082rG9LJwBNmj5G8
wYR4fdfCwfTnFXIdnPd724ahiMDZolnoZicYKZoDMQCFYjDZkc4NBhRHyQtnmzX7
H/e6MeMQNiDcLYePxq/2ufDDVSodv1j4RetKah0MNcp+4bfBslc4uIuCKjzJmU39
Wqyu59dsM51UCOgmoLDmyt/pE2mcM8jISkh1M8gUAv+jBbpB+oplGFFfROB8NMHn
0T7QjTJ1T0Jr5d8hlHlWBh1SsFnasSLSSyegcySRQKoXVDsTWWr6cKslkOttT9T4
/ka+AoIG6Nr5Uthaiv64qcUWcNndF5VwEc5RTddSBQC+9/PE96l1OiH/A4uJGwlj
XsFdvNQTe4wfY23+NBfF7TgdOA5UIQdnDammqFtfOSeHXMHEIxBFDFx2DZcHD7b4
OC9MxhM+aJqQsTs8KYJr5OjcX2bPZp2eHuO7JnD+5PA0mmVQxkuhPpudwN0U6P/Z
cnTjojSHX7stMNWCWlzDik8YxKa3yLU3+IWrsgzKQAP7fduVkTc6og4day5hRZqi
9bR5l1eWlm/tIHhoU1qHfhkHx0vDe7w9YfqN6B5+kcdW87UqaolPnkOqjdi7gAjb
ja1D1/BgxzTUcH8bUbWtl8ikLpG+nhZ/f+d+Qf003yNmEKeUp7WyqT7NB/rye4wS
f1mMa/u1IiP3z06RjtCAGyToiZWu/zRhutNvpWIycLP2d/MjGV8vVD/CvAhCBebq
GwhPNLE5DbL3zejpJFcsxNcvp0mWPEyn02G7qVeqRMODhV147sW3PLPMTe8b9EcM
5gj5jo8AtvlfAi/nC2ydHf2MwZctcB2Mh/r/8CeUoBqfipbrQ6bH38Brad1x5nZ0
Km49WycH6cqLKRf0y7aSmHyBdzuim5cM1DmvOvOIf0TYgqo47DeAwg6PeNKl8TPL
q1YETCJGuGpta1gupJvwLXC6NKUsto2ejc5p2n43+6F0/9dml+2eTyD0UCbKLkHH
jRaWtGISXuppWntlEr1BO0by9dsTHA1qGGgTGxZ61oNpd1LmUZDh885P689EWYxs
PmHhfCu9U20k8oJTdpHshm+o7f7+4T3Gn5C37J69fb9vdkBK6YPgNw1389nVz9J/
xIEJL3wYqvkrzkniOXiH75FuJ6MSEZvW2LODbEyZuR5vIX7r5TrMbZv+FlPPdA+N
YvI3iT1G8PzNVxVNescttaaRoTm7qma0FPbsA6ntqSn5sAzjR92nanh3bUWRJq/m
YcluOUosGMiYc4ZKgGdjm1/olEe7q6WifqLl3kplVZ+v+ANGoQwNjUDMPUYKtJwI
Y7RBCNaeAHHgXnUYpG0s0wJQdJ9LJzoGrK9nHRb8VfniqQswwJswiODBp1pq4l1z
nQDezOT0xI7Ifuk4DywnwxnstximZg/HqZ/SdS0rZEz9hpQV3kHaA0IZo/VSMRbs
vQ1o0D+LASR3C1E6Nr8STfSrtDqV0g+oiXqFrTfSGfSz5gEtOj3AkV3OMiq8C1oN
iUfxBxJzh5+/deBPPrQbzHebc3EwqiEiSyI6E3mLUX/kk2NJ8DsXHJ6ZzxJc4St8
4a7+XLW+cSODIafmB9oKZcvVS4V/hbdeVKvA7t/NebvtZvrZ0DPk8HqmpZJ9+kHw
q6guMaWe29AUkHkT26v9NkvlfmdBYIqkKAFewrDKXoIjkWXM0Z9wssuROQu8MAt1
kqY5O9/EqNFR2GLnYZUdTztXdJCBSglUM3O1/mabNJr6Jj15H0L6YantfjLJvTXb
kYaFOngLUHQ+quFnfsQx1QbG7xBnq+LiNJqiXDQCg69lVCu2b6d30FFMOF4Kt1QI
bouMJFeBVNhYG2MeoDi5H5bvejRFZrDZQYZ4snr4B8VCK1Dw8Y+NRgw/GrA2tSf2
WZM1GTbQIBpW2gNc/gk4CcF56/SS6G35F8vmVi3H2owYD6wIhYhARb97hCwzSALa
oDSZGtDJXRJde2GVPly4qCDHC0eWOUK+5UVrrP70myLE7JGpOUDhcb9hBSLR4EEt
Y5wTC1bOEpUNEtgNE+YqsGuMklIab154Z9Vo6sPijZXRU/a1B/vjOS7B/2hSK/wf
g6A825BZdKvpGGkPjjeVl1GRZsJRPHEMMDmWIKvwVatwexgeHXlV+RzZQjp7Xw0R
PTq5GK21h1mjpFODKVC1MI73Ct96HeVYdDTr4QHKfnc0VE2g/yeXS39+xAJ9h+0V
cNrtVURMbOOV+O3bE+OsQun5GqGc02q9omgnzCUqAqB7vxi6vfJYCK7NCQaOAGBk
dzil5X0RSOhMhPx5HlF0m/XtB6oZDESQnk0OJP5kHsP2p0qcyf4rKACyYVyRa8By
4oELyFBMXzWYigyk02wiMA5RxwnPvybmvvHEfgLxMlr9aPiw7T8b6JYuv0hYP1pS
Fo62PHK+zSpy/qmucg+BuDx//AnfhJc3+f2YV5Fkacu29g9I0pP5YBX1MGmSBs7J
P3CIKs60dB4nvUddDss5/i57Pao+eQx0AS13deMwlQFec4ipXK5yvPM9mrYYNXH6
QOhOGvO+qSa8S9Re9I/qVfeeWCh8dX2MPSe1bKBFuoJHgppEIuFFwTJQFt9tSPhK
BWjejsfY6nEFrYVFIYUkZmGykREW+lUcoDW4HWzQhBW6pCYzhgNp6lRSOMz28Aqj
37SH4XcsAq2HzyNDXGH/JtuRC6uf8OT9j9EF8qnWcFJDSoiSwZgAFdUX5QIr3hIA
MM4KV5i1JYmEJV0+yHShvYZPgIf2HiYhK+god+XzOw3UJbXB5I9GE52sTFOstMCk
Szg1cItuveuqLfgnpbhKrtWX7I5fmHGTS+CgN/PAUxuZ0yYcFhORCGl7ihdfGf01
IATTdbVNn4nibcuhK04IEekey+/rW9OXb0fh4fTHXLDGwCTuk0voMQ2hdyKPhUoM
oG4ISSQuZgzXclCy+vpPdAWHALx4RNEt12RFpRa34ug00Hzye5+eXhkxnliaoQ8G
/ZTsNdDXXpFD49duIMhcHOEmXJMp2hl+E7r5itQVD9fw407PSiCMjl21+A3a7ByG
oFuCJ6ZoSM3t+BGoShbLX2qC42WtZPFyVbu7Dcu3pgcuDfw+i5HUlmLXWKRdzyKe
uwr9p2hJjqQMY58skDWJpLfvFNXfz8s1OrfZlam/OK01hfd/Yn9kDjyXYqOSv0jl
X7D2GIC4vEKkFwZCHWxY0yGyg5qNpfPrIFnGJZFLs2tXU5MU+c4ar65VkevGK8Wg
5OGhDJESw6UR6Vmvh8UvFss8B4n4kIFmF8F6IqwC3SJPGVHttgs48EvA7YTraOKz
khSCtSBvtMrsdTYXFyoKpT7rITKxDsImVj07Au7CSV/41H00HZbn7RhRG6m+QiGs
XhyT+HT30f05EIXBJvwl51rkKUSZRf6sHeyDjhUI2UZcp6A4n6aNG3GswDBgWDgP
EshCEya3rTCqxF3uijTzM/5Lq+ojRCyMiqQ/aJ2L9udKsTQXpEXv6JyWdOLtg/WW
kVpLhIUz4SMK3FEbUIImBMet2dns/uZ3Jvvbwq0/xjzTwq1YaM3bWMO3ITbQa8a8
KTSOgLt/boHgX9T3f+N+RIBszPQeO0GlZB6yiE6FYOU3NmCWIoPX+c32Zi8gaelT
1LFdVe7xZHc6N5xN2e4Hof2nGl+K8n04Jr8Ne+Ex6Pq/1nJrnp8n884y8bRtHEYe
hNJSrlge1ygWlI0D2593ntmV/Z/3VZKEwDPs186AEdAarpeHog5URwGFqV+8QKKh
z0xl7fLgno0AHktHI8FRWEGTx34leGrpD9vNB0JG4ZIOSSLiRyi8IVDWoX0cq59j
oYul2OsI2c3NSsQr2ngWi83NxC3J5x38f3UV/NGaZ+5+VKdseFnozjzwN2gSW5Rs
SgCviKTJK9cGjbGomhEuoVTYKLUPJBRxiFW4ApoD8YM93rzBxlKZSWJHn9tlOogY
fDWgYfCocKogim5esvilRdAvSuTCQYbTzOrebIhDgre7gA+PZwd37Bszpsv/01+1
OMcKmKCqotr+fhonXo4lEmFQ73Xe9vGIpg70Q+Jq6uhofg9uusWnx/HK+EcP7TiZ
dyPwKXznV5V0ZINJg2/5XCio3p4au6iJtmhyOkerUkNcfxm1U5ki+AX5Z9kTgNaP
ucBwPrKHUJOxqkjpgzuIk2Tlvf3LR1BOhgDUs/GuNaoUgF88uuB2NJgNfBBSBhVJ
NjmRw/XdxYEk5P3OBKjTUidArhxlBOTDiOvD5d0eyFybtTIBBLelzuP/IL0bkmig
7/GTX7VwNPx737UrsxmicCzcoroZUaaMFiBKvfiqhq6N021uFfIiRE7+QjrhurjM
aX/SvuY/irEpG6xSX6heuQzQS1GTczPlNmM/m6fWwGgQRXXrKZHKwFPGbYc0iGyg
lQ3zx9jtuH1UDwpsdUO4HQZ1SZcarOgrofPblqs8yLVUtrQRm5ZvH07l7QfmNTMP
UrcHQZFTnYdXRKBcNOU1jQ++CqM3925h6++sfR/v3Aup3BYoOdw9UuY/vv6zwSV/
Ot5Y12P9txOHPnVV9ho+MVc5ZtpI+yb8rLiOMi2GxKC0EfCMDwQKZU5cp5FHZb5a
P2PefB1YAvg3W85ahpj2MD+QwN++x3AKmcNp6Wm9FybR5VIAfB/Dm3OcYAd2fycd
6Tj5wlaxmctS2VQOFv3onZ8ikYBSeMgTgrcHs35FdmLVuvSUhHcSTmRslDG6ZVHb
Km5rn81OdDZ2yT+eBNvdIHATdYUOu7t7dZQL9xls6d4kzGsWpvdf2UBjKiAtPKsY
0TYXJkHu/gt/ss5WRn8AAM1BkCHD88j3CyD2HuQHnpa8RKE/tKVYigaS9QzhO+la
OaY1ySrF8jZlhQm81gsaRcfIwCwDjF2mVrqccMZ6h3B0pubOgc4nSH9irFblQ59L
p6BoAtWkEzn5yR9QiglYxbvCh/gp/6O/VFYY3TmbazbEY9YT0wutyMM0rIUrHY6D
0LKfcYIKbfj4ZF8w1bCwbVeZwbUX6YsZ2e4NLe/1MskMeelk7e27G4RSrNUgbx8T
i4Jc1yGb6m+AK2sIcc1XGYwW6/ItXgH8eVaEF93YZX502edkcVbBIuIrn6Gv4MwG
38s/7LAw5PIbmKBIdITAGqn0lzCeBjpkLQCYMBuzLaGSdwMW8CVVkjrh6nU4fuT+
KzaBHs/j8kA0xXj7sUDazc9eMOOhsbraJ4THxy7Bkl+75g3dfRkFeGvOCxhi3NY5
9BI3NBMWYBggrgd3vY/+762sUAAEO/x5xfPBvX5gB13+UqfjZZtcZ1MYWHYH/wXJ
sdwFUUzZgDGxqXGOkh00X3N/JFK7c+EaZcMPBvgdJBHpTf+ZnpmWqqlAs6IKbgkD
XNF7h0KsKxcvomgQCQ+i6v14LbMSuYESyB208S6rtTZEjnR9W6Vg/urSQwYHbUCs
LzOp4lER8vBnysXl3s6TiBcxAa/bJSlLMuwFvrRBvTPMat2wKCkLNzwPTmRgZ6Hl
/KcwJ06YvbK/MVpGaZRZthUwZ+xZAXQvPozpQk1FXSCPbf4nr6lIbzoEcGjvHisv
FoJ7SNwWZ4bTL2RUQNkG3DqZxNJqtlxz0cNo8oDXHU7PErwA1yIMOEb1hgseh5mG
wDEYjv9m3rxaN4QRG1iPK6wpHtQmk/FgacoytxuJIcUAcRNacSiIKtdk++EIEMcs
s+imxuJnA1C1Qt4bVLyXZFAPwVjIb5Gn6R/s6UvNKlno1BQNFaBB5CrxcedeLvoj
iTdxjVfSeZ0cKqdH86y/qk8k2MZ3tdQvxj5T6ZGnv7N28t/7fPcGwmMZE9OA9hHe
enkyTVIRP339X+TiW3mhzg1Zsd5vb3rI2MUeK6YmtTEwlYd9B7Ibh1hXG43HCCEs
M5y17jRQHrCdjN1v6M050wgm/0g8pkC0ASHTdRF35nPvxHyWnFt72mcmema/DIHX
cAuuG+gJfWFkrEYIdf6V+TJJGz6Sb2DYzRqL971HrzV4moTuYmlS3o93Wun5DDpt
xAPR0usC+G+DUrLF9ZaqE2bl0imce1DNmI9FfrFEMojjqd1MrxK0TrdJYi0qvvBY
P4KfbJZy4zApQj1C99uWNVDFdYUU0ZpagDi7kezBAInvD2J8f0RkpVDnBfI+owZV
0WWgCEKECTGCjDYJhmkNZUhpd0SMpJNwipCWfpjz0m6Ty/E3i1UFkp88QUD0pawC
eJu1ol8k4dLZ6w5mYvyCtn5j4ft59MqcbCLaMbxYRk8ZRgy7GwHwtetDxGpdaOIm
YWaTp0vmMp3aa0yVElTpMaSzK0hMPKj73t7XMNjoxFOvwRCj13z8LtB51L79784r
/nz7TLBeG4QSPntYqV4kldDevzYZcuMoBEraDMXZQWowJ7nCP9c1f8BLVDCyfAIH
KdAlQmK3NV411hjQY/uJtwmImbPmgac7CcOm2AoGsKwn3IdGHy/zhfVMaTj/KnYb
rENN6bgkrmNg3gLSnpRSQGN2fAOXyXBORjIQqr/gI966t6h6kx6TDZLNG6QjAUXj
CNtIyCA9T3NNCeW9hr5R0V+RMXbAy4ILh5aVSgxkQt8lwJVaJcgfhs66g6Fa9vDw
BVnZpy4lzS2jpxNrWCVpHaOE8LXFm+J/B81BcXKCjone9tolaQJf9ZLkNIZZ0G6B
QsX/qbgE956g7tYZIu0UvmIF5qKWFAuIWf9aBcWv+GeWaaJYmzhJ+sYGctax03Of
YnfnCer9FnuyGlrhoV7wU+h4KYzwSRzW9x1XTMB0aNPCNjGuf9A42LLxTi3e4p9O
Is34GWBwc4GP594XLLml1DpTZWBUdpb1Lg6NbK9Xbb9xqBDJqUxuVkqN52tFF6ME
akXlivRfis+ymNS2rt35IHPCxRWrIkXIkq2AWo6P5/3oRZZZXl47ui/G91qluZqy
o5ZlWcrPmcevSJlE7BIN9t4zOZgDk72LAdRSzeRc2UY+gXHFU2IKPSB1QxWC4Wsw
0HOW6t8fxhFlBcNzUovvDxcJvNJszYc6XFr6j9T6dlGiURCBn7zX2eCaR6CQPjy9
6OKThyQimVBt7vcK46NjKIcwkqeKclS04/EnpnAoo/gcHN14R0AgushZCv9ddiGU
JmFo1vBnF8u2BAHyCUJ0F7y5FqhUCozyZO+iV8blMvShd2Z5XIQecIW8LnJiiQUQ
droUHm3eGRLUJDMFL0khhCUfqevfUQTlgxdfQmdddg4+TWBDlEN5clzv3cQ0tNeu
n/G2pJ09huAUV9/icI1gYQhqZz8xL7Hzwfl+DunxYptxyvU4GXG+sIMOY/1JaGZY
ntIV6VhvG6yubR6IvaoBuFzcAxEtSrA64KAiAJyVKhrDX0I1+aUbHs1Q+mqyGFNo
yCobNoGQiMOuq6nA65Ylx0V/aAgVUSgDkeg1REQewTZyKwp9yS6kn2hTyLHFRUUj
/AF1OoRjZm/Qei3vHUqKnXJtHB4O4/B9CMRgg2VWiu8GDIw9kZwUt7U8qDfOSkHB
iv7dKvLER5EvD0IKJrY8CcUgq1CMCPGgl2jYfIrsd9aBIt/Yn9QdE22uNs4m1gSF
3j7YQKiRC60LfUcIEbLy5PotbJygVqRqNnDqkXrl/miwfvm0PkvXJvLipnK+7Sy6
bCdQcWeVVq4oAvjrgfWEYyNQLHAAIuomap1FOqT4f0mGI7aVqO4KOJyT+X82erb+
/7xSA18c525dgUDzMYZtXmQ4n+7ARxVzXDdKc8FQ1liNxLY+Ze19BIUYvMSZobAh
Pa2gd6xarDQVjCwPpl1Mjmij2x6oesIxA10ucpXOxGmJ4iKF4yNNDBFMxlJFDSm7
Cw5S95a12eNYrR9y1SIimvXeKX60D0l/KCvkgUbaLUzVyDt148UWl5J6N+4V3nOV
g3EfJ6i/wSqPHijQgfit+I096Z6hGGaG+mpqn995UO3aqARIycAnl9RttQ39vwfR
FowWKpX6ELlnOkl9r2Lckk9hancaiarupOscamfXD8ojb1FDu+px5LZ5hhCCgPGH
qizkdvtyZjeVreQ4+vTspsBIxlrtf6juAy/a6QN9kejFaaQ6rPq6DdjYE5rffOnx
BFJGzz37HFokSt19cy4wlBRhlVASlE6M4NF9GFeru8AMyS2/x9m6RtQdp2qWJEXg
j7vG2svtffvNuufTklOZzD3kh5StvpVj0Z5WVyFwNmTjp/EejqAaTlTBI4lEAyE3
aYJ/4oP40Ik1uRqD0Y6Okv0TJmY9Dm1UNwN8zjU4xyVMZOVHIc1mdpMLnRwrhQs2
UtZwarsIHqh8XcRu6udIYqtY2pVq9qf51Llc27I5kk6e9mKg7xWWs5XC95bfHQGI
xq8kIWJJy0HhqnDrqAbjmlJ5qcpUA5Gne8JqDt+C1zcrvixJsawRJeSu5AAQnLZT
5ckV8qH9ORxXuGxn58Q8i4mtiN1F6PVapCD0U/c3GihL5A+dYdACFaWyafhUxvjE
qTMCJcYd0plPzGbrm2ddzGqN+y4t2CtBTyOQN3GLx5MfF/BaN3pF5MxlVFlQMwUm
sBR06AwNv4/+AMdXGPx5JzH2OXB4mWU+AfpdTH8mgR/e7zciLcz+aJHwuhgFJQjH
WFDVyXPrhw3NKPegBieE4zH7N9FmHaT6EZ9wlacQ9p5RTuvz6zJH7eLLw20ytt8S
nFnz4Iyl24LfA190EKH2i9xg5GTLBCI22dftt/oWeEM6fJHVGi/FODHbi+vYOH3n
FtetFIuharK4dGWZcmYcThTuAXU6zotLF9Dh44ct9LbH8i3SkBrDalQhwe8O1vLR
JkbpXfAbDzcxhHnEmUz2bTNp96LLOJLQymcz26wJhvHO8AWMVUyeGSTMmBAUEKFs
jx4lVhVVCOp9m9xtkl2o0BHY0PJiq6J0NAaOkH3sg5l9Z3qdaI48uE9UJOorGKxG
UKxqHLqS884/zUaVSfKTtOStKWm3fQqT09mh/7w3nrdWnamKzNe6Y88Btbk0M2KL
rE/XIJGbGRvPZWQBoE2RnP68k/dHayTJyQXCdrpiePdNWWHYnh8lCXzhbuuR4RtP
Jp1R3Pbc9buI4TrSiryz51xTBPxC519iIMlyeSB6C14qGEM0tkTM/A1iY0Y71y7+
9cLtc8RJGWqeRYTUk+7hhBUhpx7lHlv2GeY5dqLcFIDsaQnxN6Xz42ICQ3wbnw2/
e2k6MDQmYRALq+wZUtsA6Oe+WcqRYFw9jfxMsXtPdafL5sG+5Vwuz/B16jQQkUTM
mfbiDgkkF0PVUkutsT0yyrs2qG6uqIjilfJE1Qkljtepngyk7uJZvwn4GGUE11S0
tbuQlAjrDLpGgxFa4nToPvy/fOfn3mrJ8eR0X6+E/qLuK/LqysQcfA/HK/LWame5
CPsc+dMu+otQtQOg3EJodCy/Hm2qeSwqXfa/Wp9tjSOD20a2tc/qwi6CU9z/qSVO
6Ta3oMJTq1jq9bWNUJhZIlZnOvcqL9yl+y4bsdapPA4EE9V3Muqhjc011JaKSMpU
5VzDXcsmrZt5DKv7pUFroIS0jPz6tIqWkIytqyTI3K8VMqs4/wXmlRo16iJN9Yqe
gKAysOSwV7ytBjIcuGVZSy+UOYxXm3j7zqdJ5g4l1ffLJgD6SPiuHnA5ipyV1wf+
P7GOTL822vzdVDxPg8ZUahYAcEQxLBcWdBUZtXTr+RgmGSvzooCzhkuxNQkXRc4M
HIWYirVGZxUSQztXR3+eHmJ2jzFQN4AY7eFtD1+6Ctqo2BQ3cyjC7atyXzmeb8iL
FdvcO/ptpBPrBSsuiM5yj8v0Nc4BOyBc5mKVzZf+P+hY10RlKG4mGHWJTaFzuErZ
Vm2eAVPSI0CwOvugtMiTsF7ujzpFPt2pudy0geGfedzlpTKVYVkQ504M540BZGBE
GnPV0oGAJiYM0oZTWK3kjmbu9cB24s7oUrUAWn9+MNuUy6nYCrJiwzA+6wmD9Le+
wntfX5Qg5G7EGrRC6uJl7maE/XmweQds1sL8ZB4+5MR4dKN5ObvA+AvxavPzTlxw
3k1WG0RVxLkNLEBsDT8l/S4r3kZdh/K9xlm3EgC5WfNY7GWcjyWxHZxU24rANRQ4
aNlCKADzwFtZmvMYX3eC4Dfes3CLu4kLZAj7cNvXMjAGPzeS5jHt0iIMmmaOTonB
6VRNWfqFfOh0ODCQj+wcB4B/E9T6x55cbXG4jMLXYDHMYKwG8eG/tdATWavJR9WJ
znEptdwSiQ3Ec+MRnlOuvdE/gzSMRsf8OwRPGVzQD80vAmVv0qwVdcHbMAKiCbUE
1qzXgqKxXh+B3aFJ5bfVysnbkMQLicka73wCKYcGGnq6YihROr0D8HSMZQfCp2nI
9BlofKX604ghZmihVvLA0LDfiKi3DmRsUz/KPnhvEZpeT+6iUhAjR4EoCRgybKlt
EdxPLypLLmFrNWmX9uOS4BK3C2rx0M1bPqDDxHKesbAKlWKE4E6OHCUz5cykQWWv
k6dPMTdIDcy/zhq0rB2xirOQ+0EKGWSTswfHQU+ZT5zkenuO0FvlRTNho55s2eTs
JeSgkALvRM2uyC46TW1UjiqyVrOfEmTm57RPPpwnWF7/UNViPE3KS/eU7+ZzxC1z
j+K7/S5OA+hIJLXfDpNMtSnZrppNw6nNnO0smJpGjkdpZLtL9x4ZAuFPvfcUoIBS
u5Xn+xPW++X35o0FHJWH17Mm8tULRGHs6W3u3sAfMkkNJ9xgEwNU5qxd616gJG/j
NGoAe+10z38UO2Rb/R5+Dflnh/tXUU4lxc6RlETncQmr5fs0964S3Yp47k3hd6zH
hVFVIa/gTqkN00fF6AT7Yd+aMF7M3MfIiI/5yfyXRyfpODsztc5H7bzfG3rGpnXg
0zyYkGSC2r3QwNI5y0cfFKJr1PjxjhcTlTXAXBxL5JZBs5UpnWVZcqNoRuMAeFiR
Or00chL1C8RMRm/enW611VvAysDxsjnOLA2CUenFIgO76g5IxX7OP1eYsqKs8qhe
QhG5ZQ7UwJBRiwxbSBSLS6MZz5Udo0uV+5FFwmNKq/AwlP8ir4aeHDvYWqJoCWpP
Z77/rq1XeYpKoMmDWlfCS0Cjt2veEMEaM4gYozBqTuyBX/+UP0cOencbR6Tn93me
0G9S9+oavWL4PfdZTMaOVsn+WnU2H7kqfvb2uOM81r9JCuV1tbpPzSjCN0nizT8u
8TjWbeLe64fkN96bA5RX4cb5rqIotGQCp7YqKy8rFQAJDn2J6Fma5fCjCvTrRVoY
sO/HMGOp9lIINEjNWpIjATdJZbMHRujMzGaxF5vNhSrro81EoBbPgkSrWH5SY102
YAGO82oFJlFJGFkxhzUObTC/TC5/iwdTA9k7gPHXBYK5Gv5ttEHInBwHQhb6V1aO
LNhU3GIvI0d0rriBU7D2Kzw5iTdw1Qg8875Y/rKNyiWI8OSMImzRA0ET2+qYEuio
/TJoi7lFHa4JVs2Z3jbcMaP3p4JOyqiUhNJcN78mxapkm48OuRRcR8NE0C2KoetL
bEHuHlLfvK/vzicOUF8AWw39iQnzzUmr1Gl9DtPAsDzvnl82mJRDPDna3vzMKiE6
4CVqrRbBUR4BOivBBrtUQijBEnPIjjd4VrOhLVnNI1IWikAFzAo7leZW8iE3cZXE
X6Wr+SresBQNdnyvmuVJN/KEHdINfUMR6VwI59NMyCfhXvJayIECOuj43MXi/MZf
kefPCXU60k+xLHjef5GAEnsYXFTwPcS73iAjo8kkcs8LeQkFT2QQWpkz4AxxZX/G
gNfZQ8bF1/ByyaRpWXgHZq0PAiNHwYbt6RY7fm6m/KwSPv06CxvgsOpX0uZeZI8n
6EBFdvTlWnVnHHA8Pz9jXUoGlYWy2EaWTI6OddRlYIhGHmzMnanDPMxOIgh7MBoA
SiewwbCpX65a7SHmI7bLPBt9VvogE6+JbF7/e2sGv9jc5hlAKUj7rycWrGGpFMEl
UHSACyPuml/THJ8oCnGmdQsV2go3BfhCCumkeGYetyNwJeJAjTj6t5jUE2uqAJPn
CyQq//vfQBYhNuGLdbkhGPjrLy/yX6Sa8G2CsiTFqGQrCS01RfhkMQ8+3bi6d29I
Bpr+VOiDrxweyeuHazk1IdaRK63mXA/VLq4ZCvdwkHPto/WkxcN5mDnkzCDXNcAX
/iAJcsx+Kij1K6k4KsQWNLLjmZLdkN04WYmklZBxRhv1gS+UdKreD7zVPqM5oEqt
uqGZedounTBHz5FjmAwQbHT5ECpHpwvVHuW/CQ8roEpkAnkp1NXINTpM64vFxuGD
uKDkaVErtT7ncfoKw0X1z9GPmUYH3zNUSA5Sn39KtXBHflvGDuS8z6HKB9qwc8GU
l1M3Po8ujDKsN7wCIllh9zNVDF+AUL1GH6o8ZPXZIMc/ytbCuuuRVyDjRakJonQc
GyF221Dq70QQzPoIZIUKYqO4anOtwjDjBVsEqiKO6GXb4xu+4abTBEeEwfjjWyL1
DqjaJxINyK7njTZXR+Wf6dhaCrwRhrLuO/SsO5MHIiSl3SMUFIIavrzqh4WDjRSV
/JRL2pHVjOFZaU2/v5+k1mzFOdj+9vkFclpZu7tIyebJncEIcGmcU9PQPshiRBKJ
rG2OJ77cKUj1l3vtMUhW3uqiq0etVru5rZgrMuhQ1RrHMlDMlXlwImPJ2S3cjpbR
ZzieT/cH+8OLz6E15haEQXkSjEgvwLK9+mnXEIhUyH31GIgExgIJ8lgQhTRXY+rK
A6akW0E6OCqjCFlDUFL+rw2SBDj3Guk6hbf58VOV6mzNZLE+h0k/p2wkeSme0Pkg
pI8O238dLoNrsu+JFMY9N9Qx7OKRDyKC6OfhBT8sx/NNWEn6kIi5OFk5SGl3LYas
zvS+ckq5PM1PWMdnvEvH7ivCdRN/vUI/XFK3qMz9yjJzTcHdqTSFXCoQ5L+Cy+o5
y+qLNcuk1fF/3p3yOd/lwn4Z7PnBp/HEC9v99s9ilkuJ98gJkAJgmdl61oMnjcwV
t7O3DQpvDjAPDWyNZXtUywQtABGOJFT7PJAoUXq5AW9McZVcvrksOyNEiPUetQme
0zTok2KBQWH4rJ4j40vMuQuwuBQXV1SktkbRJ7zyYsd+r6Sr5wnQEFp3ne1P1rzG
FPwYVeBkmHtFpsn/9vo88WwfVJxeZqmFXllgZM0IxE4mxmdXy+hSxD7eADHo9wub
RBvEldum/EAh0g5ls++S2fIrifVVBjRUu0iWON3Qyw6WoOcW0wtDqkYfouQCq/rA
HoEQ4VsphTL770SnNYr+ctbLSNDcaXcysb2L168qdTg/bzZX+xkoShxioSgQ9CMs
pEYFW165RUgNT9aXrtKJsXpjy+vniNha3/JBqDBhNsq1/leMA2KNV5ILJbMtJqy7
v0haGQ9NdSyu2mw2g9ZsRDrT/KyBm922CHiipjJkDve10yBj7lWEN0Rt4MqYfF48
5AH6Ds+QX6s1uibg/YWg+2q3rtvP9cc0hGwCYqSPi+LFwsVsIbayhccBZYKVbnu7
FnatkDPYp8d6g+70sfpi0c40l7bi2IjyeOgu7WzhbXmoV/Mg8lCx7sHjSS49PGaH
Kg+fTCBVq4cR5bWqNVrGNxqXRuocE9wF1CXhTATl2cgCtKDi7SSPpm4oDgdaizEt
HGL2eFCU41EDgFQNvQ2eACGOZtqjfqOVHp+iH6YjG4pKshQZkmdefx+Zdik7SBJZ
6ItzBfXg1bW2mow8MFRUSwxXHrI5vreIEreDgZgOpskDrI0sCAE6H/CSTPrmp/Yg
pWQaVfot4elcpcliHhyGl2yebPX+R/telFt4BxosM3qEJz/7M63dIOAg0UvGQajq
+nCoZXXbtNWKY1Dotrp6L+k/WcInUwr0E1ZmiCJJJd+9J9KrBz0yRhOeKGoyvCuz
WPS3FVWAsWNQaSCeels+pFkWFrF/whl8xw7/Hy9I+IRiT44pmWu+vlrs7empIkFa
ZZJEEMKoc58SJvjxoPL0pNeMZaGmgMAoX+PgT+pWCugkWj9kxbi+QBOC+EeSFOJL
Lo7KifZLJQPWyJOwudcR0ihAq3WYp5e1oDkf0V8aJnyEj/FSD67vrN7dz7TgmrZG
VeGYS03xtmPa7NhHf+9KMmsI2ztznH45kD4I8zpgT6RyH5KuxMIqU4nvAW7QdziE
+Omr7DxpmwD6R6DsF/Ez6/niOgtrDMWXVh9m7ga2oyZtHQXR52cR47KO6sTWRnyO
8d1zsO53TeeXbYiS6gs32KBqH1sl2oXsjGpVEC0wBoc5Mw3CcCfSQkzsC8/VMJ5J
nxBDM1CXAFzpQoQjHY6CZbgMDVDVoXdt1U0TAQ7tKMOBdnU0bkCiau//boCNQd9n
Le38ljUeyQZ19cjSWMV/mQMDvGuhfd83AmpJ/gTFc6UlFDYsbGT6Vos4XgniazuG
/FG8HOMKnI3uPMVeiDy+3iR0pUQZy0glnw19GrbuLakCaHBVcPUOudtVcW8C/jVl
bpvVkyhm4Y7P83nMmC0dPsu7a9y2JtJZ7jbbb/PWwit1TFxva6lwBIriMYh8ROSe
Zi+jf/iZwpdr2ZnNP/2H2HPX+PN7ZlgCzHHCEvyVEr8zBc7wTAhR+1wbQHPRXjax
fTMHoJC0QZtFinpOJeLg7Skey7Y5cbbmZv71pbkXqWWritiaPD4FD4FQn6mTqgXb
X+nu28eqgTaMJg/M7PQmOjCnCDWbSBKhQb+pUFN43PMbseqbeYB/Xg3gh4xwRaTj
vFh7Obi5K1O8cg/nMTTaDRt6QzG9Rje7tFqEEgdYDJGH42x28axsPT1hX8x6CLIz
L/tzxcbTQuey9JNNpc898MehHuXbE6jpmOY9BkrVN0qLl1mknBw0Skn9/Ti5OdKP
ylyXwIO7CQzlNIWmFDFZco71kRyU4t+ADFoDW2Pe9MTCqZE3COJPjGVoAsYHfrE4
Do/+ABoz4+nq/+lMsS87bMOZ7An++RwrbKMABDlDOFZRIrTyLla5tPX4Jad70ZrW
KRSzrVF2amdFEqH2wD7qikKTD2skmxSpylFZD/gcgKHPNSPVZlzG8ZzTW/DZtev2
CKO5SwNUwUqzCzdWjhdJPyTp/B3Fj2jIpN/Y2l2uRI6dL3fIIDIPw0J4VbY+4SeT
vXaUpY/dIxqfpwUIKZs1Lw632FJh2MThbe4lW3jZR0bSudbEDVpgZa/NiE1K0s8H
UVMyoO3/kiH5B/VnJgcJUDsV1lBz38Vpz5FiXnZuuPbBhvDIM2RJFHqiF2vop11F
SKp75YnKO62TW5urHFRAzVMNg+Mm5m7Kq86XgbL+aDVBYFbTSLLGpk7Nc1H7RtWa
k/KVlQVj2L5+MZDoB8EMKQQ31VsiVKdOYLAg5IEQNddTxwlQ4Vm2wMaZo0vdhH2a
e0uDwJHo8xLY7Dswi7IX5I507ozroS4gzs+T/YB4IkZp8f+MKLA0rDu9cbVJNKO5
tvIESumPu798XFlSjFvw0DpTuuyPzmoMdY1a38ntDiILPIhrreC5Ko02XEr5XJkX
zl08F2PXj2fk85h8p7kDY1LSids1NsQgjkRjjhA0diOv50sL/2aQYUuHurvXg+aR
Lziu9tHBzuCAykEeR2Os5A6xtigzxJe5q1+KqwLWqgdUx7eoWJi65F7MWVBkGqf0
8vF8wM5HVJI+Juax8ZhLbbpPdDs8Jc4jo55NBqcf/JfzTgNMADG77tc8cyQT0xAl
gZV+Z6KJ/oIwndAxCHOOBQgZIEZedvmXdbctwXoIhM4KLdVouhfKUI+5vhXgQU5m
V2VDuJ+YAFTn9eYLd5lP78Pf1Iclcyfwq5vJ8244GP9ksbEkU1yQPivbhZORqe4r
Jwq4o96bXHbKTmdRnxAGBFl3bCFiGGCvyjig4YZubA6WD+fCS8Noj6SXoWWm5c7D
666NqIQzvfqBhWlYiMjKfeAfGk0O0GP1TgOoxTa9/3MLImC96eNE+WNjYHlvdj5t
FuwQ8xcM8HtNfV21M2B4U6sl2veDQ2Ngb0PXP9vmUfuQedBFWDsfXZraFpsGui1w
vxlPNR+eiRZOrW7PLL4bhDLWdU0K9yh38j6B+/OWZJhKuqaEEhSatk3+3RyyVUhB
cYxqLnwlYZ40OlMjcXBA3Vd2iDxLtvvU3TxjOctMzap3vBVGAYDJE5kRMsp1w4FS
dx3jSFqqRl84YzORqbieWtE657EJjMvVoKSHCFuy7MTWf3kaS8RVmeksp/c/1e/h
2jfHkbuk5bfQ2ImcFIWB/h/IFq+LSS7oZmn/bQGwm2+PK0DSX4rPLZv35kGCiAsL
UFbBWlK/AavdarwVX1FVWmYvjOJCdR7QIGg1P5v5FJdyQHRzoRJI/oUJSEEs2XlT
bs4abYX9u+cG1NrP8dPGc0JAQqrk6bO/AA+C1C8h/6z7etsdi8NMSdbzNGDih0IR
Ts7G+QPko7WLn175x157mnIYfXVAyxrqrwMGRg3aWOkXHEgonBkkDuJZSIb1fnfE
a4N6hisYnRozPJx1Z6wcPu+qZB7QNUQkH/pzbYp4ucaNLfdtJAvhyjB0uEEF1xbA
EEH0PREy8WxJ6guVC8bhga72BXULunxaiSyzY6VITMjZUkBRFZPfs+ZHTXCn8cvJ
qNWXauqunfMlgFJqrXIAnJdgT/0rsp3P8SeRWBRK5xr/9WBy42/sj/6ZOl8nIsLG
CRriSQ/jSBHE1i1J+Hfpp69G+4aWMQFHlPQDCJ8EDhQ6KqbMu5YzrvZciRx589UM
rFl48kFt+7G8Dd2/5UKA2mkpmIVj0lTx6zI48SpvkhSAvh5ya/8Dsyq7S0IoZjB7
PfgwigTjHlFZ3tT+GTt6ejWSnfvjsUL/FNwcBxuBNBj9GwZF7QxfHrakKqGtLQ5G
zm7oTtwakL/C15y89fziZmZ0VKETphR+QGcuSDG7J3vhLhqm13jxLs/6E6dZn8cC
aHG4YpCFZmfd4KdAQs0sxchCsg5LQxc9JDlC0puV+CeeyFFEpUyOFgmOGOOVVE0q
uLc8/2jaY9mTEzUxvgBQqTyjaK8P85sBbjjVRXSPhHS/wy1PY9suenNbEqHieTsM
nNQIOHGhyS93gWIBUPZ0aqDYgaaD453OO0HDuWCdRVTwQssRQwihyrLWz9qmtBK9
fS4MxQi3qn+pfP/OuzvuWal8R+fMjP8Zatpz8O3IIE2jdOyY9DhZorkK4Bfm1N82
MvhYSUPdtCCYHiIGr8oGqe3HUO0a5NrL8I8FHqpYIEKavSkyrmJxGCHY3ey10ugD
aIM5r6zBnBB7xAjLMknzRfyBhIjRy7VDimAiujiHzeTkct1m1gBnsT9QcCVbKd7h
1ND8QQ2HFhrg1DdwsAF8EurqcNo/MD9J3H180hTPB8gtDPmqWKL1KwT3lz64Aa5c
WLOXLbJVlWnwAr0lU3Hl/ITADlKb9yvpvdgzmlIUakkpPzE45EU8n3SpFwfRYVGk
rvldQxiJQA5+RBckbCXdWPRgOkFPGUxjJRVH0yryeVmg2Bl7/y+T+sGi3ZvG1H3W
DGdvxVp7EMmweZihVwjlEsOeZGgKPqrYWyo6NfwL7kxNvwPkTWdrgYcTqZthfcvr
xHy3uDnTKA4RHobUfEbYwa/eFAKglliqEpFlorIxJ3VgLNBciLIi81oav5+jOHue
SmrJXHYxXny5KAaJBbCRCQj3CjoYMUT75ujULpvTQGZIucX5xzT9cmUVnthwnhqt
kzRKWy4S5aA5NSoNtjjikN9QaR2E8/DjBRpHzXlIHpjT0BKgtKsXPOGTdnw/xBf/
HXRFgeAMiMCnRo359R5E5h67KaRcOENi+tiyCVXFcUmipt6CXDI98nnRfviKAMwg
i/GuYJXhVcMe6waq9+2mNZWsHBhIojUA+rzXTTHwDTctiOy5EWIG0cNHDemxLLKz
s9R3CbFRfqoa2neEh0r56hm+amgq7v8Ca2AY82Da/W2SsSviHD/1DzQBvrvgolcc
NzlESTNgp+mwzZqYebZLlWMIkoyodbwwjp5/X7DZ9WPDA1euongPYORisOTCaTi2
WXfUE2+T8zsxJylQTQuwPd+uMQYHE6ZuVv/ezk0jT+lfs1wMafVPXt4kMyaklwc2
fwsMuj9ADniRHjeSeTG5dmekidz8klGHBV49K1FS8r8lQicXtq0QJhHx6aS7lJjw
8uLvF7Gkx6tLID5jzmm7rJgbVAKW7ljuxN1okujgkRpYM17//eCRTJ/aefLYeS3r
9A8lGeK1T+WSkYiaJo1gr+FR9IWwPHxGpX2ZgC3xCnvbf2NoAJwzoYcH7U1btYR7
VGNZn16BEOskFuFsUkpcsA323jXLH8QFfzaKjqWLHIQrDPPv/PrUwNjYWpZ2sOID
18zZrNlTtyEWjw18Dow+nR8KStYpdMCy0F1hJ0NbPheE3VQi4cmi8lhQPB6UYZF4
2PUXrLVmGe23lIahaX1Laf68tdLlfnTyZ9H/7f4LKtlW6Itsfu6j+ZYwY88pVCcm
8cJ6PJC8EQIbMWsiILZeyPt208YBadw9rZKXWL32YXjOIBC+DbeCypVZSa4/R6ii
2/tWE9TpckpHE5LFTMjj4GvM8atzV2Iqvy5es1zuk8k=
`pragma protect end_protected
