`define CACHE
`define DDR
//`define AUX_MEM
`define FREQ_250
`define PICOSOC_UART