// data bus select bits
`define B_BIT (`REQ_W - (ADDR_W-Bbit+1)) //boot controller select bit
