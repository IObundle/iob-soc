// Data and address widths
`define REGFILEIF_DATA_W 32
