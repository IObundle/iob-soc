
   parameter MEM_ADDR_W_PAR_0 = 11;
   parameter MEM_ADDR_W_PAR_1 = 14;
   parameter MEM_ADDR_W_PAR_2 = 30;
//   parameter MEM_ADDR_W_PAR_1 = 28;
//   parameter MEM_ADDR_W_PAR_2 = 30;
   //parameter MEM_ADDR_W_PAR_3 = 28;