jroque@pudim-flan.3533:1589398075