// S5_QSYS.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module S5_QSYS (
		input  wire [3:0] in_port_to_the_button,                     //         button_external_connection.export
		output wire       cdcm_conduit_end_scl,                      //                   cdcm_conduit_end.scl
		inout  wire       cdcm_conduit_end_sda,                      //                                   .sda
		input  wire       clk_50,                                    //                      clk_50_clk_in.clk
		input  wire       reset_n,                                   //                clk_50_clk_in_reset.reset_n
		output wire       clk_i2c_scl_external_connection_export,    //    clk_i2c_scl_external_connection.export
		inout  wire       clk_i2c_sda_external_connection_export,    //    clk_i2c_sda_external_connection.export
		output wire       fan_external_connection_export,            //            fan_external_connection.export
		output wire [3:0] out_port_from_the_led,                     //            led_external_connection.export
		input  wire       ref_clock_10g_count_clk_in_ref_export,     //     ref_clock_10g_count_clk_in_ref.export
		input  wire       ref_clock_10g_count_clk_in_target_export,  //  ref_clock_10g_count_clk_in_target.export
		input  wire       ref_clock_sata_count_clk_in_ref_export,    //    ref_clock_sata_count_clk_in_ref.export
		input  wire       ref_clock_sata_count_clk_in_target_export, // ref_clock_sata_count_clk_in_target.export
		input  wire [3:0] sw_external_connection_export,             //             sw_external_connection.export
		input  wire       in_port_to_the_temp_int_n,                 //     temp_int_n_external_connection.export
		input  wire       in_port_to_the_temp_overt_n,               //   temp_overt_n_external_connection.export
		output wire       temp_scl_external_connection_export,       //       temp_scl_external_connection.export
		inout  wire       temp_sda_external_connection_export        //       temp_sda_external_connection.export
	);

	wire  [31:0] nios2_qsys_data_master_readdata;                           // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_waitrequest;                        // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire         nios2_qsys_data_master_debugaccess;                        // nios2_qsys:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire  [19:0] nios2_qsys_data_master_address;                            // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire   [3:0] nios2_qsys_data_master_byteenable;                         // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire         nios2_qsys_data_master_read;                               // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire         nios2_qsys_data_master_readdatavalid;                      // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire         nios2_qsys_data_master_write;                              // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire  [31:0] nios2_qsys_data_master_writedata;                          // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [31:0] nios2_qsys_instruction_master_readdata;                    // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [19:0] nios2_qsys_instruction_master_address;                     // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                        // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire         nios2_qsys_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire  [31:0] mm_interconnect_0_ref_clock_sata_count_slave_readdata;     // ref_clock_sata_count:s_readdata_out -> mm_interconnect_0:ref_clock_sata_count_Slave_readdata
	wire   [1:0] mm_interconnect_0_ref_clock_sata_count_slave_address;      // mm_interconnect_0:ref_clock_sata_count_Slave_address -> ref_clock_sata_count:s_address_in
	wire         mm_interconnect_0_ref_clock_sata_count_slave_read;         // mm_interconnect_0:ref_clock_sata_count_Slave_read -> ref_clock_sata_count:s_read_in
	wire         mm_interconnect_0_ref_clock_sata_count_slave_write;        // mm_interconnect_0:ref_clock_sata_count_Slave_write -> ref_clock_sata_count:s_write_in
	wire  [31:0] mm_interconnect_0_ref_clock_sata_count_slave_writedata;    // mm_interconnect_0:ref_clock_sata_count_Slave_writedata -> ref_clock_sata_count:s_writedata_in
	wire  [31:0] mm_interconnect_0_ref_clock_10g_count_slave_readdata;      // ref_clock_10g_count:s_readdata_out -> mm_interconnect_0:ref_clock_10g_count_Slave_readdata
	wire   [1:0] mm_interconnect_0_ref_clock_10g_count_slave_address;       // mm_interconnect_0:ref_clock_10g_count_Slave_address -> ref_clock_10g_count:s_address_in
	wire         mm_interconnect_0_ref_clock_10g_count_slave_read;          // mm_interconnect_0:ref_clock_10g_count_Slave_read -> ref_clock_10g_count:s_read_in
	wire         mm_interconnect_0_ref_clock_10g_count_slave_write;         // mm_interconnect_0:ref_clock_10g_count_Slave_write -> ref_clock_10g_count:s_write_in
	wire  [31:0] mm_interconnect_0_ref_clock_10g_count_slave_writedata;     // mm_interconnect_0:ref_clock_10g_count_Slave_writedata -> ref_clock_10g_count:s_writedata_in
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_cdcm_avalon_slave_chipselect;            // mm_interconnect_0:cdcm_avalon_slave_chipselect -> cdcm:s_cs
	wire  [15:0] mm_interconnect_0_cdcm_avalon_slave_readdata;              // cdcm:s_readdata -> mm_interconnect_0:cdcm_avalon_slave_readdata
	wire   [0:0] mm_interconnect_0_cdcm_avalon_slave_address;               // mm_interconnect_0:cdcm_avalon_slave_address -> cdcm:s_addr
	wire         mm_interconnect_0_cdcm_avalon_slave_read;                  // mm_interconnect_0:cdcm_avalon_slave_read -> cdcm:s_read
	wire         mm_interconnect_0_cdcm_avalon_slave_write;                 // mm_interconnect_0:cdcm_avalon_slave_write -> cdcm:s_write
	wire  [15:0] mm_interconnect_0_cdcm_avalon_slave_writedata;             // mm_interconnect_0:cdcm_avalon_slave_writedata -> cdcm:s_writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata;     // nios2_qsys:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest;  // nios2_qsys:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_qsys_debug_mem_slave_debugaccess -> nios2_qsys:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_address;      // mm_interconnect_0:nios2_qsys_debug_mem_slave_address -> nios2_qsys:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_read;         // mm_interconnect_0:nios2_qsys_debug_mem_slave_read -> nios2_qsys:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_qsys_debug_mem_slave_byteenable -> nios2_qsys:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_write;        // mm_interconnect_0:nios2_qsys_debug_mem_slave_write -> nios2_qsys:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_qsys_debug_mem_slave_writedata -> nios2_qsys:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_sw_s1_chipselect;                        // mm_interconnect_0:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                          // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                           // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_sw_s1_write;                             // mm_interconnect_0:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_0_sw_s1_writedata;                         // mm_interconnect_0:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_0_button_s1_chipselect;                    // mm_interconnect_0:button_s1_chipselect -> button:chipselect
	wire  [31:0] mm_interconnect_0_button_s1_readdata;                      // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire   [1:0] mm_interconnect_0_button_s1_address;                       // mm_interconnect_0:button_s1_address -> button:address
	wire         mm_interconnect_0_button_s1_write;                         // mm_interconnect_0:button_s1_write -> button:write_n
	wire  [31:0] mm_interconnect_0_button_s1_writedata;                     // mm_interconnect_0:button_s1_writedata -> button:writedata
	wire         mm_interconnect_0_temp_sda_s1_chipselect;                  // mm_interconnect_0:temp_sda_s1_chipselect -> temp_sda:chipselect
	wire  [31:0] mm_interconnect_0_temp_sda_s1_readdata;                    // temp_sda:readdata -> mm_interconnect_0:temp_sda_s1_readdata
	wire   [1:0] mm_interconnect_0_temp_sda_s1_address;                     // mm_interconnect_0:temp_sda_s1_address -> temp_sda:address
	wire         mm_interconnect_0_temp_sda_s1_write;                       // mm_interconnect_0:temp_sda_s1_write -> temp_sda:write_n
	wire  [31:0] mm_interconnect_0_temp_sda_s1_writedata;                   // mm_interconnect_0:temp_sda_s1_writedata -> temp_sda:writedata
	wire  [31:0] mm_interconnect_0_temp_int_n_s1_readdata;                  // temp_int_n:readdata -> mm_interconnect_0:temp_int_n_s1_readdata
	wire   [1:0] mm_interconnect_0_temp_int_n_s1_address;                   // mm_interconnect_0:temp_int_n_s1_address -> temp_int_n:address
	wire  [31:0] mm_interconnect_0_temp_overt_n_s1_readdata;                // temp_overt_n:readdata -> mm_interconnect_0:temp_overt_n_s1_readdata
	wire   [1:0] mm_interconnect_0_temp_overt_n_s1_address;                 // mm_interconnect_0:temp_overt_n_s1_address -> temp_overt_n:address
	wire         mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                         // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_fan_s1_chipselect;                       // mm_interconnect_0:fan_s1_chipselect -> fan:chipselect
	wire  [31:0] mm_interconnect_0_fan_s1_readdata;                         // fan:readdata -> mm_interconnect_0:fan_s1_readdata
	wire   [1:0] mm_interconnect_0_fan_s1_address;                          // mm_interconnect_0:fan_s1_address -> fan:address
	wire         mm_interconnect_0_fan_s1_write;                            // mm_interconnect_0:fan_s1_write -> fan:write_n
	wire  [31:0] mm_interconnect_0_fan_s1_writedata;                        // mm_interconnect_0:fan_s1_writedata -> fan:writedata
	wire         mm_interconnect_0_temp_scl_s1_chipselect;                  // mm_interconnect_0:temp_scl_s1_chipselect -> temp_scl:chipselect
	wire  [31:0] mm_interconnect_0_temp_scl_s1_readdata;                    // temp_scl:readdata -> mm_interconnect_0:temp_scl_s1_readdata
	wire   [1:0] mm_interconnect_0_temp_scl_s1_address;                     // mm_interconnect_0:temp_scl_s1_address -> temp_scl:address
	wire         mm_interconnect_0_temp_scl_s1_write;                       // mm_interconnect_0:temp_scl_s1_write -> temp_scl:write_n
	wire  [31:0] mm_interconnect_0_temp_scl_s1_writedata;                   // mm_interconnect_0:temp_scl_s1_writedata -> temp_scl:writedata
	wire         mm_interconnect_0_clk_i2c_sda_s1_chipselect;               // mm_interconnect_0:clk_i2c_sda_s1_chipselect -> clk_i2c_sda:chipselect
	wire  [31:0] mm_interconnect_0_clk_i2c_sda_s1_readdata;                 // clk_i2c_sda:readdata -> mm_interconnect_0:clk_i2c_sda_s1_readdata
	wire   [1:0] mm_interconnect_0_clk_i2c_sda_s1_address;                  // mm_interconnect_0:clk_i2c_sda_s1_address -> clk_i2c_sda:address
	wire         mm_interconnect_0_clk_i2c_sda_s1_write;                    // mm_interconnect_0:clk_i2c_sda_s1_write -> clk_i2c_sda:write_n
	wire  [31:0] mm_interconnect_0_clk_i2c_sda_s1_writedata;                // mm_interconnect_0:clk_i2c_sda_s1_writedata -> clk_i2c_sda:writedata
	wire         mm_interconnect_0_clk_i2c_scl_s1_chipselect;               // mm_interconnect_0:clk_i2c_scl_s1_chipselect -> clk_i2c_scl:chipselect
	wire  [31:0] mm_interconnect_0_clk_i2c_scl_s1_readdata;                 // clk_i2c_scl:readdata -> mm_interconnect_0:clk_i2c_scl_s1_readdata
	wire   [1:0] mm_interconnect_0_clk_i2c_scl_s1_address;                  // mm_interconnect_0:clk_i2c_scl_s1_address -> clk_i2c_scl:address
	wire         mm_interconnect_0_clk_i2c_scl_s1_write;                    // mm_interconnect_0:clk_i2c_scl_s1_write -> clk_i2c_scl:write_n
	wire  [31:0] mm_interconnect_0_clk_i2c_scl_s1_writedata;                // mm_interconnect_0:clk_i2c_scl_s1_writedata -> clk_i2c_scl:writedata
	wire         irq_mapper_receiver0_irq;                                  // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // button:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // sw:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_qsys_irq_irq;                                        // irq_mapper:sender_irq -> nios2_qsys:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [button:reset_n, clk_i2c_scl:reset_n, clk_i2c_sda:reset_n, fan:reset_n, irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:nios2_qsys_reset_reset_bridge_in_reset_reset, nios2_qsys:reset_n, onchip_memory2:reset, ref_clock_10g_count:s_reset_in, ref_clock_sata_count:s_reset_in, rst_translator:in_reset, sw:reset_n, temp_int_n:reset_n, temp_overt_n:reset_n, temp_scl:reset_n, temp_sda:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios2_qsys:reset_req, onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_debug_reset_request_reset;                      // nios2_qsys:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [cdcm:reset_n, mm_interconnect_0:cdcm_clock_sink_reset_reset_bridge_in_reset_reset]

	S5_QSYS_button button (
		.clk        (clk_50),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_button),                  // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                //                 irq.irq
	);

	TERASIC_EXT_PLL cdcm (
		.s_read      (mm_interconnect_0_cdcm_avalon_slave_read),       //     avalon_slave.read
		.s_readdata  (mm_interconnect_0_cdcm_avalon_slave_readdata),   //                 .readdata
		.s_write     (mm_interconnect_0_cdcm_avalon_slave_write),      //                 .write
		.s_writedata (mm_interconnect_0_cdcm_avalon_slave_writedata),  //                 .writedata
		.s_addr      (mm_interconnect_0_cdcm_avalon_slave_address),    //                 .address
		.s_cs        (mm_interconnect_0_cdcm_avalon_slave_chipselect), //                 .chipselect
		.i2c_scl     (cdcm_conduit_end_scl),                           //      conduit_end.export
		.i2c_sda     (cdcm_conduit_end_sda),                           //                 .export
		.clk         (clk_50),                                         //       clock_sink.clk
		.reset_n     (~rst_controller_001_reset_out_reset)             // clock_sink_reset.reset_n
	);

	S5_QSYS_clk_i2c_scl clk_i2c_scl (
		.clk        (clk_50),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_clk_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_clk_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_clk_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_clk_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_clk_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (clk_i2c_scl_external_connection_export)       // external_connection.export
	);

	S5_QSYS_clk_i2c_sda clk_i2c_sda (
		.clk        (clk_50),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_clk_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_clk_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_clk_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_clk_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_clk_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (clk_i2c_sda_external_connection_export)       // external_connection.export
	);

	S5_QSYS_fan fan (
		.clk        (clk_50),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_fan_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_fan_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_fan_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_fan_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_fan_s1_readdata),   //                    .readdata
		.out_port   (fan_external_connection_export)       // external_connection.export
	);

	S5_QSYS_jtag_uart jtag_uart (
		.clk            (clk_50),                                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	S5_QSYS_led led (
		.clk        (clk_50),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_led)                // external_connection.export
	);

	S5_QSYS_nios2_qsys nios2_qsys (
		.clk                                 (clk_50),                                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                          //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                       //                          .reset_req
		.d_address                           (nios2_qsys_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_qsys_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_qsys_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_qsys_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	S5_QSYS_onchip_memory2 onchip_memory2 (
		.clk        (clk_50),                                         //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	TERASIC_CLOCK_COUNT ref_clock_10g_count (
		.s_clk_in       (clk_50),                                                //           clk.clk
		.s_address_in   (mm_interconnect_0_ref_clock_10g_count_slave_address),   //         Slave.address
		.s_read_in      (mm_interconnect_0_ref_clock_10g_count_slave_read),      //              .read
		.s_readdata_out (mm_interconnect_0_ref_clock_10g_count_slave_readdata),  //              .readdata
		.s_write_in     (mm_interconnect_0_ref_clock_10g_count_slave_write),     //              .write
		.s_writedata_in (mm_interconnect_0_ref_clock_10g_count_slave_writedata), //              .writedata
		.CLK_1          (ref_clock_10g_count_clk_in_ref_export),                 //    clk_in_ref.export
		.CLK_2          (ref_clock_10g_count_clk_in_target_export),              // clk_in_target.export
		.s_reset_in     (rst_controller_reset_out_reset)                         //         reset.reset
	);

	TERASIC_CLOCK_COUNT ref_clock_sata_count (
		.s_clk_in       (clk_50),                                                 //           clk.clk
		.s_address_in   (mm_interconnect_0_ref_clock_sata_count_slave_address),   //         Slave.address
		.s_read_in      (mm_interconnect_0_ref_clock_sata_count_slave_read),      //              .read
		.s_readdata_out (mm_interconnect_0_ref_clock_sata_count_slave_readdata),  //              .readdata
		.s_write_in     (mm_interconnect_0_ref_clock_sata_count_slave_write),     //              .write
		.s_writedata_in (mm_interconnect_0_ref_clock_sata_count_slave_writedata), //              .writedata
		.CLK_1          (ref_clock_sata_count_clk_in_ref_export),                 //    clk_in_ref.export
		.CLK_2          (ref_clock_sata_count_clk_in_target_export),              // clk_in_target.export
		.s_reset_in     (rst_controller_reset_out_reset)                          //         reset.reset
	);

	S5_QSYS_sw sw (
		.clk        (clk_50),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),   //                    .readdata
		.in_port    (sw_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)            //                 irq.irq
	);

	S5_QSYS_temp_int_n temp_int_n (
		.clk      (clk_50),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_temp_int_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_temp_int_n_s1_readdata), //                    .readdata
		.in_port  (in_port_to_the_temp_int_n)                 // external_connection.export
	);

	S5_QSYS_temp_int_n temp_overt_n (
		.clk      (clk_50),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_temp_overt_n_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_temp_overt_n_s1_readdata), //                    .readdata
		.in_port  (in_port_to_the_temp_overt_n)                 // external_connection.export
	);

	S5_QSYS_clk_i2c_scl temp_scl (
		.clk        (clk_50),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_temp_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_temp_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_temp_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_temp_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_temp_scl_s1_readdata),   //                    .readdata
		.out_port   (temp_scl_external_connection_export)       // external_connection.export
	);

	S5_QSYS_clk_i2c_sda temp_sda (
		.clk        (clk_50),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_temp_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_temp_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_temp_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_temp_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_temp_sda_s1_readdata),   //                    .readdata
		.bidir_port (temp_sda_external_connection_export)       // external_connection.export
	);

	S5_QSYS_timer timer (
		.clk        (clk_50),                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	S5_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                    (clk_50),                                                    //                                  clk_50_clk.clk
		.cdcm_clock_sink_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // cdcm_clock_sink_reset_reset_bridge_in_reset.reset
		.nios2_qsys_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                            //      nios2_qsys_reset_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                    (nios2_qsys_data_master_address),                            //                      nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest                (nios2_qsys_data_master_waitrequest),                        //                                            .waitrequest
		.nios2_qsys_data_master_byteenable                 (nios2_qsys_data_master_byteenable),                         //                                            .byteenable
		.nios2_qsys_data_master_read                       (nios2_qsys_data_master_read),                               //                                            .read
		.nios2_qsys_data_master_readdata                   (nios2_qsys_data_master_readdata),                           //                                            .readdata
		.nios2_qsys_data_master_readdatavalid              (nios2_qsys_data_master_readdatavalid),                      //                                            .readdatavalid
		.nios2_qsys_data_master_write                      (nios2_qsys_data_master_write),                              //                                            .write
		.nios2_qsys_data_master_writedata                  (nios2_qsys_data_master_writedata),                          //                                            .writedata
		.nios2_qsys_data_master_debugaccess                (nios2_qsys_data_master_debugaccess),                        //                                            .debugaccess
		.nios2_qsys_instruction_master_address             (nios2_qsys_instruction_master_address),                     //               nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest         (nios2_qsys_instruction_master_waitrequest),                 //                                            .waitrequest
		.nios2_qsys_instruction_master_read                (nios2_qsys_instruction_master_read),                        //                                            .read
		.nios2_qsys_instruction_master_readdata            (nios2_qsys_instruction_master_readdata),                    //                                            .readdata
		.nios2_qsys_instruction_master_readdatavalid       (nios2_qsys_instruction_master_readdatavalid),               //                                            .readdatavalid
		.button_s1_address                                 (mm_interconnect_0_button_s1_address),                       //                                   button_s1.address
		.button_s1_write                                   (mm_interconnect_0_button_s1_write),                         //                                            .write
		.button_s1_readdata                                (mm_interconnect_0_button_s1_readdata),                      //                                            .readdata
		.button_s1_writedata                               (mm_interconnect_0_button_s1_writedata),                     //                                            .writedata
		.button_s1_chipselect                              (mm_interconnect_0_button_s1_chipselect),                    //                                            .chipselect
		.cdcm_avalon_slave_address                         (mm_interconnect_0_cdcm_avalon_slave_address),               //                           cdcm_avalon_slave.address
		.cdcm_avalon_slave_write                           (mm_interconnect_0_cdcm_avalon_slave_write),                 //                                            .write
		.cdcm_avalon_slave_read                            (mm_interconnect_0_cdcm_avalon_slave_read),                  //                                            .read
		.cdcm_avalon_slave_readdata                        (mm_interconnect_0_cdcm_avalon_slave_readdata),              //                                            .readdata
		.cdcm_avalon_slave_writedata                       (mm_interconnect_0_cdcm_avalon_slave_writedata),             //                                            .writedata
		.cdcm_avalon_slave_chipselect                      (mm_interconnect_0_cdcm_avalon_slave_chipselect),            //                                            .chipselect
		.clk_i2c_scl_s1_address                            (mm_interconnect_0_clk_i2c_scl_s1_address),                  //                              clk_i2c_scl_s1.address
		.clk_i2c_scl_s1_write                              (mm_interconnect_0_clk_i2c_scl_s1_write),                    //                                            .write
		.clk_i2c_scl_s1_readdata                           (mm_interconnect_0_clk_i2c_scl_s1_readdata),                 //                                            .readdata
		.clk_i2c_scl_s1_writedata                          (mm_interconnect_0_clk_i2c_scl_s1_writedata),                //                                            .writedata
		.clk_i2c_scl_s1_chipselect                         (mm_interconnect_0_clk_i2c_scl_s1_chipselect),               //                                            .chipselect
		.clk_i2c_sda_s1_address                            (mm_interconnect_0_clk_i2c_sda_s1_address),                  //                              clk_i2c_sda_s1.address
		.clk_i2c_sda_s1_write                              (mm_interconnect_0_clk_i2c_sda_s1_write),                    //                                            .write
		.clk_i2c_sda_s1_readdata                           (mm_interconnect_0_clk_i2c_sda_s1_readdata),                 //                                            .readdata
		.clk_i2c_sda_s1_writedata                          (mm_interconnect_0_clk_i2c_sda_s1_writedata),                //                                            .writedata
		.clk_i2c_sda_s1_chipselect                         (mm_interconnect_0_clk_i2c_sda_s1_chipselect),               //                                            .chipselect
		.fan_s1_address                                    (mm_interconnect_0_fan_s1_address),                          //                                      fan_s1.address
		.fan_s1_write                                      (mm_interconnect_0_fan_s1_write),                            //                                            .write
		.fan_s1_readdata                                   (mm_interconnect_0_fan_s1_readdata),                         //                                            .readdata
		.fan_s1_writedata                                  (mm_interconnect_0_fan_s1_writedata),                        //                                            .writedata
		.fan_s1_chipselect                                 (mm_interconnect_0_fan_s1_chipselect),                       //                                            .chipselect
		.jtag_uart_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                 jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                            .write
		.jtag_uart_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                            .read
		.jtag_uart_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                            .readdata
		.jtag_uart_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                            .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                            .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                            .chipselect
		.led_s1_address                                    (mm_interconnect_0_led_s1_address),                          //                                      led_s1.address
		.led_s1_write                                      (mm_interconnect_0_led_s1_write),                            //                                            .write
		.led_s1_readdata                                   (mm_interconnect_0_led_s1_readdata),                         //                                            .readdata
		.led_s1_writedata                                  (mm_interconnect_0_led_s1_writedata),                        //                                            .writedata
		.led_s1_chipselect                                 (mm_interconnect_0_led_s1_chipselect),                       //                                            .chipselect
		.nios2_qsys_debug_mem_slave_address                (mm_interconnect_0_nios2_qsys_debug_mem_slave_address),      //                  nios2_qsys_debug_mem_slave.address
		.nios2_qsys_debug_mem_slave_write                  (mm_interconnect_0_nios2_qsys_debug_mem_slave_write),        //                                            .write
		.nios2_qsys_debug_mem_slave_read                   (mm_interconnect_0_nios2_qsys_debug_mem_slave_read),         //                                            .read
		.nios2_qsys_debug_mem_slave_readdata               (mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata),     //                                            .readdata
		.nios2_qsys_debug_mem_slave_writedata              (mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata),    //                                            .writedata
		.nios2_qsys_debug_mem_slave_byteenable             (mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable),   //                                            .byteenable
		.nios2_qsys_debug_mem_slave_waitrequest            (mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest),  //                                            .waitrequest
		.nios2_qsys_debug_mem_slave_debugaccess            (mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess),  //                                            .debugaccess
		.onchip_memory2_s1_address                         (mm_interconnect_0_onchip_memory2_s1_address),               //                           onchip_memory2_s1.address
		.onchip_memory2_s1_write                           (mm_interconnect_0_onchip_memory2_s1_write),                 //                                            .write
		.onchip_memory2_s1_readdata                        (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                            .readdata
		.onchip_memory2_s1_writedata                       (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                            .writedata
		.onchip_memory2_s1_byteenable                      (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                            .byteenable
		.onchip_memory2_s1_chipselect                      (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                            .chipselect
		.onchip_memory2_s1_clken                           (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                            .clken
		.ref_clock_10g_count_Slave_address                 (mm_interconnect_0_ref_clock_10g_count_slave_address),       //                   ref_clock_10g_count_Slave.address
		.ref_clock_10g_count_Slave_write                   (mm_interconnect_0_ref_clock_10g_count_slave_write),         //                                            .write
		.ref_clock_10g_count_Slave_read                    (mm_interconnect_0_ref_clock_10g_count_slave_read),          //                                            .read
		.ref_clock_10g_count_Slave_readdata                (mm_interconnect_0_ref_clock_10g_count_slave_readdata),      //                                            .readdata
		.ref_clock_10g_count_Slave_writedata               (mm_interconnect_0_ref_clock_10g_count_slave_writedata),     //                                            .writedata
		.ref_clock_sata_count_Slave_address                (mm_interconnect_0_ref_clock_sata_count_slave_address),      //                  ref_clock_sata_count_Slave.address
		.ref_clock_sata_count_Slave_write                  (mm_interconnect_0_ref_clock_sata_count_slave_write),        //                                            .write
		.ref_clock_sata_count_Slave_read                   (mm_interconnect_0_ref_clock_sata_count_slave_read),         //                                            .read
		.ref_clock_sata_count_Slave_readdata               (mm_interconnect_0_ref_clock_sata_count_slave_readdata),     //                                            .readdata
		.ref_clock_sata_count_Slave_writedata              (mm_interconnect_0_ref_clock_sata_count_slave_writedata),    //                                            .writedata
		.sw_s1_address                                     (mm_interconnect_0_sw_s1_address),                           //                                       sw_s1.address
		.sw_s1_write                                       (mm_interconnect_0_sw_s1_write),                             //                                            .write
		.sw_s1_readdata                                    (mm_interconnect_0_sw_s1_readdata),                          //                                            .readdata
		.sw_s1_writedata                                   (mm_interconnect_0_sw_s1_writedata),                         //                                            .writedata
		.sw_s1_chipselect                                  (mm_interconnect_0_sw_s1_chipselect),                        //                                            .chipselect
		.temp_int_n_s1_address                             (mm_interconnect_0_temp_int_n_s1_address),                   //                               temp_int_n_s1.address
		.temp_int_n_s1_readdata                            (mm_interconnect_0_temp_int_n_s1_readdata),                  //                                            .readdata
		.temp_overt_n_s1_address                           (mm_interconnect_0_temp_overt_n_s1_address),                 //                             temp_overt_n_s1.address
		.temp_overt_n_s1_readdata                          (mm_interconnect_0_temp_overt_n_s1_readdata),                //                                            .readdata
		.temp_scl_s1_address                               (mm_interconnect_0_temp_scl_s1_address),                     //                                 temp_scl_s1.address
		.temp_scl_s1_write                                 (mm_interconnect_0_temp_scl_s1_write),                       //                                            .write
		.temp_scl_s1_readdata                              (mm_interconnect_0_temp_scl_s1_readdata),                    //                                            .readdata
		.temp_scl_s1_writedata                             (mm_interconnect_0_temp_scl_s1_writedata),                   //                                            .writedata
		.temp_scl_s1_chipselect                            (mm_interconnect_0_temp_scl_s1_chipselect),                  //                                            .chipselect
		.temp_sda_s1_address                               (mm_interconnect_0_temp_sda_s1_address),                     //                                 temp_sda_s1.address
		.temp_sda_s1_write                                 (mm_interconnect_0_temp_sda_s1_write),                       //                                            .write
		.temp_sda_s1_readdata                              (mm_interconnect_0_temp_sda_s1_readdata),                    //                                            .readdata
		.temp_sda_s1_writedata                             (mm_interconnect_0_temp_sda_s1_writedata),                   //                                            .writedata
		.temp_sda_s1_chipselect                            (mm_interconnect_0_temp_sda_s1_chipselect),                  //                                            .chipselect
		.timer_s1_address                                  (mm_interconnect_0_timer_s1_address),                        //                                    timer_s1.address
		.timer_s1_write                                    (mm_interconnect_0_timer_s1_write),                          //                                            .write
		.timer_s1_readdata                                 (mm_interconnect_0_timer_s1_readdata),                       //                                            .readdata
		.timer_s1_writedata                                (mm_interconnect_0_timer_s1_writedata),                      //                                            .writedata
		.timer_s1_chipselect                               (mm_interconnect_0_timer_s1_chipselect)                      //                                            .chipselect
	);

	S5_QSYS_irq_mapper irq_mapper (
		.clk           (clk_50),                         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_qsys_irq_irq)              //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_50),                               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
