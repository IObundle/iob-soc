// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZuqpfXossQOiZDc3aK6OfoCguz65spWO1n2ukgenq/3HAHdCtPiRpeIeDrW0zIQV
MPjSFZI87EIaOI89fnLapTXNRpbgugiHhhAdN0GWWYVHRxoSgsPmKi1LShgKfvFO
i4EGuw1uwFej5UjLaEcS/ka98MUkqVIrHmLsa7ahH7o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 51200)
eQp3rujyAynplaOvLcSJOGlCfBVBBHkY+HzgBx4EZSUo57AWDA1XhA9Tf80uvrM/
Grl+Pez6B0+C9f6Ax4j+WE92XIo+Z7gdv75dz2SLY4nSG5dJrH3Z/mncJiryITAG
4Gl0IBiGZprsCiVVOyStSvlEyZl62Ofw/06WZcjp6mgRgViihTTqdkQEYSHYjx1P
lev1I8qxpZxi3PNOmQeP0H4rjlNCt0/by8gYNV/DHme5kFqlNBmn0R03mO31zB2W
TYLm+8IpsoRV167TKIBYXPTG6PzcqlNjpBljdieP3skflu0tc6o8N/Lnb4N9jRhF
ChvJozR5tgYWfoBxMC0qITKcfGkLHkgV7ssT6LzzOBWccPMnVnFpFYy0PFkihLFZ
RHgXv5gA8dev5sVoRPz8fNSUDv/g+HM78lA9PAb69CW75QHU/B7nC8pkq14sjlqR
QilYsG0dUpwDuCOYEICxyJIrDzX6mF4FUbCOaN3aKUwc9S+A+f0QnrsCDjqwyFpk
3prfFgDlcNd17DigWdM5d5kMtRDS36N87TCuJSKKDIsV7t6e2CFeXOJkU9OBW9rJ
fY1PBm2qdMz5ihpJ5tjOU+0YhjGzT4vVCLKk54IlRr6mScYAecECTaX30d68zzRj
7ZGtiU2/Hwyj+FqsGs2Wb4xlhEZmGCbbL+BGJGfVL6GshI2Z5BzdDyXYKxP6H2Ku
Mw8/RohjNqGsrWfV8jbCiO5YvuNeev9XDGZjud3fxcXr5CBV/7BslstWXmRbYM6v
mYWqGUC2FbDK2R3PujLM5aVHW/Wg4Y4HupjgD9T2sjWM6PfCoOSelIuD9xwVzg/3
EZSYy9mQurjDGHQ2M8V+9DvQyWSvnBmJcco7hdzx4MIBwUnowKsU7erTZJJFjhnR
nZ1RneyMLJ+NgglDHZ14I+rTxK/oqpmH+Rfqn2KzlXvJbZZkAKzenhULvdXtyB2T
gHex8Llp+gLim+PJOJAQA9RxUQ2ngtSEO4RTEasg/Dp2luZPBxDkzSCKMKoemvre
fJtA9NFJNx3YZoZx7hpwMcCPGoLcx8ijgAjMQdQdl3d8q/Xtr36GbebESGd5nZbd
0DRlkFyNPULJFlgSs78LEHIbFCFg4eWQCwooiQJ+Srnhdvs5A6O83adD6BD7dxWo
uFo1uaZvOC7yXvL1UZt/R8Z6tE57BriUGRKIk7movZzVxcwWuGI+MkWH7E5BDEIv
bVDOnadgfS/IE7BXvQg9AXqwUMeUFe/WinZSmpm9MZv4T71t25kOM6Cn6TvutO7S
pOk6QoLh8Eem9SsZxMyqtf0Us7EJgHOHBrfa/IWPHYw/a0Br3blKkye4S+dN/OH2
ttjtsRxJljeOfMYDpGboNIcKyyMzHNhyYUMjbAeJmdxREfyLSvlTEKJcRLGOGe5B
JoIwpMy1nm4imR0+VAHr0S9HkhjhpIJwbOhdYuEtp27Mhc/FImKhvkWVSbXr4yao
Fi/i6nnT5ewsSVh3Qkcq8IS+yi1U30K5ctcfAv2O3dDuEBtVzBtDjX5EfwihUWl5
vQQ7sRxDApL1jJ5Cnr9lAvLe2SgEUwN8h+CfWzHtjY7Yu1Ya7N3OwcM6lVTh0G30
f3JtjuTZoUyzlpBOzI2tYjrkXjbMHRcAR5Q8Z5OgGzW+CvfmsCgAnfEb5VK4Wflj
+KPR8+luYhpk6hDHcS5MaK/5zc6ipfxxqKVR2wKXkZ6kaV9ocZDJ/VyFDprqQqKV
8jaIz5Mk7NvRTZ/47eTnqdrNQ8PbbxsinjJUYC7Cw0c+Ox/zNHQ5Cpe6wwGdZgNG
giwtkzROBmx+pRyGAwNXcHaMkE4APbZILD0qSHbCkQnkNWOWIGAzfakA9X28yNSu
FyIoLsDNiVqNk86t7KiuApJOg/oM37AKK9MP+usk6mE2Jx682pmuNF7hPw0fagBG
COCWpPvUr4XCgmo1aOv6tpAv3rs8tZsTs4OFjJAI45XtVkg3Q7b+dJIFGwhBLU8q
FE5zK9zfSsQTLezUdkXWQolKU8MiuVH7mZt+AMxH7hw2p8HDWeuOYLX83J0DSHgG
hIXycXJ6z/UUYhs0S58liJo6OfbFcS84fmrOkVbL3JRZS1tdv3z4Rrfv+SKfkfyn
2q9qqAtqPqpQQoBRiWAFDz+GbHH/Fr7ezzCb0/wOv+GTeZcVYHKDmV7IDvsfrRWn
tqq2yVu0zaNiyhguKoWpzm/lwjZqrj268UbTvDgtvhA+jBYwkCXwwlZZ8IhncAZ7
SjQn/5EvLUaIMql/265GH37MnIuKjB91zaiLRC1EdXfoVCCjsbtW09sZcnVq/+Bp
PTtQcZHu2m3JSY7FE+KDlzr9pyIf0SH2lidITHk24+vyxzlSzSw4l2CPBbC5fT1E
PBgGfpBBattVN5WyB+/Kg6cyOt/DThLRL1gWdxZEb168TZJpRBMkAeEd2ndD1zTH
lr0teD1wOl+ZIhUIMdEbwTq6NzXHjGrF3n3OEIu1hH8u6G7N4nar9gOJ9vyOWiNB
jLYt1o486Nxyt5FK9AP1qDHaRteF8udaaP+gArxNPin9whyjsDGNaWmrCs54LgYj
iqPZzAoiik25MIOpHVb1CRdN26U8nTTGPDCEXB4xVdE0lTozW10Cm2hLcz8yE3cK
BqM+aBy+y6QVqm54zCYV5atCoJ1NX5HCw5KM6+bYo/hHsdNM55bhQ6M/IZ5Z5lIC
pbEP7PeoOhBZy3yTc1fCDUNW/eYXFl8In8mMYn0aZTCA5ntHsbpRo8p5uPBZeqJr
Hqplg6TB2pPTRhzWO+HXsFL4iuSbVg2HbLuwrt9H4etSNoT33L5rkDFLnHkS/Nje
WkC2iay3Lyedt471n6D26gUxl8bs7p8tYSyghVSCujjc0BW+q31zObGz9YZ9BABx
NHkmMPAdra+0/VWZ7qEfrKir5GV24o6nX+dYrZmCio6kRkCfNXkj8NOU1UhSPg2M
G4fcqx1MPz06rQD6BSeZ8AxTql9fT/p/Cfxya5s0A3d8+XcZjV2KLDaiQ9tZJFYM
rQtyE+1suf/Q0XYJCm6TqXElwsRbkgO7JkUYfsEFePgmXfK7w04WrROPeIrlNvqS
YYpRRHF5K3MSH7wlXnXCOTdG6pIBZckTdFRWRfC3HmIixwd/zW8Z0ypU8l06FsZQ
sluL2og7Z6cENsXBEVNJW0oTndgcovCSVXjD7qqSEgo2e/lGInaWwdCgp0p163AV
rLHa05D+QWq2j/P4szPqUWRyV3POeiHtMj2KLopnwmvwMEK1ctMS1RO3p5zJQw2h
s5h8b2KmxUwHN1DEIY98uwP+pg7nnqDRpPfZfadhUJZ+mi+AuxzjkstOQqNxzbkr
sdSex+zU+XVBrADK8DN6NMVfI4ZXJwc8N0KxoAXEFvIexedJZ6c+WhWtilUl8toD
5FSJpYgzvaLttfrFAx1WTR/HB8+eY3+R86LwFI6Rg1MzeAAv/OvqSBR29EjxTslx
q84RrDaWO0FPogPB8f5xOa1ePljbz6uBfUoDYH3Q1cFtaNcN0OjldzwLuxe2BZDu
Rb69e6xl6lScLwIR7hrxjG4oNlKB3lLmuo7jJwKktWNM3tJ0DuoxEe7wYuJBhUdn
hXcHQBYitqFB36IfkXuX4ZMWmgCNBzLKozjM60ov9gzNzysjIBeTsmXKPORQpZGG
/Ttmh40jJ9Q1QzzluX7JefGdCTbTvewwTvZ0ZbPmOX4BcpnQOcyGjoMCsjHIQ340
PF5B9ZcpUS8gi+fqpJ+kaS/ooBZYStdFF7cOL6vSwx+U+azPGRl2p0NPkZlLFmdE
DEqo2yLJV5Lg9j1KVBYQ6rFA3VOxlfdSVFufNoyja1MsiB/8uKeXsjqnCPzv2uAi
k4+ERxts8AfPaOBG9T2oqyjxWjouUU0rGL1ZCiE5kqE6JwCSE0YWL7lP3CYCjn2O
KeGJplHV900e40I42r4jzzVBHHH+HrtfVChhdeslGLGp3o0XnTfoTJsmzlBzkC94
yaRuZRw5QbG/1Y1FJRqpQ3Mole//IykSYT10rVJjcQGL3QAZeSclzfwotjwUY7KW
xYMWD38qv3W/6Qhkd4McTJiqJI3C1xbq/yciFsgvfaE2nmRJmx3M9LGvaHh9A7rt
jA3WuIs23sqMtJbgTdKAX9hLiz/7b9zTrhdLj8gm8jMcZkl93txf0WTyXrelN4ch
Cs5yK2TmNHjczxqjKlUEBNVToAjWEyqZC9vkXiMacyLpUPMhX1/PUNk0W6DuPZPn
nhfKd6OYlm4C3nBQxUJ8+9/5bx3jDtl6I1fyiBLIZFSJ8XdSo8vOkVVS0pWF/x2Y
JeM12hMOwraoq1bDv5otBkVSDUGRoCGFp4RUuoQbkAXsxMxv5o34EgTRw71q7aZ7
AbqXPfBz62wjaTznTM3zSRLpEHzdDaHGp3innP8O5en616pXH9KwJDKtC2LeJaFa
CznPJZ0BeuEA30QiuAuAAuTC6Yu6k9m2TqTfN0xoaRZmOJNskEnw08eAmF16GPy9
QoRSzzZs49VeUiII9/E6u8P3wuZSpYo5cu2WX2Ku8x3h53gV/oZR2nIbGA2/zQUU
wAAULqDmSSXSiSNOJ5JUeSHm9OovS/wKhzDaglpugo9sqcAELUwDetjilKxnU/E/
Ty9/F16BGqFMrdbryuY8MYkqWWaA0xtimDjt+OM7Ym+zb9Bi4aEXguSDsXnRcr9L
wuU2IiF4rlNGG+pcYGNzqWQZya4ahzSkDb1Tem7pThCI55eOVuQjJwOCgxvvctea
WqZHchV2HOd057xPP7Odv/VRZXv+dkkhv32oBnJDjPKu43LXPd42FJRKa4spuuSe
WRiWvMUaxSkEBwIbaB8nqqaxO07UgeaLHT808p6dOeDzTBEoLecJ6JRVfZePzC+5
iLaYGTjPEhD6HLsGiecfy9lZPZBjEap9Kr18QaQQWDhbGYSTlg4oAifSSZCEC0tf
b/EKpDZ0AJRNTGD4a/z+EVfPuOEepIKnLo8NyBHq2QD5urihAjiBsUBXw7X74NIX
snuw7gpcDMAPtc6Fme7r7WU/jHfqeqWMsabENZnrekOUYR+Jfr4kEdSGjtSaBD98
Rrsv2ckTcPimVJHx/svlqGuYxahlMMC4wtW4kNwpev13VTtRpbkaxRx0ahQ+Vv2e
a2xUYDSTHPegxc7u/rpwNkrU/chh9bw8uwhfzA8zINSn2jWm0DdihYstvO1xvuwx
2m2rnYh/fVi/DtUNzpFFEVILR6GWRQaWivY4H1EeMCRq7yo7SvxkrO9gVNHdzwop
GERFyZcwNnr0B0M3d+vy7NzZhI7v3dpjImvowqbwlXNcGzVLcV8g4sOFB1WiUk6E
y61EYXUxuc1syLMT9QLmrWVaKYr5+8Fp27tHO6+hsc0s8fY8+lyjwTnjDQRXDh7Z
CHVslcjMEUfENba016vOGxjj/vX21IeV0Xty5RDXQn2xcmKsrrEXjJC8oZ5zUMtJ
lXLLkrXdnAtOJkT3AYLRlebc1f76VGvVLEN52gT9fVfYTtbYhsTekgFdcxkp+DdI
4Rr4GDuvSmsX2wITuCFtGCtQw00B1NSTkOz33Lq99yscdUvjjTv+kES5d4aa8nin
W4Zd1Pl9lbwk/5/gr5sgH7IX3sAOe0tpCDEraybHhDwNK36vGBZTb9XzblL9JZWV
g0vV76ljuBfUEv0uEMp+FFE6wZmoJLpmmYlqQ09jmpoimmY0EHhddl4YsPmKGlrg
QNM0P71l053ptw7lkFwS7dymDDyBtv+LOrjAC0JrPVkgsSNeWahvClu6MuOp23lX
mXl8St+Y+ZLHZ/QsmFzMSMR9WJj3tStjj3jvyRcWMW0yUUhPCz6JR1Eanub/W/l3
VxWAbZJsZ54GzeKEXjff4qXUE6IvYs7lUIhN8YIztjGyzUbwV1r5qUyYy+wmKOrN
9N+lmKRKLz2cz62C23Xh524J1jMamC+D31rA9+kq7NpznKAIaxz1YT6raXZeJUUS
nGju/wLkT1cNUqKeH9lxzOnVZ4sBlPEjuTSLyROg3Aw/oj+Z3YFloCOnFJmmW9Ba
Ng7BDVIn/kPi6B63MT4OCyZOp7NeI1nzsGpuw4vx6jr5fa8yOSu+kOqlH2RWRp8a
SIV70iz9zRCYeCtUNHL9HzpklDQg6ItNf+KBmza8rY6T53TELoe3AEAFq3d3WMsk
gQgIAtwyjovi1/oTeg3kOVCigXOhPOLLfcKIr9XKxzRBlXMroBnHgIMXLVSI14wx
J2apaA0CtFeANpBHJF0+OSsnTeHrVBij6U+kKAswaxT5ff6K9yc3hoZIYfOywmLY
kxWHnoE7meVwZvh3KwfneIn5g4qSQCKkD5jEQLvi3QjVQUiPGQth86gWFm4ct2Np
VWIA1qMgmO+I6pXnE/nL9zUgdGE85chnlNDKyv3d3kdqv5u4R7pFF9Q+BwNvTbjl
XBEKdZClnkD7K3rlEd5DM6VamuV+taq5KSLv+20/229j+Bi5vkfZik3tW+11pWBa
rzKrUdTypTlX+s5t7OBKGGV+kNQEg1ryDskaz9kJLzmgGZXo3BWofAmH9mCF7TU0
JG4aTL+JjrxKo9x1o7fB30GcMc4dbaZEO8Yylow/xJbZ/Y0rkmC2PiM1JK1qEeBN
VYX2O3fOCWwzi8CP4hRaihvtf9ihTKUBP8OYKA+QSBpLxYLacHDCxMr5AmZHop0/
sfBpTzP2oNytmXRm5MzRGlV+zoYx90uCzfyDDn2Hsxb/jK4eEk5DnV3QZZzuj1Mn
1QzZtuRRJdGFgTNJjDvMeN9J6kMfGc7LgQz6GQin4yet4dAU6AOJpj6RssZzAsEA
9eXhT1r/aV2yOLj1vAovERQpwCMksnoHtq83iOE43NKEudAYeqTxBq4M1+j+/Qtj
SyAJmvwMx6ZrHAx7/0TvZb5USdSSHvQvwwXfRsTuAuRBh/jsHewyWWNI1rwCi806
wyGmvzg+h/PnewsYnjV9y/B419sFJXuUnSJ5uVpo4SQhWGbNp4nfy3/3C7k12914
T3YQPgS408DfLI0qWVsiZMYAns61TGWrn0m48A2LLDW8GxgZBK4/DDXpRjBew8wP
oyRAtc66MRNV5Dviue8voC2yImNreqRh0b15s5/VrDMEhdniLjD84/eCoG4+fl6s
D/IizEj3WU7M43oTsQgPnJG5ad7hDwNUZoRCEQRk1aq8uHFLbf179kooctJchtwK
+hAqVllaoFOVyeQx/dQlPf/W/QHKIcJ7gtdS8JCEJ7AZoPNJkK03cY3HeDj/HnPB
L+/0shbTLXXIxCXI4QvKnjg1hFPpqZWtWME7vnUi48042moycHBmNLH0owMHlEAK
ivhllUtVJe9vjWVoeYlck1d6z/uR59ybqwtJcEkphNWlGSmT6CLVWeceh84HeFys
SngRMORg1CwZ3Bf0Y+ze2UDdhDyFg3c78NTASu5D2TkPGs9EjrAOncrwDywtv+dS
rT/Ib34oOcaK6zs6RU54Qd0zid5sggh+riEZC/ycEC2XPDHmooFNRBUhC6iCFKxq
lWmTsv5XUwGTAow6I9sMUwCOBJjqHmDxqJ9gg4Z0r6NFww+kG/XUj3udk0dzH04o
RX8/89VAPDUrdpMchK/eKn09Awbkme7U4xXH3FnvYv+IhzhcxDtW6/ReA/ihRFGM
D1nZcy1p+qpZU7sz8H39mkk0PablpFsPP92sc8Xw/hK+W9jEbfP63oJEy9120DTV
wUEBb34oCSnTNrq9PLwcM8iQYJUpfxUer0idalM7b5F16BWDiuYamK9W4Qo3H3kz
KE9oCncpket58N3qf4JQEEs+Yp7pQgxZfEPSn6tJizyaFAAtkqpTAYCLzNJc8muQ
wkxTWpQiiZz+qCpq/Vd/pAfCSo5l1ACU/rgK3zWlQ3n/2a/iQyoPwpxaRfUq36u/
3aZT6AfY6lqYL9PkwU4V5/1ldmVxdm5T2UBR2WdCCfOAGWn/yJLMdsVp0IoRIu2a
IPRMBPxcmsmC8OwmYe4ntNxU1k3HndokWsqhFrEZWazwp4ch4oSiu8HgAf6bhbqW
/U4B63QzkbadW+bFKsJyXlp+UO1sd9fR+IgsUUvsnPtm1QUdj55BXg3UEzkxk09j
Lrj8TuU2sKXeEQ01tEXLlZHfyThpxNVTPBN8wrwz+usqyc925u7ynh0E95Fw2EH0
u5azhdxt/7ZvYIxX1BjEt6arbT870YAgrguiDRtb/JkTz0q3lq52h82ai9kjGoQ1
VGvl/UuGMBp15dNepFW4anqxZVFDSqDVVXjIJcdkRfF5xexQCR4hVw4rbqwBNDvY
XPLBhTj79PsB0RcyToHLRNMgxhnJYLFxgxiYpn+QzM4jPySDKQTGZaMPGGSm0DIA
PjWpsX1LIaDpzwZzmtm1SAhXnQYdLzwJAk/+ZYkspZ8HUhEcO4/REsjnFS+Vy31j
Z8HPrfDC+BY6p5nWXmPLdwaN0qpRdT18Vry9noSHn3JxMZvoPl/LwjFMOXRajrVa
EGtJBsoF+/Fs6W1/XwIexXqPyloDLxHyEiWZmyJ7i4fzJ5nXAghpr4YiieddYw/m
bX65pLjFi03muW/4HuLNbPU7hAfjLRCpwLfs6xWZemb+6RCCJj7GtY4L0eYBLJ3E
ikINg9f8Ad8VgedXTB+N+HtG/VE5h/sPCdvKSaI66wNClIE9dt4FKHFz7FbI2gQS
mER67/Y6m3RcV/4Onuk8WGxX23fsJhYSsLbWfL7TAS5I9wOM4EGbFKGz3ydN0eo/
Ory8sL19eAr23yq9JPMzWDkqrMqmGIXop/LhhFp/xRlsSVBgcmNxG1l1pNectwrn
vrFTrW5e42Ze28Jxxu8nMzvBntfJ+yz8Ux4B1wC08qrXLCT64qcYiKLwuaeuN3oL
vAz5tume7sQEfnhCn58371SeS+MJm6Qf2F5qusVaUxjuOyABnQYbRE7y9+vuddKI
fhfDpW8tH5OiLeRpvLrmWFdApBbqdZKuRfJExo4im9kaIezWbhAzzNuge0wbGHOP
obL8NGFJcQhKkJ+ThH8FEuSQAPoeTlOaPpHEgNnc3a/9bMhUgsb7+5ITG3ZVHdmj
N6tNPBTDoKsowxYseMeCp61UbPl4Qcp9o10P0VJRjBc9y7AZx9pZIy2s8P4GY6hr
+Pz3Yz8UN7SOXm8IRTe7VzMj7iyPFkkeHw2Nagx6UbRzbrEBuAek5UVwnGZ8Ok/1
nUl5Ih9kWJVVikgDQ+ptXUOBO9kqh4ujUP0KFp5FavXAfxnU5bC56+kpVJDungLr
zIv56YVeeyM+RIQnmjTLjR+7pW9HrpmXD14/rQ4mYSjcgumNoCOEYpbO3uT4eX9W
3dBlhioZQNTNLWl4p/9g0jeqLZBAm+xlJme3eoTrl8uvKTIEYnMxhSn41rz8y4qH
VVCyAYITXbJ8jziZvXN+QajwOU8MxQhF3dEOMb91w3wus4046Rs6nDaDe8pr7S3v
c0/0nlyWYdVpTLNyK0TqVc7QEWUcVbduD0KZb0s4jxn/xCw5sLmo6/F3dd/LtZbf
pTwfVLgEpMEmu9HZs6yZNQnw0Urztf2N9VUL5dNr73G9xO2iobYyWvl7s2DESqT/
QVSFIWh4AOiCNGybGIVTCBXkjgxoAsBsN5ozcC5vwEYzgMRs01Rofvl9yx7fWYsW
PHe/ejgmzCNaCOBR0xHHuzjsGyqLl5RZj0yVI7jQCHhBxe8H6NJKeXXUEdY4mcaR
Pk31m4vSFKAK88uG5yYih3amBQg9StLSrHH2KQ2HxdfVzc77s7wNtCp6lnT8uW3T
VMECGN1qBgQbeI5Qw9G11DWoYSIAi3kWkWgfRDpCXowJw0XDkWhwIMwijUEOkmHu
3ycZOCDYSmRRsyOwj0nESsRXlch8OwYIODdK31nGQVj/E9sFN5Lz5/oZtLUbtM2B
VQh5HmCzz9CyxWOCw7WjAGu4kW91KhjpRQpbYpn0RF/dXIg7IdzYkd8o8hPJE5KF
maAYcfTFwHbbxjZyfg/KYGEMgMvs++fxLYNADtCNP4ZyynJlMS0FFLVJDznqoWRF
3SyZG/of7vf5sph42Vg03vcQqTrxc0XEZoFnX7l/R4LeJqsAtGe2l2oNBOmkgNqo
onp8W4dmpPrf2z4iCKqrCpneA3caxPoQuskrJrUymHGf+5gmuQHeLcfRzXPtjac6
y1bzlWrGzuEX9F5/61ZD5LnxE7Zl5k7zdCkSUrUkI0ht+W7NKJfybIjIVcEhmDi9
2Rzv8MgW/7l7n4ZV49RcX4bdecmZlUrUuIPrGLEgF+aQktPS6cQ2vQbqNy/qrN2k
pGkV7wkdZMtRTDVt6TPyoWquWPPUDDnwO7awhmLlLJvbxa1J7GPieQERNOBT9isD
vGd78lFgmtfLvVyk3rrgZOhtCiSMC2cQoEdRr2UKBQVTqNVBr9NH4vkg2rXvd1hd
wKw1ZtL3IC/3Np45OWsNjCHzerQFzSrkEPn1U0rlYlVAArgazQPMngyKzR8W3PmQ
UVnK85vgs1IoUl1U1g7lVQCEa+Fej60//D/nsIFhcaov0a/T03kzDS/U9bltIzeJ
1f53/jcsFW9eT62mkNW4jZ7Iojg8evY4eMZyMD4N+HCn+DPNQ9eoxY60DR3yr9z7
9u25OoTsFl5pOxqrqKSiqCFX01uVv//CuvOG45x+Tdxoo6kx/otkXK9DBZ1F6tl6
jx05i3fTPO4Qj2G57QarfPgWM5dmWcfBukVt/mfzdKsUzzb6u+oTJrEmypW+PG/l
5MLLy6NFRE1tzX3fosK5UURdcNQIwme8QLcQDMpkDCAqoh3TVVT6bHvFbg0iRfMi
dgQBx5Jgm5DLvIdlWxFk9cEN2L4FlLbjBLtJ2jXF4hJTbdQ+wcU9IcERRbhEdeWT
4++Rk13PcUPcg+z2GdCSVS9212lwqSN3qcoVwOV578nndSCn5VhSUeZ8sw1mh1U/
pTKQqKLDSyjKMOK0gWXGwNG8eYNvQz15yIC0WUwN+mTDJ1tS4S5hm+u3bRnVbYfh
xC5kindmJHRJ/8rRn/ZjjvBDMxwHnyzOWBjAbMakKRMFYGLPvy6fHP/Sxxsnt8bp
hBtgkwcUZpBWtPPhkdFKNR0Y7OOVZvWsZG5uz/x1+WEznj8JMRIwe/REN0LMHSx2
wZiIdcF8OQXVspuAE5eUtLdqrxUIjDR/+C3PNS9NITuyxPI1tSUVAMkOA3EaOBXB
+75OrkYY94CyaqJVjxVpZ8Da3QM/TX4JVpo9XCDQXE+Fo5ckyF8dm6BAHsQNNdcB
mFFUxrSJWA04me4N523jlv3oZpbTC4pdYAXrE3bD5MN/xxv1MkuKDEU/+nfNkbL/
F714sRPJK2NvgJ1m2CvrUkDnze2g2maDK4tgatz/EI28UKi1nKGOA7kzsaOPnYuJ
4nc5y4bTDtfA/U7XBivNT0grqZnjpXPGpDHg/j3t71NPOoPfwN4kSJtNJ8pJ+TC8
NudIP/y9PEH8A2SxNrvu4v5zw+IhUZydL68CYvQOaqbdrYUQTTcriIT3eDlluwDW
tUY7jBME4x0pYafioM+VwzfbQ9kqonzoXdUdG1dVTifTaEuA4cjQWlDLPndppR1x
qMygIk6a5cCt41dSVZ/QZECRQDLLfOzZawZw19uzqoa34oyl5eQkkLmKSKwaQy7t
vs3zDfoQJRCXHI4BmXnoztuw7mLAEVOJEKvti+rdITo6UuES8dJfZcnLumvUwiZb
1N2wk3qa0y1IT5IrGMbIglTECC+EamUsGEMej341NoZY2oV4hqLAttF1m9HAYd32
fJhHRyqHGTIpXfw2vaKZr+XGk3eX8+fvLJzJ7zk6SNyd32O93Mrsyu4inhRuA5xd
/y1XVUEN83DK9AqWfDR85ud2i7w8GW0m78ZPzzrBXBSd/XhjkzS7G1PmJFisjntN
Unl2H5fLVkpp2L8boU7Pfwy09wrS5HgGvSFqbDMRsF3FCvQXyz3c3mDpeUWAj52h
roc/zxApFF9tOm/bM5po3rfh5Hy0Pez3xOjUuSSz2doEf0q+jsroOVhL1bJu0gKi
JxMBYJEj7OadbQXcs3iIea0eiYMP9iDZifM19NVF8Wc3rjTYX4EmnJDm9oxwxWTS
T88IIk/SxrRb/ebXLazoLWM0liIPGnjSigd8/7pIgSCalkEjZflBgryGtjBp/lpz
tTY5u5jVauwk3CwgFBsGMSr4b/jhOzG8XwUfJSWeVBDvZd/zDREfHSYzydxvS8Nh
TE+LFWlDD3QOH0g7OlZ67lxar66S+j0Z2nyMXj22LPzxd/sg7G0mbsNcdLPjlMFV
VBp1Tsnhu1QZJSCwYhWEf2UtH90iZHJwe0icXMv+2lioHgLt9g1DXo6+a2vqPpWm
Njunhkz5sqH/X09UrK5U4ciRjUmSaZHNjUrqLe3u7fQn05rDLxAkyoPUK3kX5YiK
53ZPbVR/DtizgWtRqS7D2PXd2aijVHmEqsrw1miXxgVkI5dT3l2AdTbf5bznnqPs
0V5ENZCLigcAygsFXw4PuNhAnpCKOmKS+v+JlbxklR0R0o11XyYF2xfiyEjlbHWc
+AxIF7eIoCFybADFdVv6jHou6OEm56yK3MU/BnHpkOnRpf5rk+0gc14c0APwrHgb
2MeOh/umx/Hk+bdY/9vEwnNU1woCpn7fXBLqi+1ZxhhjnHjB1sVNslzpIXV6nCYn
OoockB4mLlCO2Xof82NK8yYtXlM/tZnHZyi/2IpG3sVIKaIVBhmHiRYd1NdxRj+L
on99Q7ZqKWZuQfXoqbkDm/kAp55F6WBmU48vGx5EeVj/ecYDXKsyc2jUYTbit0Y0
QmovXn+OiuePlIE9oPFYMIxC0tkWgRYsyRMJuMU3nGGgK6ymAtk6fdSalF4nbiE3
nWAPuJ9PqFvm7+Xl6vG0hARoahUeeSHsv1F4jpeUShZYxi7xta85/wGPIZJFfqSE
/JLDx104PitpnooDfsivmaLwASsBoS5AuPGZC4rXR0Xg9l4bfheCp1uwDwKpVzwv
CIRsCLKAzACnSvi5Ntk1gMLUqnatrQ8WqtKJ9eXtnA7SnDxZIRkG7Y5NznNqqjHH
O2gwN5zmhj4+ij5cGpDDLljEanE23Xz+wouSc/odBhsWolZg3vKQT0j0xVD9xd4k
dSUsP2EfOdltTyVLSrFiuEipurFpxLJ0WQGABuX/4ZzqsgHj4B0cbvSEpLv1VH8E
vJR89RD1hR9Ds4UGrvKuW8fAmJ/BITdFhi+t6+M/YU2/+vomWmxuA58aCadIdf2w
RukkraJR/GJxZBgtDDCzA+42NdsYfuXx5qGfBpwb4NBlD3zycMmW/6V0NV1nSAkw
O8ZYCaLfzFhGnIKNfRSX0/Fm+dac3YipRUw11aLO9h1e79CsPAsSWj1EWILqtgFN
HtcQO3MUhMiVEr0nloOTAJsZlhEKjT+0WJaQNQVLQXlmsrZn9fcbqJPMwcZO7mWj
Gx9fuFUJJhEcUdWxYiXm69zQHPc4hkX4WdgFALkOesHgEj8usdko2twjbYk2zq2O
6QwZ+k0ZIO5UmJZ0Tv3m8Z/nfDD3+UuXn4LKOR5CNfyy7Tl7vAc+15t8Kfc6Iy/s
3H4tVlegAw0Ir4lTHuHFEfrtTINEizSrZagv9qMKwRhSlTuJqmqZ3jBr8+FVkNyB
q05fScBW1pBvHTM5fVd4Rm1MPjg7mgWzU/JCRU9C25W7ARsMaP73IGks92WiCmhg
4noujmAnKty3wVTqPDXGdwFcPsl3APFEFWQkt7J3t+v+oXuIGF4l3i8FbssU/03z
/y1NEX08B5kM3a3zLISX5oqZ1T2/w/Yc1T8Zy2wOQqwutCaBDva51rLD+Bk96CLn
7A807SZu7VFYjzlElqqxXfxWOPBMYYmE3WNKFCHO005yReBpBccazXZ+xkYCR4hO
ZWd6bls6RMyTv8GW2ZhBwcX6qGsFd2yKYnHPuag4v+yiqqDAirEMOjUO9kn0R7Og
j7HofTQUapXv+xbRN7sohOpzJsYmZhsS4fB1N5MiIlcn0lebOiCZ86z0uJ+TYp0h
L1HMlQaQqWx9qzoXkvLuD38LE9DRLpP+f+1+0Io6OH0vmDYHrK372y1x31wFhJA7
X6s0L8bbn8aC1QsC+APz4IhwwqBm3NpTH6RDBvaABb8A+vi3V/ytOdaQPHhr7ZWb
rQGxK/Q8LcVT+hav1/c/hrebYW47OS+68rCqhGbq6ClfDyBdBYOZZicHdEP5J3TP
sZEDoREMFqd1rgRCFUSBeiB4BC/mCrlXVBzj+lUtHyDz7Y8s5pVPM2oz3CfQoAbK
ucw65ojj3EHa00RVcP18ZIy2zIikTjR1n2PHXnOfukL2zZIwBFHpZziTjaXVSfwI
rpqRVV2+H8PF62o85XHT7r+ooqIDOq4Q7GBk61IgMwptKeg5Mp/eJJ8WCoBNPLgM
GohGJQDfFnv/JUC6UgKvTbxBHBCa7skJ4EsWClRehij0Gd+ljZRRCCaUTUa61zQx
INm8lu8zbBGbn/gcn7selM43UXZyEeareiorrl/uyqrPFWfCQt6qOK0iJaDXg5Al
RkPD/DGMGNXQS4NK3AmZyc082N19Sck9tfu8VHWPVNJfbItiD+AaZvsLWis8SkhE
F0wqOYzRZfLiGzrl7ScduEUcXDPP2Nh3J0Mhn/iQ+ICMx/eNiTx3nZPhMMcsAl6h
SFP4PZWrW3DI9eYeIlQog3dA1abU4FXO1Mm1kLtyuInUxWZIzwJfvWxZVZ2Du/dh
q6JakRT5hajpO6M4b8Ed8KOHCsURqR5F2LR9WoRZEOIcQpXL22XiKx/xCl2tI8fL
QVj/rVpnksTQSEHiw7R+KgdxE3ryNXZBYgSKLgCYkriQUjHwM/sI4MWj/qQRnF5U
JXA2SpDHmeeR+uGJ7CT3hzQEX3nI9Me7+JYi2Kw7rlEGX2OvnZrGcpy1EAQPitiG
jtHgfQfYP1ZVsmwAcioaEylUC25WzTNP2tOBaoodmzTdw0EXLzh0CPV0hLrBQJHO
WZlh3yYGUyZCsUhTHEiln/7wRNJzhG8UKKCGMiIiFyIDwK7c52SRmgtblSiNgiMj
/kfE87hfX1ldBI3smcErbmC/12Tlrtp1FS5N7gZ360lENowli+Um24bxdHMIi4So
V0wbgt/Dzwa0xFziO7A/5v0orSDozZQUa4amBFw/R81L+q2ib9klwn3xjCPWQleg
hOsqDHEIuCax4mXmb7czRutwMww1Q5xQpCIW31VItUFRCSxwcD92uaTFZPr/u9eR
yhKw81TTKDZMRl+f8NsAtTLp8BKS6SfUKyR/KLcHbmsAJblkMYaIGStnoWEF+lcl
Ur04jnj2Zwmco+Uo6hv8UKsvmu6aIssjzts6iSFoQYD9RWHJxTmQMl0jpc6YVwyD
I/IWom57+iL/eWdvkvl8mPKvOLU6qQhh6SPaYrHHRtudBZgpPGUHZNCTjTG1O3Rn
PRvC7cN+v1wYMPHLMGXxoKwayTHBNsKRIbid3CuSOBSjbdSTw+wpm9NO9xw3AVwc
bMAqSzajU3PzRllQNt3ChGloTUsHgwUyLxehoQl3oPppN/dHPmra9UBCG0XlGbtb
1kQAbT3KOlml/XhspqT28J7UryMFN1FURHt+hRb1HPpGUGddWpVKNDROoPA4xSJI
gA066RewEB377P17pR2oYWjY3U6hTc6VkgBiHfXcWgMJ7cTDa8Lq7TytJSoMZo5z
kxyMLJQBFub6FVZOQPK+p9TaxeIgflV+U//zrLUuHzo9PLmdPy9Fw0364LEcqEW2
PSayuqqxcQImHY7eK9GWx74iLinXG8EXNGNefp5aQfgEAcB8dSX+4JLob3HEVSsx
zdB5gpjYCdA4+isvCsFe+rZB0bBiq4Q09hbaP75VUzsn5VutEmokff8DIoclDv3k
TWN62wL98oxEor9RdRIxKC0U6/Yt+MX5EmWmcmw9+Ka6K4w1JsYU1bBkmm/jv/SL
yIOQeTQuyTcqwED0TMre2N2pDPBPdtFGf0Kz4RF2F+BSYtyseoav1uk5ES2SbJcV
bxF1bNEY1LGTiJeRQ6+ceRE572D48ItDzjzKFfTGQ7TCCjraNWinfugi6urreKPw
eEuHXisB1Hm21jvlpv3cmvWTZ8ZcmfsEWJrAjcUG0CSP2NC7y+XnJU4dmVaibkEk
DxWId2ubtat+h8dTKGtGPxrGQeG7d/sRb31AfwIiG7SnxDlMsvLICVyjiDN0CkMf
vUDMFMoN/T2ZmD9QbTTxO8vcZqWm2ee1haUiN9pb79rHEU1yOWNXSqwthPqHAhY6
y1WufHhrOTrbtsTQkFbP0/co+309JZltRnrulhL9MPc89Nu6aA3VMCFJCCWP+O1i
bxKWUBnwoOEJpqHkkroRJyv4IVReDKDso9ocZkYqYOgn771PH9aaIePqFngAlAY+
0rVghFe8EJPux3bkpumw/I9BdCmjFW0QDYLjsyO2ryg88xuA/rdkpuOBJTQh6S/4
lUNGis8N9SIAc5kYv5Yf7MdgCf0E0GTdIzr+R7ZoS2EspmIonuovsgMGZGcOT6rH
mzwHosn+cwu1xnEa/QWXAUqOhls84yU6ajY/vO9VzCZUgHrc2f7RxwKoua36cczJ
czyXllZRLYqyScgeWY+OZog1XwmOLGke/+puyzxdBXZbWMo2vTOi3vlcVCApZL0N
6INGRLWQo2bFZ4LnbTx9ldsCYAyKFndD/qO3HIks2pHfbOWOnmtrQVeQVXRu9Arq
ZkE+eWeZLm0mbO6HcRlHnzDpslAWsTTqBiuKNBDQMAg0kEjHE6FLJYHdtbLGNsAS
s9c9QkMVaBMEwjkdeB0CV0/Z9dF726yjQjuzuBw6EgNb7gFjkBGAvgpiS2jDVpoa
PPW3SdRLkSxKCu7vNP51XB97CSgc8tVk9LW0S16dmaisDfh9uKPLJG8iXG7AVMRU
cbyyCZGijtdLpgLZJC4a+ss6U4eGDvPFBy17JA+qQCpRbP9lUu80eeBbMnjeh17P
HH97WVgYJdaNCILZxU7F+Mc3RXXpalURCbdgaHABzutdOSwBA+VyVrG6qhZMt75j
6ipc6DV60MnaDrEMLfd6XyccQRTBBxf2Bisn8bKWb2rpXWydWLj1dmI3/jPm5ztS
oBMTEyGq79hjccJL54PtDRsO7OA09oEmgtHABZxHG3UUxXHQVc2z2GgmGxdKg3gj
QLXiPSJve3jEMrV5sK2Lh2G2fDkqIJrJBCob3IR9URb1bnhez0rGjKcWmUew3/eo
CmpIlGTEWx93QYpMT11hPXQSqTi4q0G2Ij3Th6saI9KIlFelaKXRe60WFVtvyWz+
XH90GoWWuPuoIDhg+KNqQ7DVgY5D8vVZCcSTr+l/XXBLDxzY+HMUE8heplbwY8nv
EOkm0BP4tvazb8Kp4OKdnQf8R6Y55iV+dAti886K8QqR+LAURyfDS2h3m+Ar93Hg
ugSyyJRuZl6CPyEkiYffHPAn5eB1DMtiyIq8P3afgddwjJH0r5ibkXx5O0LCFHe7
+0UjlfNfKfE5ZwKGmaalYJKRA8pQDdRVqqU1ntFZCjiMKvaxdDlAoB7IWEeTs38A
FuxkyEJONiz+xzCSAR5FS0yBTQB2aP12fsxCluM1KCws4pc7glC/MSJvHWFtn5bb
FvCCSEGt39MgVlfwF1JJ7HR/mCko5kTrNPKECKtcTxpZlZXA4oCj+frDdJKUV0cO
7ADhnwRNH/48jBwnW1n4woPtfTTVpcUvp78hT0twlqSP0NEaVR+KUPl+ifAiI9eX
7b8zBR5lpbT74W3Opg6A13BCuGp8g4/p1fXblTyj1Ea26dqeFShMkzsQX2zLbAYQ
/4Vepon5AZY9qSpywWociTlPOQzVK68Fns5DP1qc9Gu91UmQNmfcBKKMOtVzMTJF
KkHGdUcbA1+1f6ES055g21qhoYAKCT85rb5Fzj97QOS5Sbji+Hl9NIcrKv4TNG/b
KT/7giYkBlKkvjvXw59BWx3igLU0R9UPsh2P/yHVAntqgvK+g+D5CV9yhKlzJuHW
b02NXit+wNVJFwJFdlTYZYLPeT9B9KVH6I+qjyZ8500K7AjSDgXs2/MlqpHmT2dq
YqMtxWUnBoPQtzxq0I3Ob7vk7uw4AGO2rSLIQvL2A1SUEmtDAKF51LVtTwdN7gCr
3NcvBfbe/i74RF8Rv6TadTGdDT6JXtyjyFphVxeXkLyXdSUV70SxaDNlBTDsym+Y
jLyJNgTcN1CLu3Fx7vaLtXcqXXHesDWC+1gWAX1vElef7LMc9NrBz7OPWnWJ5cuW
t17RAReyI8J/EheEvbC2PY3eMwQrHAdDycjUOzjw0/3cLCvPKNoipV8x6b4rt2yr
nNain01tE5dkil1n/ipSQSVQmOJwREvHUvrSnA3xbpp16HarZCAoXF3cBMS2MPbR
/vVVlik0EasKy0wHky5r0qv+YClUjIIeVK0YNL2XqTQQgHRAFYtz7KwucZLD6qwc
PUZ8IQ4pOuCFAzzD5ou+fAbKwDqfBjpP9EqvSmn90jYdtF3EiOqBot8UZtw3SNXZ
zRRgnHumEC/4E/9koGyaII5R1tZKZbLj4tq2SSTLvZ3AvTorsLaBST60ZM7zy6Vz
UDv8TxIsJiAKDbscejZHn1TPcfDvD+qBif+vtMCqKhiCryfLbviz2fz/xtFxdB+S
bpYTveYSPxwjoieJa68DZehvXxgEspCxHl2SA5btQjJVq4K9m0ElW0YdfktbVphm
o19kNzR8XBDK5i5ReuDpnCqtx+T+vdNZRztaOICFwjw1lDdnqXe4CMeh+ZC6Wd2U
kB+CtH6KhHL3FnajaySTxXedLu9x3ihgEus2kuoK97sO4gnli1L8WE3hCT/4Riv+
93b35ojl8o6TqNJyubGhUqmp5WsXRGYxaKcKfAm/MoszykhgGN4bC4AT41Ji1lc5
4ilq7ihof0zlpS5bk6bXsQvxmPOlVrT7lPOQboiFf/BIXdK8hThbpI5XHRQi7pW2
aG749cYfcvhCx+bubq3t5IJk42t+xuHyPYO+MlD1glmi35UU+dbpxoqIeUaFQYZo
9igPumCKe/0p3RzXt4FtMPmkJWRUm+VPfBbdkfh7BI9KxTWUxtWcT0Ai1rJ4F9qr
QfYQntZJRuBVDBF08zEaWUwAin9l2whTZXbezphbPoX5MSisbduI67BN4DtvhIvL
TjeZVZQFDlm9NNElvbUV+41RU6bzv0PaO7NwUKFoVTlbZpZ5u+FFF72WRrgvNCbH
9tHfSW1QGOQOh1TnPsp9CB+VPoVfPeEXAYoz0QsC99pKEgGkmg9hXeOQd3Tq45M1
UC+kQAeP9rHQ39SC2yNVioylsWCoMP8D/u4bnFx4MTnFgRx9wfkQYemXMQ8XdO65
VpmeWKBteBAKYwTOhWiBY7KeQ6onriXe22uuW60GoSSUS+ETZisBh9TQX8TYNjyk
UhMKUEhT7ezXcMeqifcENXfVraKyIgCqKvBv359RWAQmh3V630vKPOcLirLvTDSC
K6X19OWglVNvGLT+3uwi4WzQQ887pJ7RPSzmaesVqydpV17mhz0mCMp1D3iKrSpU
zb9U2zhvY+//Ve7m1wYx47OEuZzvQKGLuC14Bsdi4wyl/Thke9SOFhpsphiPwMF2
UQVz13HbtRFvEHcd+fC9fD6iddct9VSGBPIRukNG4St9p72rJXzoN55dm0CUxAFZ
i+VNbSsEpYaC7CJgcgMWu/r/qaREk8ZjnxQFrfM+ZTXn+NSn4kMU0VVEJic3kLQn
d+uNnVng92pO8HM1UI6cLXCnqcFwZOnhzS75Uq4mZjs86B2SB7b0MJoHHeC0GEXt
e1nISGvTBTFN0lMeygOxE3MOOGdOK4RTNg2dRuTX+4HN4GevkFlUoiqlPwdoEXPc
PSJAUfAgM2xFYLq6m/koutit3WFZzVik3hVAzaqtW/jx0f7X8VRL2dog28iU3Msk
01uLD+xdCWXTiZ0wohIGpn5zgW13J6RzsapJIqR2aMdPvmmg4oriDVof85XPY5o7
2wIOTCeS8cs912DbUz9lgFVWxd5VuYN4sfKh/5WtgrKWYEhGQzQbxHuvKynybQyP
GsHi5COOvZgt8MSBOMYp7OY5fWidXyCm5VDESX/9ZKKaNYw/yfHHc+LFSmySuP3y
KzLi54Cp4dj3gzMlxvSImlrkPflgSTgknoa7RST7sh+htnOz/EVo4qI7TRPC4oFy
vFCNWosDlhreNGj/QIlU5pxNwBU6rZ23RIXXGFhFugoU30ab+mN0NtGoqo+LOfXC
VgXYwbhajjh5c7oI+5MZrD82sHRp4PCKp+yy/LgkMaIVamNaoWDMVASxIdEngAJ2
EtkqYBF2fKth9Sso3/b+vTOb10xV85Ci6HoJZ9oJTimkobWhJLznLQUeyRH6IGdM
rl1NRdNlXJsFSjY8PymdYikPsnWIl0U4wdbVAOTGsCx8sDwsFnQA33346PjgQ21+
VtwmPf3Ip2iGcdRN/PtVt1/WEk3iFdxajAQiE4CjGurCo5KVOgI2vLMTPw5SuhjJ
VRdQyaVuSIs66Riy3evMOnzolz4NTiGELTYngKQ/ubGKxIQHsAUPksZ98AE/Iyue
rrI7OCMpZMjUcKgLbJO0lrA9UHocUitdUizAJ/TTW60ERpj5lklveF7pEKrNqN3G
/FBXEHc1lGvWS42S5CNIQVvlj6oQYDOvlfoIbw8rrxqA+WnAufXu9wjxzUOs+DGF
aHoxDJ9CFVt9E+OCZLXoF1rL1z8GJwaJS+JGEDMORdcHuIbMsnRO5wwYMb60M5R+
FnMlculHG96XZDXDNWefGlFv5MrcdvZTUsgYZUC6W33L+Xetzk9Z6I/SBM+asVSZ
lmY39fBb5Jp697rrCGupWy5C66PkfYIP7Ny4i9COb7aD/LiiJjF7bK0a7+oodMBV
MAh2yuLE2pV3+ZC4KU6JnTUDPqLmwLXvz+5sgvWHed+kOkosM/nMWFrKcdKP50mr
M1PaPzm0VFDxCTElNpqDinGHVBIY6TyGjuGu9X29gmYmD2J812DXQPd2SzQQudWp
quvVsuma7a/KYpkWPrCdJXawpYyjn6mx0gsczmx4+JogS+nHU56v3mIjPw6QUhEy
V22zrKe1RLHu/ErLi9k1/TKqiCtq6w95/5CoBfTicYQdDldHm0aWvy0gQVRr1q8k
ebTpSfTvSuIJNaRfSMRiZgKelkq/fqgf8M+x7qGHGI9aUY82V71MsPh7JeyXvkvw
HCBHdrZB3w7ufSI3hJmLF0PcInHNOxWuNMBY26c0dQmYw2S6j9PG33KgzZGufNEE
6jrSV41vOm2YCePgcrya/ZpGyMD+nhCuyzzINkvoHy++MNc4jKkI3hoiLRbWOKHc
BvJDzqp/HqLOC8Wf81erRMo9FKd7HoHIejCw1H74mjabrrqbYUp4D+wdT5OdIJpn
S20vBptX/GDdweBDaKm6ucWtxNCOsZvp5HIv7OvKEZ+RC8g5jE0N+H1XB8Fupn0K
DkyXt0zMe/66K3wyrmFaNFxAIdl0cSvAu1b285ZZZuf/HdHS6kLwh64DGyCVC7WN
KlYXUSfBHIoYQ3Y3IPFAISVzZ6Clf0g7eP2rYWLF0k4ALU8INX3JzYF3IguTc5cx
QsX0UuqH9IG6sl40EMLZfB3TdU6OlxeClD+fpDlbhJDuHHe39+XQyQInlUVmEThM
tyKMqCDMIgZoq0vjhXUIrykxqpbd0XncCSCGyQ0EBsyyAz8HKNZF2wt9iIO4KMHa
ManQ9k4HfuixXhExVmd/QawhTUBeDpNCcFWIVHmZ3dgHnKzV+Yi35Vt85nmlWArf
ABueigUG1UQfIR7I1DE0xy3/oYGEK3rufKZzEvNQwatSaSFbBYpwgSc62qk5Y9Q9
OmBvcvK/IBOgIhmPJsG4pWobIls5bHNzIgw8o238gUJv29eaJic39XlQUT6jk1p7
Bf22fjCY8xA5Uii9W4MWr8EF7LO3ewZOKjfWneifSp4FYOMskbmkPF5yCSMJRnsB
x9+BBSQZ0ngHiR7QfV8uIRDmUsPFG20x2XTV2BoGXqZX+FSx5y1Wj/YmD7vYgpF9
4jPpMz5883Jm4dR3lzqLb4vs9Mrr0thvcDtzevrINcmsAyboQToKXdulpKRDEIp5
unrD18Dyvri0S3KkeCasfSqOf9eeHmNH8pfY1+Z24GHAhldq7njQhnug8K+R2q/7
oiCI52labRKmpJNN24wxoUMFyjeNtffc0oprYbwWSSuLVLh+A57eK3aN4sgfJtdK
356II2V7lcuV28CQAIc8aYiJ1ui/oL3L5O9PzxGHZ38x3u55F/zFsGlAQSfmr2cK
2Fjvy+Gt5OKrOUsQUQ3f+Waot7Z3tVhFpjAkleqvpVjsahrgt3FnKF1JZ3K/aOaL
wQhqpX4cOBPvlepyhs/asCDxnKSodXfVwM6tzIpSB31kxI4Fomqe1RBQ4DxdvU48
5ecv5uMXsX6ydedpZpnKpwcDhmJkGFhrBr91fkG5t5a0a+P32qBYryxEQuBapKAV
VX/+g8162xdOrsyQiKi08xa5/hZz0VZo8xPA7HbXfRSMHuXie0gwEC4cV7csbjMk
wS7AIIqT9A3ZZa1tFD4Vn+CbDuXGh9LAkktdxdm2gOKAlBsUyWhruUVOXB/gA3N7
fVxW3t7AAiLU+wUKcI2aNIkERbZsKnuY4a4LsqzlsdoFY93yLX2ijUPFBgYWLB14
RJgouVk4iPKyNmQEh0aWQtEnoeYx0RM7qzuX70Dz3oKSJIFLQK6cdOHiigMUKkZS
9xmorGJV8fnlmvodIo1oYQB5eECptElMsQ2dWTUUSUTpnSpsE2ims2mI6Bv0DOq5
T3vyzEeJKIOh8yS2ZOElklpL19Gces+zkUg8be7A2CyUx4ENX1q4cC9xqop0zlDp
S2ZZ93Ikxk81ud1IE5V15PD7sTz2ALQKSOEV2PfBmif+oPAVQcdVavHgc/4MC/bN
VeHOPcjiunrzVoxP+HOS94WncQulvTeUOT2VjJ9WaNytiHfVXkXE2EmUG09ekLk9
bWdIcQVWlO/wEloZoLZOoe92zEa8bia2HfP07blJ55kDrCkSbkQTIvS4pEEwbe/r
T6IdLHbHaTUI+uPZUAnluOndDupbckqt8GbB5jwXb2AihyeGIz3vY6ce+ceP1NYS
6EyQxOpPycIjJxsOF6PjORym38COGdnScGeVAjav/HqljjdEuTiswDHej+GsQdbF
HafhVbDdOG4c/Z3DTrehla7WCtGcyqVZ5zT0NMeNhXQpJiF811IdYj97mmONoIsH
djD/y58WbAFry+7VO/1NOyN30Yc5+boCN12IddFeCM4kvOID/KFXcvbTV5ik+qQ6
5pU6HpBQk0FHPwscjthQ2YU42ugqmH3wc1ygKvtfjEBYf6Q8KQ+/WKANcReY4R51
PQRR78frpVaT0NjwJoaLXCXpIlOAKL70KS0Fozjm1RCMBl7rxuZPJcteeJbbxsMQ
PAFwCgP4UbaIWAlDcrm8J4SXtnddEFmUDNslkqKZ4Lsm9ouA2nc4YFlor0Hw+5Ai
a7OQOBauihFRArgIK7HXPAq0825UfYSDl3SdbgJ/vDARPGA1KQsTdyhheyL3+UKE
y9GT1MXC0bxeoSmSnfx/nSQe3EDYGeyzbtutCpScakhb9MW0UTZMG1e50XQlCluT
0oZhOwDh6Pjacxw8WorIUinf0b1AU766fN/Sqsi4I/NOO+0UAeRNdkILrem2ZVmY
pUm6zCPzwgV3QhC+0WUnYzrVDCZkhaxzvI6MMrP+b9eoTLEZ64Z2wRCG1xe8a1as
IHNw/OvmC9Wp+0PKimOyOl7BUhyP0O9ktCqA4NZdRhlKjeKJG0/1LAosmaYYs5Wi
D++T+kJyrO72Cx6B1CAbGCFbQRqgfMAOrrb+ojDJjTk7owBeFe1EBjhlBR34ZK3/
2+/UZEkNTtWjj6zH9VDFwjDnuBRNeZM3CaOLYEn41DJ30VWS9fP4I5/EHBnAn4gW
nGYQ+WSVqd+wxUs0kqFj44laVu4F09GMusVZhm+9j6NpU48KquZBEShmUDKaHazM
YmtCGsUfJtOK/hoKXifw4iWwdPToFO5OTgaCil+dkVd7d7c5VeAqcFoZZdd4oUTE
/Yk3DyPGEJsQ7YCalq6J6173p2EYfD3Bg1oiuWjev2cm/+vWyULsaMomHnEoStx8
geSb/cI5s/9JHeZDsydeJqw3DWro9urLLIj9TEFh4cGblXQp3dtU/hsYKCaTK223
4ZdmEPP4L3K0z021XuD7cAhtuu5o0W3XAow6jgorNl2ULI08hVbb+WzmqZ8iTeMn
Mz+5RthruCdQFe+xa2MxexExaH4nznI8yyRnzm+PdCAfqf859Fqkvfk0R2wqE1bN
Icv+W3NYKCpHROGKFvJCWyOTF0q5NV79KMy5gIyQ9WYpWOpTfPltnbWV+WAjomyS
Rhzc296MJFvRlAzFcV8/J45QJ4dqVu8NS77CI2BFxzTcrG3DIT1aAykrsDtryKJP
i0kcu9y19euR2/EWqpTHInwLZYSucG2VjTTZxZzzeXaP8AaIcHQgeA9A4eOeE91Q
UVeCm3A7eq4UJJ+hvx/JOAUgP/5ww6+gc+C+q92C+80vclBVj5nM47DL12qhhoD5
OPkMv7mTFlVtwO4IQGlJfRqo3oN+bKGIXv1HIe/x5aGGARNSR7rVZX40tspC33tQ
+vMaFVS84vnUECjAq7C04ggE/pafbRR54O2bZk9XQWGhLOpvoGR4U7iJVmjfCsVK
ARughRAWuNU1zfXKQMeirLXhfpfHR83qTDOBLu6iKzD7ddleyLD2xvSMTL56hDXK
rmBGDnXPf/vhh9t4pOgK4XzslheOgFfmtfTCpFWVjHwIiJ9sdddrgkBM86+/T+M2
conB4OxuLYB/rthmOrwFyKYH68DGhhET+JGzV5E6LwJ4o9OEGbVHbuAmmBfOfQSX
Fv2OyxQ8STm7WE2U8xPyUbe+H4fxTjKJWWbBtoy1sUPVlScbccmaK2kt5vhLugWL
4IDJ6L8ABratRTIVindOBHTbCOaZHweoJddBP63IiuKLZ2D0VWFwjjUU51Hsj/uE
12b3Jlc7joCMNnlaQoafci+SbpGfNSQZSxhl5kEMHaZRn4huvmeDs2rJRvuEtPOT
sVkPGPAC8ZO/45pE6aY6GsBtM9xPfaHU8nXRMINZx2fCPx9aPlfGnAA/BXk2r3cg
WtJzJPXVktew2tbLtIyTbGrnhksKBYSlJrMbe2aChC/dW+2dKFRr7KtBpAjoEt5p
RqVsK9ximyQxrubRkE9DBJhNxSyGzDEIZ+fe4GEWuO9HvLRJD/XaLbrfGQC/Qdbn
7R+d33VROJ5yCGHt1OUvn9oV8lD+IaKqpQK6SNg4FmMrNVizK7UHQ3nMKGOiWO9h
K49ce1Q6ldPT6R0aI333jlsGEVuRT2H9OujAMJGoEhEX6q7U0e4CcD532MZISS5C
tPkay3U3KtRcwGTcq9hBiLCaZGXUaETHnl7rW4KoSXgOl2Mxq6aaZmJfu1Nqdjfq
ZjqV186FGABmQdqkXSV+5MBC9yp8ESpZuMrWDdeckUuaVjk5pDGvNRDF9rOTFenv
llM0DwcfiCGd8/OQTUAc/JT0i4DqjSsEVYe/XJU2o8jZDUl0uzK3TOtQmSWisMKk
fLzEOG7MSOdHy6QCNPIyPn1OB84dCgAf2rHDTptkDTL3SHBYBaVz6MUpP5k8GJNA
LydQLnmffbHqZATVqEGBowDax9rXC5i3DcRCCFPOSJXgaT6FACyXiqFqyv1Y/8Yd
O6s6YhIzfEuY98KBG2H38PKhUyw9uhGol3iPWx87pS6hcCb5MHQk2b7tReKiXp6O
dOypxjJvNIGKFP235cxoKpYNYVr+QMIGwkTLUZnhHbly5g1Hm2205y4IT2HY0R3N
6AOlkz/l8PJwPZRwyo+tGEr70QhMIf//Y8xesrRoxyNTEU5sRFs9BX7Xc3QCQOAw
YZO5tsIiNxTM/ma7J7S0obpXkxc0eIwwHanPnNjnP6IjNX/1vuoiGEEnQRmNpeoj
Plo89OJftFyqwH+C+RWONwrLwT/HPkKExdC8eBN/Q25CvHiENKdGjHXlAqGO20O0
YMC/4SREfyqr3Se37KD3phokHzkmSc1l5hp4kFZmQDvC1O6Ry2vdQaGT1m/uEAT3
U2PuvidNVhhzae/IsC078rozEPah2kapku3rBrs2zoiHuTZLLoSEM1Ge4n0YX5oO
ref0X/N6/XoJRnuQqq2c9jVjkY1xE2yEbwJkQ7JJlinxIM0sotZLvkoBkITB7lur
E5m0P6kF4ThPDJ1zbUyM97MbKHFW8lT1QMhBIF2gCyw4OImZv5eJwELVsx0Etb7/
FOE3PaEroKoQamHEn/Hh1jQt1gJym0/r7uaJQGRNUEPt+2pB0GswlongL0HAuGGz
N2ZCGYzXUJvN0LIABhrXgsHZWrH0lbrsV5aiK9VGEoKLdUJm7gQXMLGDyEr3qVQn
oW5yeE5u+eh+6W8NaVRADqyltUW13zq3V8RgKZtbNbM2lYbOgmn9PTkgkqQ8MpSL
WX7d3FHOntaiHK2gud7M6PHq4tsPMKSTklAEsie1PXURRBKYRxLYHTSWuVo0N0nF
qRM51M1zFCCPAGXjewbWrJsibwFTwQxmYWHR52reGm49TNGIKvELQR2KSCXscA6+
yfYUMYJUYzPdzn0T0zTMng65J8Qa/Wtmu7WTVRDpIn0cn8W6F9phac5HrDAokSkN
wT9VcsZPmYYc3ZJZd1k7QvoDQnLJMzwIjpoNvuZtPnwXpymZ0GCF4mD/7XqqY5AQ
StTJ89SRTgmla1212Wq73G//AT1di6c2iLLbUELx9CzTVNVFJLRgUCh8DdQmqizE
9hosHs9mjnJ4jLOoWhdWxCpVhquzaYAEfRFVfoMJZXnTllvDlXA2T11CqytEZf0v
iH2a4nKgBN3rB23JVn9PMDjeh+IcOMVd3gHp+E6+kTTxe9LMTTAxXB98AaCRzGQZ
LWTT7XI5ph9A6UbnxuKsFmowDDEo2L2yVWIwN4c606HyZ7SH99znJHSwh0nFN0Ok
72Q86vYj2dmlF+7VInR01DOGeClNyaEOptOeXwdIQl/Jcp6/oYrH1sxKdl60fBAE
Q7DXxva5+iwOjfTSwYR99zCMn5nQiMoqRwdGyhD+UGJggz04XbVy7hEg9hKPWZIU
7hAhqnemtsqZhzXEbZ2eXlSvlzHpcRsnLZduHVo1Yf064POa/HDuqbdvLg5FSLXR
YcBQlQ1i9+qtrrVVVtXxOk1K1saMO0DZMImRugwXHnl8e3Ak4UTeC7tliLrvt7JB
Lt63NXbWE8gy2l2X+F2+Krs0uEE1OaK/DT/QulCjJEHLGwIrzkzyrIpPmQ8OPd5I
TG8D9uCmS7AMM8EfqedULWT5jY79jAcuE55xS+pwdkxz60gUMQYEiigSaJ00J3Z8
BSEYVvFK4EJtaY7+GpcQ3+CyNBzw0f1QAV+/iD/Z9YQbSNyJQWPgQ8vBiSPE8tEy
9k0W9rS0GskT9Gk70zKhJ14pRb7VUvn9y7aGlBJ9/9X89e/jQothWLtGqlmKI013
swwkRWiIp6qvKevZBi3/Jj414J1uk02p+U70JbaQyWoFqSu6hPruERTYSz/X+9iI
dvT0YMODDSJYx0+h/daQVDdrz7VcN2JB+DUIMNhGKvCmoCxasTj0qWuOM2HBDB7Q
mW1l5XHdqe8kiyzvqgNFltKbVJ+w4tlE19BoXAjj26iNjty2HlKEM30QXgaEMPFA
sb/XY9Xfd6bQSujQO7JAgyzjnFXbpBYiqoojpalUJIerYA1q8I2vxlOkWcUYckZ9
A0CXuJ1BIGly7u4WGlhbYjvi1PKtZ+zs3TrepHq+YmiqC03wntdyyDYHaAUjq16M
CLXmLVsv6kFI5W+5wft5gLI2e/CZN+0mhC4e2DAfWyxgmtQh2aAJh+q87IbYLeTZ
VajReRvc3SQPftnVBNBHGtz/kELY49pWmhGoxtsngxdvkxMWe605snEwQQ4mFPCX
YQGxdXsHuSM+/VlEyTzm1PxcCcyOi/a/8zsf4hLIMjxaQzL3xy+bq5+3mK6b3taO
2nRajIOPqOZFu1jxS/J+j40nXTS1eDyt1bOJDW1nCjRVLtkW7PVC6yGZBxuVsFxN
Z/eEnUH9YUTF1UZUCHttiN5PB9r6MHKW1Vks6U99N1i3MfLE3ByKYBzGofhRYiEx
vNirid0sdVAPDxzSerP7ANJG5e4se5W1OKGszmLIsutwQOzYR/fHMowIqCqTsPbf
I0dD4geSkNdpaa3LyFzWtmvNoxTKNt/3FGzQ2EH3+NOVR12E5KYQZd8MtiPYUurX
n2iD0vQiTh/rJBQ4NB464cY/uKAqlS/xBCTG1kGao+kEXzMFe4FYKVSu1xGx8MCe
9wEeyBP4sMWouE2jsZ8vW8QRx+0hGSv746tge4wqXpsNmrfWaso2oKAQ957jeBfa
xRMliPLjYeXJ53mObs2LnfwyxcyrrDimpC7g9y+Y4lwsEdbBo9em+Gf86q/pcsaU
igSgRyPQpRqNXeMszAxeLKZRq27T8c57w0KyeV7mFQPiF03rZSWKoM1rAKyNlC6g
Hr/AnyYYYVMpdK2ZgXd89OIDSJFc8g31laDSQQJzf02LfNcL1zghAJL0IjCWT7PT
4Juikdo1TS0xiJ0nWeoALE/joe2pHhBdUZj9LvdXOD31hQpo4ZVZTLfB32DWIeTf
34Ksir+mp+mbdQIF8lYaqBncEaR2mZE7DoNC1t44J0l5HYtMSDbVQOIHow7grsxE
FmtE6xhMSAlqC/g+Wj0WYOhd3b8OetzANt4xLM43StycePpEy+8kSgreOThytJgu
gd0wcbjj1a42Cne38exDI0x4uaQ4AQE63ExNucEnp1QqR3g+D+gbilw86I4CowyS
/of+/SpS7WEsbuWS7Ax9xZ/bvdLpJ3rR25zN7CMxFoaHzmNuquwa6sT789BK25dB
t+M8Re8DW/wXiTRD8IhnxMPRHXW7qui1dpUiTM7+Ab5wJ+ye4RulP+mOpKLMcTPX
bbBdgK9Mo3S9wiF/BtC7y9QKDkfirZVyKA25k8uSL+lgssIsOCWN91Da0VAKXoKI
UaX1z3CspdgY1PjWDH6wXipQiJxfsEjdxLfa/xUlM4pkxQ2hMtD9Vy8QsOndFmMY
/XKl70CM1zSpc+gXkZTtLtVvrVKyrtHNHOapS0Z3Z1C8TKi0mvo3fCrUTGGalsMQ
jk8D0PdTXkv6iaPK95aDwPS+OF/dY4EU1V8dwR+oXZACDnTv1LzR0xY94d3YHfk7
cEQyHPDpLv1/WE5KmM8sf5F5a+/v5x9C7jCDr0wFEJ/jHES2+n7RVm1K/BqSLzEV
dtqB7mpitfoU+ppmrIErAIfYYOUhG7haAsbzCmvfb1BYW1IlUg7ycn4vMO1K6cI1
qvj0jRxoVUOpQpFPhyMlWCjojI29pxSR5Ss6/SkjOITWhGFKKsHbYEkzt+m+NVHs
gOIzyXdJ1WMIdTEwofqOjCE41NvzOBboRmVK4wqknr8i0IwLwir9mSOLMyyA/y7u
0rgz4q9q8c6aGvP4FIsywY9q7eGemevEdg40rk46qCwK5e9yaocEhFUGqKMNp7+e
uawO4zxrbM010izv8jRr0/VYWhjS49cbqU3MKVsIYDrT2Ao/4G187FMVmIpURuGA
/5HzwpyYTe5qNxsXeo7g4lHBBClR+gj33gfmo0CuP7GQ2IG8ORKDe4A35DN+2zLn
746CTc6U6zLtmRHNy9A24bad+Np64pCTMS6FD9vOWwyjSYx7r14+ilpr20DWKQQ3
2sLGWxShvq/R5Qi9iGRujVa8f9JJvSXe1dhJTYrGLOrRtXA2kPtz0565TF2NGsd0
t+ugh4k1m6dKYyNJLcfNMLBhZXr8JBe/syJWNbDsYIXzpXhcmV6jGojPShbZOYlU
Xey3quGyZce9ng8wRmQt5UQvMV4FVQvC+Zy2vWB3dE4x/V2/PFlZm+IZHceCtrtz
53+O/KFPHn401/AROuiJHfSni00gSWN6eQkutZ9jAHB5SVrAPGgCLW5ASNo9edqZ
jjRm9Xsh9y5LQ5ikjQiqqPkMOxmVv1sgJHQbZJFOc8Tp6fOgtqukh1KsE1GMM4fA
wQodiaxjX5eegED0iEAnT6n96DDfZp8tOsloS2IHfA7Poyj734djdxcx/Dn+/RHz
iTtzgNx4iizeJQGJxk+FwivXwM7cCkMHy5J2euYrkLwkutLCWzr5TaTX8gAe94BU
zTd7iTHUiEkCPQiFErOZ3mR5vahdit5JkFHaYTJE9ywBa+7q62xLJIv5TGSbicVJ
x3A6ug4VQzH2i/J5G4w7X+giQgDLchlglP6wQkB4ZGiq8aNA7XXFun929gfarloz
yjPU5OAOZaatUC16EBMP+7Zzh1XfkdKiYmT9eei1zJ5Aytg2Qhx8p+cUlW4yk0rZ
siTL1jgaAe563m1seVtiVgvmurqgJxcbbo4qvQzZ6tqF4lTO/pTJHJrE013rgF7w
kHmgIe34YIRqJBEkwp8ZopZ3snsJu3eYGSfndmbefJrcuRqi2IOCXNTbSfxXFmVE
u/DQCjmRMrzKvS+n7XydHLK8xtVkMXflzG7EdR5fOCANWdLLfRGFP8BumycqITMb
KKinavaeobvj7f15sLSacobDSPfeE3emDASIlKADvYKb4EzIOt8NMRq4tRq0DRBE
sFjdZbfId14ngbY6Cbxd1aFEM0hnucCqZ5Wn3OxWRfk8sjcZ9gCgnshofioKDImP
ms7AH8ILLBZ6tEC1xqfGSvzN48WQbAgC+hUm6CjwlV4q4mskNDxWBg/fxmLDifOA
C8KVA51wFqqpNo9l3aby3222HFlXPZ5yqVtjuxI6SvSYFPDsNaVhA+3lfj82ZTuW
ET7fTkrsurmIL664Eoi8vJ+WXqQYTq//SQ/KgLH/LhUFCx7nO3FNYk3YIo2nTxl3
1EdFpQTK2RwGICnq1L24BdEB+6oZSWI0eCKV6CQ/9Ck9sDHqov/mZoL9V7NNUxW/
HdSUgZOypYiQ2FqzmHkmwwqpsY/0tQQhMTKrVLSHRd4EbGXwZnmkSwkmrGlwDqSO
kxlE6lzpfDM9yXkYtIQ7t1RBnhEXOvtVRv6p5sLYNq/9pNLa88HZknq8uagvrLYI
g92fETDJFZEa1mlvmnWX2exFCWrwHAElCUFoI7m7R3HR7Wby3Z3URbWLOPEwF1Se
kTKp8p1mjUkbMlzH99lnHDPdLuB+jTsJIJS0kBaEFnfVZPYQFwP+qWirCqYlJ5OB
8I5cfXbCNuS/UnLJEsf4cQOOEbS5reSwHqyxqkeTE6bg2rDu/4zuZ8ss6Z7hAHMT
Aw3xQH8+dND8cRJ/broncLpMBtFhOeygK021/h7/6YiWbQyPOoRjAd+3KrB8qUlL
6qORWP8bmkPlz80gHmTzWPbhEEC/o/PfoWrEZFtUxeEPjA1CCffjlN1m3fVIaxzf
Mv3HCaPYjhr45FFxjmPfst7sczdzTwlvLFJqmI1YukUyORBv9qP8qzpuXYtkyUX6
omXEsqrv37ttS3BI23Ej8NzSWi6j6MAFNTxKUm0BblnlesCEv7hi5Rd0Q5a9zvxD
DrRqzEX70wMVuAEgjmJcpxCtmbnSwsh94fQDTqeKKGiXrGv3QXoGpWStU0VUejvx
d7aLtV617P/9wgWsTDIsBYK/3E17nya1BXwOAuKz1iz20PmpdBm4hCofIEvQFjb7
nLU9hdalcamyGsk6P0vsUTkOIEhCHAI0KJ8JBANhbf7znyF+U3S3b9xII+yIyTz5
bBPVuyaOVp0z7WgCrhbvMBhoC1lXImj7hVwJuLQKbpC6DuRsGfCF1ojOWDchwuYS
886gt9d8eZ0Ng+rIrVPk2rzXLuFDPSjBOU/jRE0CzZJmltgMPPoxMnCu9QcUNLhx
bDKy7Gj5FoSHQojqlH6ceqokwl9Pc4JR9CShByKCPQr/RmczlSBZemDv1WrFLNJ7
M6E7luZ2a4eB8cKA+yLgJ0ZTJ6hOap5jyPaRcgFiCUeltg0xgmJswbb5RmYaQzHl
PpYS5g2X10MGbGRcyhuUetG1NmRDmaCeLHFzc4ZRLlgBDx69aGt8WgLssotY9rkt
ZRy7CRXzOfceYCmb1PcvorFlgivsSoa8HTpROCxop8oIe6O7TF1lgEEmm5fo05Jc
RAo0lazdhGW6ATnhHgQfuifUTMWNBCd69kDBhxIPPCXQlMADNOdj3n8CvZftiU0d
rxnFmY0CvLEzUiogonOrnHNJlDBH1kRXPJl2sy1UNhK5+5nHZRe6gyZbUV521f4h
Zu3u5Y6vrEdU6cut/iruOoyywwThj440342dsMKPmzijdQbuhUu47AZ52cugH8rL
RHNM9Qph1mdxgiJ8di3z46+ForrxbFNJEKkPoIDDgw/+egv7mD1eQotPUjJPXnVs
cHUCQojMltQslbClE8yc2zVbizmK1nv7b2TIzpTciY8uK5SoyrkHRnVP+bc+Co95
CMflOgfoI5ko1VcO1/H4jF4pSpmhKEQC0WzYo3PnJIf4fWmVEm73+WS3aNXPRzq2
rmW7c6lpq5CabqiIbGWKQyiTtrpwLyTl5WsI/XqYHLWbqjEHgwce4A37oYBMVDH2
YIgzWgXVGlTD2omegjmvdw8vCZy53XEYmdjEtbmWmuZvcuCKw/ESSdzTyxEJ7ZZl
ZGWvBORU2pr9Ot/0NYQe4Jb9b0SPp1zRKaErLdlPqFMwRQHhUlwtAYc0VRs3/XDU
12gp7RxFmVweXOjlJLxJk49YtguvsUsxyXwP2nwUGryBBqXiV/LcNYGyJAF3oVBK
bLXfVw7HC+4Sqw/UZ1mMRIhUoDr04bUKbLSPXrVSrpDXttkqvyHBd8KCuf0/REsA
WDcphUSG6Wd8icTHmF8cp3b1/CqY5yOdH90+hZMa6pegust541iOWEYMjfvmE4DX
bshfy4dL5aDVIb2Fx6LYfMJHWkHXcDtZ3oUtyxWxVWyx0B6QkpYhcaylj7bDIZZa
nUk5rBWPqUqYNkbbuYKpIvVQiIfzO/0OZgVhuKA+vqGkadARmXVkgPYwfZYCfVXF
/oUGLnWG4CRdBFAf04gjBcVEEUOFjwlGLrUl9p9svKq+tmXnGjImTaR0jKkJXqGX
gHPox9TJBsP4Nn7oN+itm73sTC4CiAHHxS+fN5p20wzJ6qdVT7QeBcDBAFJQZiss
w1ND9xRl8wxyaBLxJBhf6YJIDThEEgrElRjHehr2D1jqnA8BEc40QZIEzX3Rr8vH
qeJiIXevxoCjC1h9SP4EUn1CmnKpsQNUCVKlx8CwXz28hYQFRiRmxxypNlhPsyhM
nlHAxvMBdQjULHsCyvGmMWR8//Xs4vJB2WRy/Pss/8vyCmvoDRDMjjNLPUmG1k7i
ygqsf9sT7uQc4VL8EDoCvnQ41QgE7wdGAtvEmZVfD3bjG1W1bFOasNujT/D26GRq
Y2ocgPnTJQfhMpC14fdhIiFEEQ5bcIxgQQnCLO8PZRUDo9oShPGN8AyqFnupXLKA
XKxipoUw1odlte5Kf0rLdRHeUTO4et3dGp68cm8hoGBIYWofKzPFATYXXmFXuscL
HD7xMQgGA/zIoAhy00bz/qsui1a7Zdj/hE6ASxZeFuhU3JXRWFltlnWJjmIddGS8
5jR2oL/55SlecG2C549e4/RBraslM9NnkWpd4vaO2RkWgbGnoS81uTg7ec65Zmdi
WOJqeVBIkWRdIdcx+F0HBpylkxYC3uWMmSRIG3MDVyTksf43H/SvV5P26YBHu3sh
nec/7TfRH8u8N8ka2rmOEgUSUU5abLvo4J+qAqYfD9ncmemdE6KmrhSKFivzOVNY
OeKLKQpCOIabbDcEe/rIVuV+LcE2JxXevgmBfFVxTYtSMZ6sfxr9LJuQ5w1BFRyU
YLHPilR7ezHdBsJcKWBZp1+1ebW+zG/+KkVdgo7l5njUTbNLR1MEKqrdjjbNc7zI
WA8H+wEjIE6qKIdhcbdqBS+SX/GKO1bKRlWDKmMHxeMGVAnj0MoZ+obUFJTdwjte
CqkXGo/Nw7ZEHZTp53rfwJGNmucUFHTQXhpc7JCZFwdTAz5xL63L/ofuz7uOVzgq
qzHiHrtGxyZpRiNA5XVoVwQH7U2AyBQ5LNZtNT+li0Yx0cfn83BUqzEo3q4xypMk
zgAanRjuMhuzJkvbD2svTvvk3j4MG31KO+61LAE+qaOs4fMgPcHQ8OpDbKYxOqT0
4AB4MhBHDQcpiF10lr5maBtT7HtoTgCBf5qcdcDsPJG1qdUauUNKiETGNMNoDmxG
WJBAUpI0BI0r391ticNU9IgWfCNEKppZ0jVSJrTSLOo5nPLcsBrdjOyRKXqOZTW0
/XILg2Z1QoPn0mM1267bcJSUnNQ/0jPY/y+VNHj1pPKaRq2XQ6c7lpYypINdlMzU
LncTgbWGzq9XOoFA0DPGj4OdEtYVx3kkPrgoUD6nMCxYRnPYqpyOcXjmc6K3WwNz
rxzi4ljMoMb0IeAK6+SgmrwMwEFVQSKoJH1SwYCW1+jQH8OtPET6P/sZlZJpN23t
GQJcH3xKXIyo2z4Exuqc3LF1bb+w7rHmxn56SWuiXe4zIYh9kABFlvNxq4YKdncG
fgFZLLmgPSL4Oub191ZhwzrVuUuV1PK4ynzTcmkUNFvKRF2p3S4U1MuV2dkQjHAS
CVFNA5l9a3pSlBIUqT/NXeyY8eALOrJ6NUTQSEPpdgIdt5WMOwf/YORSVALtuUeF
v9+zTV116g2Tec1+bY92DQbcipT+Wc1ozejY+3CpLAiJ9+JTNnuUJD0XnQx1GigT
yDNMeTfd8nIoh+rcjX3COr7NpR3/BIimyb/t1PIgChYzs8o9FwFo5i573YPLpAR9
MRtUNdtUOlcr6Foos82jI8sRW20bryBe0LpNew2Byp4fJgHhfK/Yf05/7bOlkWYa
Fe1dEffwBzYJf0BX9vSi+EOZobiokroESPGvOLsCWpS0G08bTOn/fHq/GY9RLdc6
92YEwW4fXfosJxSlwEvAUPIGNE1RagSFZTKhCskOl1ujML0c5W6RZI0Y+GF5NaTL
GIyCH918kHwMWBHNcrLSlHsPpyOtlSRjZE1G25iz6gEH61rFmBNSlUm2QUd2Lkui
1QDlf6b3HAjFxUFqgCDx3d00lnp1v5gFd//Nm3sgYFfld4AvqbOouGkwvMPhmJnN
IZswQRgZU9zp7HBD+dya4Y/ePRGLRmAmbuok/27N4TkKQwxiGcyBeNEuzuQUYSfE
PCCOAqqLVVmCSRX8M4EJSxW480VHxecUKk7HcRCVSpSC00ZVYtX2iKcJIR3SfysA
xDjzW1jemsFuzU/waYRqBXCy24zNQSzps68pIyIVoQr5xKeQYcwTLN++Rh2qCW+6
u9hwgxpSeQXk8cTkzW15M9e5D2s34LYQEfSIxt7bjv1cznAh5wyGIgvg3ikwailv
STYlgn8zOguSi9AUxSBiHR70xdrcDDnoVQsSGoZLx3EJiiK3PdTDGH8Lrdme2AT5
XUcqMRapHML4l6xPDJ0EhtGvuI2fTM+XyM8B5wjZ41+UiHaXvt04u5cohMtBduVf
8yG90sjnrB25/QvYtxAmzv5FsMN/BcI+5AWaBBVOPCQJooo425v29oEgWNxNLKqH
vc0GkpBBFMfN7S+Qs59qBU4AVjXeZLGDQ0HVApn8A+PqF0Uuc7to95evzsnF+Avl
0w5u65TGh0ukX62WXp5Hdny0BBHIgkoc1kNwDM9/1VS/nZAFt/LbaNQ63viifdMe
4l5FBM7gFlm//+yFqMX4bWtO7wCVL2xBWx81T3bPi9XBanN2jwTqnCrvRj6/eOOB
B4QmRrVI4p4EKvkzf6hJ0/2S4wgW4nC86C4IC954Ci7Gs1w9Q+p1WiblPu1VHZqN
9DPljTCZXZ0Vj334TDmCfrdZMbhYW8ZAYsk9BZBMLu5XbUlQrTK54rY28Ak4itcV
G5P10EtksxlNPq+rT29sGtAi9uMWbIlxdedyTbLJj12SNTsH9UZ4JEe+7qFQBTX2
RogWIfHHNXokzp4TYwF9rYk4GHVNKeXUvZ12y76hHH9EQsKvkfhyyDfu0C6x+q7g
1nKAoONdE/vz+AHry9L1otcSIVC04vG9l5WwEJ+ihpTWwkAqMqLpTQklmsC/bpJW
GB8tES1dSS9yC1g6NCS+CsK346vgCF2w2iOb01HBdOdUsA+yNFglj9r+f25fQBxP
aO5YybkoW35WONnHDpWTQk15md5KypD/TXVgdc3NqK19t3uHz4TjQZ61atJw3BGC
C6Sw7tta/5T+wc8f8T/0KG4WXPFkNp1g9+GN2g10IlQ0URhHVCJoaVsbx2essxaC
EDpp8LcARKr2vaT9ZnPQ5Mcy/6OsfF736CIPaztUctDWATDlX5dRoRRfTyjehp99
sGFjGJK5rZxnWSw56TKIOgs2a9i6WIBAQCA4C1FHHURqYsB839TJG5c8g8SS11bD
SHQ4OkhDTxzTK6m21o1AKCjnWKa8XD4smHmlVTZtvmtWSoOJPSTkuLpXDp+d1Xkq
Ndkqzm/vv5gUwrAejblCxgsBru6S39clYqYdz3XRWl3vwTBHEOyOvKaZmzlC455c
BxJxDvFNH+DJtrBoKbiwzAsKVJ39UuH03Spy2AKkgOPh96WL5URoqg8kbPnQfT1Q
WSqsyN0RGwcsgIAv/4de2rDLTQu63DcE13jtb4mccWIKG914YKbPzxUJKQOm870z
xVQz6SUH7WMAm6KSEn2abuBe2ud12c5hjkSWg90/EcvOIVUSvaOALwkiyMIcj2R3
4J38OUJ6zZSFIQZeJPvHAs+Ujie7tFYUGgyYenrtf9gJTOyIMPrdMS8GCL8qYXqG
mbLqADqTqzMFRBGWyDWmHL+ffPj+ng0PJYoc9oBou0BkUlWwibcDASIcyLYvg+Q7
XJo9/ikdBob8d61KUss8h6Hcl8REumxQhQsRCmnGSriFeCPfdir8gzxwMtH//73t
gHtQ2DaAbXB5K9ZuuhhjKjdf1gFlLcWDFaOVOOLz3y1GS595YBFxKsw/6F/mgeLz
GJWg0DD82nVfEWfSTOp+Iz5BDiVFzbzaMjR0+mczsuJuJV0GtvR1r5ErwpQd2wRS
38VbSTwdeSMp5ep228gmuxOST0nh5xPmHsObGJ1LYSwiKNtK0ceRfkOLBcE5umYD
JNxV7nxjAxXISmRx4JvEuwaRgLD97cOGNflyeBsC9SmhhLS7gMRLErRGcFye9zSA
+sp9o1YTT0dubrt6L1jIsAVGrwJepPI4byTbKxMSeo8V8jDQMnMevrmMjjRCMxTB
SsmxjHdIDwECgmHUlnPt1wLXkjOZnj1remsrw/dZQJxi6wFeTf19zV5uzDR1H/kt
i6EOXV6a4z8QzE5vN+W+k2MY+IK5S3sLSDFnqTL+SgmF+Sk0PofSFVNUff6IQLag
E8fPS/H3GA2BwTb/jHsvmDOqaUd5zUMO2v5Uh6iKC0vJyLqXHHJQhUzeS4f9TWTJ
T5MwMHUlFE97utuaRl5EctRdO7cwdhyi7wzEWHKpI6bFW+iDAvziwQN5Gsl7OOD+
s0si6rxaa5/xopRYAPrhPgVV0L2FhDNAQQh2LsVUONHq+fI4zh+o1BQrgm/4HKDQ
tEkuIJeZOI2aLvq8nJn9H5eysb23LpKsPQSLuk9ZMTRXb8D3YFuqV5PN/SKmUhp/
L9BzWrGTPejvI8aDO1g3GVJ+0rnLdGQTpmCF6jK7NDHOv2FlGTWt1KZYziSaCZFE
de4fu9J1PwqjvzOdfuWZYBj654KS8SitVlZHWnu/85T/SBNvuV9gnx0JOWqEhL39
THKFaO1cJtq9AnTXIWSlHWMm+LK4uzn5aI1L1CJ/493v8c5C5IBP9HacHtrp1uy+
Inua6mB/KLjX+2K6CDyZVQtcA6JaWCQkI1Lutm152cafLmmmt+bFbPyarzIhP43p
jr0yyrGbzkkP38wbuMCk2MnJHcQhXRIyGYEqhjjrEPGq+H0bbj60nFVDZCCDYOC6
y7/1QN4KixO7GssAwtKzVsQLsU+xdVLE3ls4Oro2FpM+yJKDZzfHCefa0wCgW9yy
i+6Ah3ExDiywZ26lZUvOFio/zCNeKiNzaeSYWQzZbF7FgFh/4/goCiP5UHjOgnyY
bBUZiZvYRC68AWYVW50djqtuaXvkxEqWqej/p8F7UR8vfbh0/mZi8/wGDX1+gA1a
UXBhbiGV5GhbauAfVvItUW1FkflB3eBrdfn1baGHiwBgkIufMCEgsfBkH8whzGLd
AiHgs5s09CmCojJ6z/xcpGlTVR1eiKXS9Wq45uZZrtRDuLaYKO5srIppPktq1RcO
ef4tDFfNvO6PeQ/DyD3Wuyp81tMGqUui7AIl04hTW8kDp5g6HMs/3dU6k6x2XbQc
dyQF12W1LbzFCQd0MopSuGyEEBopPXEQvLA6OVUIGZ8xoc7mDRjgR3eGRgRaNBUf
pbw0BJqgnL88Vsfz46mHVF4fVTww11Joi/YnyI7G8B6m4zGLJ62TXcUpW9EPGRFc
DbK35m8YM2jjXwkDGA0q4Xd6flJKL6NSaqov/OwltJehwNSruRh16lCJZB6A7ySN
aNLbQZEjdwj8W35rMU3vhXgXjBSNJuHbD4O6Vbhcmhw4HS2zXK3li4brjWPWhZXN
WscjbC0UZ1HS+5WvZZsaZ/p/u60xtQJ2laQnkAbbUU93J/J4+Y6VMsRWp8aq0SQK
gpc+nRATWIwI62AxbjL8M17iWO//tcbhLG0TRhNCZmZxE6zgVtAsvOmWcX+uRjpo
Qr+c4JCbV94VM0kKuWhyzL9HHe32buXXHNrltV17U+8ccWwrByNaFtIrER0lncPQ
E64G340n7ZaKAbBO/cE2qPrm38g70qYRfMhJuKl2wlIfee38Z0lPWoub1EmITJ9L
8j8RO74Vt+siTSyv54p1kELPJ1WgGmVPlWJsbJfG6KcSxCTEs3y4pfNp75VKp3J1
nPCI3X9AoVwn7xAEYtlP5wjdH3phqFin//X/uDSdK86CNb7pwqZWY7CwRwvbFJZ7
BlYX9Cgi1OKKtdazoqkPfdtJOLI7vxzs/57N9GotSvw67z/a6gi9/o+Z9rsU6Jar
eiDOqg/rbc4qK7AYzIW76Rb4IGkpLKTxVa0F3W2i+4HT03sk/4WPXe/vXP7XEm3c
55L6Nv0xEienhTUgy3kjMRS+GXGrRqta9RrmB3vmPY/I8pIv4oF+ScHlTK6uiDOS
4S6USPZv8KC+7jWdj28NiVeFvOoqgDISVqq4DRCYX5TrXDQGQgPpoiwO1s+ws1Ad
Xi3ZQumO1s7J0bAY98s/F4V14HU0qMT2xdrWIQTLCB85dvYwCKLdMba2LvkpXqsD
0Eex7FAdeU1SBTWZA48qMuSCvnzgC1gIkCnliexB1wz1RS82ohNokrMbdEnbB+aX
v1kDh3+tjue/+jtYP/g0cZswwNf1YkJj3se9HEXcvlI4/lUsGBKqyIFoIai1F6w7
acjy0byqS4nerNhVjVzQGUVOUBmUVQDdYtoLCwO11ttmey6Ct+6CVWNb/p9HzGrc
tURuDV4OKrK3iuWtUI45pRWhgzbkRWgAhiDB8VQVcDpz01EEbADWf15bYqLuOkrE
lKlQexwZLps8BmqDrLpIlaKVWJopfMBoWWzmMr3qrvqms6CiHuV4LwXCE+UHc8cs
SJbS+L89oCzu0phNUFiQfA6I9yPChbZVUMfeHde0Q7XLfnU8bWB5ZOKuY1bVYh4I
651gl5cAeBXrmv7OoamZ3dlws3DnRNuZ+fZQEKyvwzNQ6zDzDzi9It351/4iJ7PA
i5GfEWzN8ACj07dEl/DFJeu7+0uNGgFzlzZlJAm/soi636+iSYcwqPEXqpCSp23Y
atJvjLRnTHFkYPfCpWYm9FWCShu7F+TnF19qeL4M6bpSLXIWxAnBdvUcHw+HjXuB
HFOy/KQolyO/xig5vBoe8NJXhCoNqlW0M8wdB5l/P4PSP7ehrY79uyKGK6ngT7nQ
LNsipYCrLVLaOzPZBgToBEbTxnwHDhWYkCRmC3fJM9dl9xYmkQ5wTtgp2hb9EDqs
/TMJQwjNnw3x3s+5eyBthE6iC1Xnzli5O7n/EXArkuaGUDGDEGQl1pJE3vTUUvOb
1bWXFmdvuJQCO3M7Eii/Jpo2SU6mQEmSBMtLwt2oJZ+N8Bm5OjbPFY4EN1P061qu
eHkfe0VrkgFnAdMznzbFn8eoo+yqBYTrEWh9NTu4VaVj2Vnixlq5y9tfq3wVMmgM
AcN8dH21YDlvdddPluhMKhL+dRmYhmEAnzxPuYFccvsdBpDCBh8E8dZcWfaTxakS
5O1kSdY6XL8ixFOwrS8FqARwSrCChQEMxrmzi97BRb3rZsbF+F7zK3bxQ5eSlvzC
K8PPZXc9DNaQ2qDrb6W0LUUuC1EYirYydg0gkRvort8nz1iKpYD9SVy6BRhzbkLJ
sUecSZXj3DWp/8p5Ndm/2/6jAmudxZN9ci/MCTixkImSv/koVomlaie7UDKrbqHk
wukXIjwQ1Iwp2lIW9/AeNBcHXScDEYXDEdCc1h/dZXArw5MFhKP2Ynmo0kkfrb47
KaYFZy3utRGGWNGgdLQdi+xO+5MbyCcGlSr39dJwSUDOK3TzLDnEc4j8uxfytbaF
BjpwDLBmroHoKL+YpY25+6W+YVEnjK6WZJ015PXHl+CUhTbTTv1ImRPL0xLibIQ9
g1+tOYhBtpnUVnIruDJHYNhkQIjKhUcIgmXb/0vu5ETRktFRhpNHiIDaDSEfFz2C
D8A3CbJAWnSJj20I3P5+nm4OMIKr11RRI+YClWdmX1dQwZeNY01WGqjCLgvXh5ZQ
VS6F88kIzUEhFInerif4Lp1Npv9EpWMdExgOkOEairHgfGGpszK2Zwy6NvGHSQkR
p89nuu2wpUPSDL8YZwsxHrMM4IcneD9FfXohBlhvgL8A+26aBoE7xvvf3qmKEgTm
hmbh83+Lu3yixV6803FG0Cr1zcoGd087++t2bjHO1VlA5HWq6voZ882QqkIn6pDC
kEdSDJAWgilbv9pl47SfpPqrFwDhe06MhFO+qYRSZc1ITg2AWa4Y4unwCYVT8OpS
1bUL57b+e/CZ94+OHlfKwUTuOSw27H4pPYPkBjlQIpX13YVlMIeEPyDkof2O+udU
UOxDR3O56Zoys+S5PeJEE0c1EmTeshE1y/8JVLVS1vEK+Hl0uYGEyYoR7waPBmMW
DcBSLyZux5Va/lLNySZZePa8D+LbgNaEy0EB+RQQVQhOHzwzGm6Z7iLFQDRF6EGi
cI1XTOr9VHuTd2eMFEZXpWZSr1cvQPPkNxVARbW23myEismTSCcO9MFoiFfX43k3
UZDCeWspY87uqm9ef4ygdGuE8Q7a+YnFnRqOhU9xndkMnUbJs90yQwnYNlXbfZdq
o60JzIk+NrP6unrnq4PhUtrAHNr4ESVFMgJ8v1vbL1Fe/2Itb8P6jxLzdJQcA8M3
5IzDIY8keL+fudjShWiX4v5+BZH3YR30aFX1kPpXrph3oT+ywdFyy6GhzhtFXmaN
N6Ywpd45GEHRJruFjLlpgGMQacNNTsLWZRERfwLKT+V3aW+LJvLmdl/KJ+ZO6WlN
tCQVc44DewQvbIBQMW/FvvjJzYH6T+8QMsjNM/YGcCNUxWXRHHjqbsPNPREWpRHI
9mmbBbEPcEN8T9ny6iMTZOLc70wsJSZWSi+xdK4WACS9KhsF1f9TU4/SpSnEv4SU
ENZSeV+GOC0Hq732O2AY9yC7RQ6ttCdtFl0Qi5pczY/ntS89jRimd5GktMko6K+V
Zv+qugvt80ycqFHykjo3nWZT6cCWV//D+3WLxi0cpCrcdja7fCJPnLFvvq5KtWyd
0zpbeCvftZdFaLcrMHWsNr9LoK740h73+h73bLn8Rg8QthYQWbA9eLLAqipazqvc
6VFkJ1h11nELevrhL6JXEmedTTcCZWPu5G8Tzq+JjvbRDzw2pqzN/fEHCFSDxypo
nMTwVrmQNX6kbZos4bcEOV/8yNZtDJqw5YCz9t7jOhfwhOLlUIvPx+YmP6fNK78V
+9fVOHV0gkcFx6+Qb2SDjwQiXQ2f0doYVjTtF6f1UgEp268zS/OBL9voGtHgbpig
pz2R53e5pgadMxK2pTUX315Du5KujJ7i3PO4f6JCwnToO4G/gPUBHLjDBVS0ngB2
84JEPAnKgikM7UT2LaPxuPlwXTh1d/EZGpOSVETHTsRjPY2Nrkw4tG4c68JL1ub/
g4/nrOz2yvko82gYFKvmfp3fSPg54RvnVAjhUQ9ZmaPtS/aKUt2mAy8Yce0uYga3
0lOWK6lPzxy/WYvChQnM4wskW/53mLwyEqHC9RZqQsqJ8jQgmn6HyG93Y3uNPUP9
l5NlGPdIAJNnQkmBYUxaGd3ZoCvzW6E4c+D6iWUxOeDaY5IGASaCQkKI4WrAS5Nv
rDQD15qe9+ZlOzUL6DqCEkL9Trq7oztmnRF07CI/PcyxwUlQFkie282GXSQRufby
J0LpCSkeW/Xl7d2onW9yBAR943TvmHpj3CVU9czDYVZ8A2RRPJxFoKWhwDtnHuD1
Y5x8K5kxRjX1rEwz4Ew6k7gmAQRb3+auN0TO9bXoC6Z/O274U30ZHlssUl0N1zOR
XY2uOBMdbqPvLEnF+jafgoHinoaJzFKv42Wb4JY4xmGrxoFJansIblQdmyiINU2x
etKzTjbOLDSyURt3HD3Gv9KjY3w4JLwF8Os9v/1xMeAEFiR2XBr2qbIGjUeDGnGW
fE4ZOLiiSrnq+Q+h1COLKjl0cBPLZDnvZzudtip0uMnH6wrnazcLsk5NzpF4I2RK
tLbTtX0d4lSAviu1Maq5Il5uXZN+hVv89hayzf8C8mWG+h1MGLMrC+dh2iu6NNWd
uf1xJ8sjiQFclv5h1lGGfK6ZgiYMUVgsXEvPgrMjEWZDGgHYwSa1X3koj40H4f1X
aoisfWb5p3KuU5E9tsyJFuauAQ61xakZH+8d7MJFoTzS6OqDyfVlyuLnQJcj4HvW
kqG2Q3MritpQiZlz7nPvistm8stI+8KNj209VUgvjjX6dG9Ku/RgIW8g1oRRD+og
9cYelZX6QFOi0B2u1v3Qh0abtlIpChVaFYAAHje9x2tN+GDZF+r9ubYy7jurn7LY
dtx3PaoElNJDMkUaC5TxWPWsOulLP29P+yEid8fh/SrIDBf8jcYxoE1Ff980U1Ec
Xr1iMcv0jr4jb9BJP8xnDna3dGXM2+d6hJJV7mZkNbV3U/ODSSsd4riFKmd1I28B
Xb7xWz6Xl2vsdVvw6JOtOIl3COrCSA6k+Oxj0+pdhu+RTR/RJ5rlDHhYqx3F/8aD
+zKAEfVAwYwu2XRZOmONkLmvRK91eb8G9O5dFqVaSakLlz12dPB2LDzqiS+to8Qf
TMTDnNhcwFgvwGHXJ+PD/0aSq7Ed7WEEtxK1we5dDMi4Jhj9E3+h3xzoYD7zsD04
Npm3arl4C9sjBMmbdm67KFKHMGMWBFIp0AXgJBdpKvP/Ji4yMei7vE6l7uzvqrHs
Ya6238AMRHg/04SQFGnFrnlcknXZwTNVEUVZL7A46LwuP9ixSCYBEbB6yifXczQ/
goOsz0ke4B2D6up6TCLceNyLN+iiOZud/Bu9hu7gBRATCfWhKceeiqkPUDnidnxh
7mylGV/XJW/zcmaqtQde3GFSfFfJci+NhtMijTW3+xRk+fzsD8lDJV9l7+X5bYVW
qR4sM+iKYzv0vIB/iISpUkAhIAzIbWya6YvnQ6KoBoJm2o+9njRpkN0+53rthT92
Zqrzqm0yfP3xM3AyiuDEIwJuOyurDVtNYkleaN3A6n6PdGQ/OdgyfFMVUCDuniCi
if2OBcglWFCR5GjE8DF23Dqy1Vt3ZtBYZt9ffEtnHXuYbop5ci+hTH1M9HVnJHwq
NbpJOYXiMEudXeZqNZqK/OcehcJk9KVt+ePE/ckqX6tyEl6K4VFqW98hRvT2pYzw
09KLR/nnsGdN+0AA2kWYwk/VsTx5CoYSD9FRAyrKLd9d8L/cbxu6EeJ72FoNeSv4
EkNDlCTv5eKiru3+gYofAGrXJkCKSuI4umdjOHsYs/4MsvXVnTP0y+Y1sOCFo1e/
t0RaAh3NxAdGMUdkcYGpbTiWpChJxrkiziZlxCQah7lh4tHmG+kZEc6QRHp8KAI9
HLm7zo/BKh5g1sqLPQEmdazOovyOOzPs99esPUKkuIPVYXeWfnLixeXLatsm8VsP
A4mer0pji3h/d7rdBg6H0i9N2kPm6MRZdYovlHEvra/l8Vx5WIHFL1lGCrwp8ULw
sUCaTBb+jLxRq85n+IoM/cOQRvZrY89Wk/GWBLkpGhIHhV7PXBXgTsQB+wQbolqq
ibRZIaNmR3DAbLjF49HOBuAKm8bDzk8XVDcpxfXL8QP3zPmmHZlDgbEH4lbga0a2
tjZBm5FTO1dDMciiFD7xzYGDyXaq171iPd/qD3F2o9HiqO1w5k6EkTMPQumgkLlJ
mz459rXF4ugEST+9cIV4ae4lqYMYHCHJa3Stv2ows6AD9ylEhCIQvOIx27weSPoz
39iQnkCAbYudhInVCGkPpWEm1vScQzPEVah4utIku4lmmpFUX8fRSOA065N+KEXP
uVDHPrvPxyYN3/AgOBXG9kY/apUELFMTJywfuprSUjHzn0p4xI07vkJ0DTD39LsP
zf28woe6hNwDk5E2fKFuFrR08aqbBuBYwkYXt/ncMSVLppjw6XnVJzERINW+jDnN
olnqTceASp5ingawNfi+1ATmK2aIpWiu1l2+FywpBG87kW3yPIOKAgVpP1G/LtMQ
VJAGMUlqzkHAJMaJnRDfTLzyhiIfSK629Xo2+JB999LWJ75CL8PbpXyHb2N138n6
6BTZ4xXj3NWW8vvgsuPE02mOA58NQi1kFWpsFuNsCAxqW7d1vr+ahXxQTaUUgwXc
eaK799PLxRvo/FjOVkPM870PLz4gGjqrWXkw/9RQwucjtrWkTTXwIzKD9+VvTsZ8
4XdpzemfKN4wc4k7vtkSeUNxGY9t+okNwsBpaT6PxDbsypS9pbpl+FZNIkibgR7l
nUVobj5fcAhxoDYUuQkrrElzeRO4nQ1L59EfYw2JOGV12VvlKe1zMnWsrWZsZXJn
UUYT1hTKRkwvQf04JSLOm23OT97qEy876q0aGcLNll84mbxGnv5GoG3SYXJKPu1V
d+AzRovSH17GJxH/55tKV6lRoudwqaTN84b3ubpv4+gifAOMBAGlfMAS2genu0bC
u6siCuTu534Eg+9igwkFBrfHdKmQOkov2kjZ/5/qnxyK0TpWZXc2HLF4h5hippLI
ziKAH1eza1oWXiXVnIVStfWgKodBdXHOVn58TMRnpzX5BmfsMO6EaMmSlml5SFV5
t5FEPt18DK8GfTBUiIuhVa9t9HuPoqofv74nJuryky0+Hnm3Q3sxvPLwSgNTM4Cq
47dLrtT8FXdkDYUrA8SVED0Lh21sfD4ZkYXoXf0hy+MG6KlPV6CsiRrvw4aMQMA4
TokuFOg1UMmrJysenigRNVwRFCfNAvlWj9KnEMysClp1YeMv2OPBcvAGTuTiVNF3
bqKXujd0xVMXC2LY+NdbA9iKIICCxCmJRQSw3uDSZo/HhevPCTvFlRrI/AoPhuiu
tZalnITDQ2wf8iTJnhfg/Smd0qCDv5/gEVU8GkUoXY95ZdS18ltSx3T82YBYxazo
t187ZjLX46NbMvOS9ALJe0yDHZ/cL1AWOiP26UniEnTDBFPrlP7S4F4dp6HsXqS4
tsdA6j4v/k70UUd6SmTEmf0eibgzmOT3iSX/E+pnDfQL4vWsd6nCeCsNTTIwB+zb
XwdPiFRVnkhbnBX6ZLGcdv+Pr2jk11RBELlL4cBcvaw76z7tyFPQ4QDqZGviCmSG
z2aldAPPB1BhqUvdn5z/cBU4nWLkZ8H882OT4T8S+5zLFGE3nrxMNfa2SG2yV+vq
0XLi6g0bAfCndPIMuTFDk9UG4iRa+jmkZcuuOc7f8K9HyGI82xbgKcor8x/PftQE
tXQM6Bntw3tPuX/QHCs5SNhmG7nJ5bL9NZvD/Ka+TizDJULnpTCOHwAjAW+VZb+F
+OlIqkPNjyoS1EKvdDtJEURbcAnX16pyqmYh5snFen6B32sdg9AVDy1liGuw+QQT
+8GaMu+JBgW4VCIARYd30OIV4czqhpIhVC79ZcIakw3hrFi5VHsq8tqgPQUHmSbD
GiG+PD+dNv1ZPvnnpJ9GspSsY4nuYlMMZ95AoUQdRP000NUwuWE/I+cFVMAqnJQ7
g9BaQGViYm9su0UBu8BD6OApJl+VhBFghtXlGlv8nPdJyUIUIy9tjgKunMXGunhr
V8jASOwVAzbO8xudGXBYDpdubqbEqoXH/jHXLIcnrP2D7UEKu/bzT/zKgEK+/IbI
pwUwyvhMJImtcWuiEduAuFweYJIzCFQSFVWdsTRfOgQadr6O4LVd7B7hvRGk8YsL
CPZgPjExIgsvSrcj8vkuZ7Fm7LBIYt/lOhzBzasraDdSRW7F7pyzFpkvIA3Vt9QF
GQB4o0lTokfy7mh9u6Gl7AnTjR0KeKeUu2wc6/2yXL0y6f7HQnXMOrJAJE4RqP7q
GarDAhmDZD7NdfY1MmxBgG3RmcOMvhIzYmYCV1fzkU9zg4ZBOhRLAyXizHztq+9v
kMZNaiH6AskkK3Hm8qaTt8UdkzL1TwvXqdBVA0+yrMUll73qJEYX4Z2uDJF1AM5I
NCwJnjYjTj+tdJL98KcIvwTMDYO/BWxIVPv/qCpdPAKqQr7cWGT1kj3vuXrZqtXb
3eNDAfJmKv7ElSNEsUfAY9bdc3pkOm1Uga52ouT9cOSOZXZse+VLNg8fpKIQpUrG
F1VHERzeVoaI+kUMGZetBQD34BOKB0GMKOYlsnpVldgN1U/76TCNDMDkZ9We2z7W
Z2cXFdsoWCahlzjBNWUYtmhecORM2f5PxNGqLqwnAM/6sQeJOeG++gWjuKQZB5rW
C+kkxs+xHf8p3wWoAAbg3LUYc7mx/EPl6X4WrUJxw1Fw3xj2OaqcFm+9tRc87k7s
ULSs3NaX7HNjVYEJwDS58w4KFLVOCu0vXsZMgtc9jU53F0sM3hDWzo1sIwfGORsV
WvfpVInelLs3xcdZxGRkjuCxIwtfgGxAGW3tlOiBa4p8KFQqlu4JyxrO+qyjQUYR
H4fh25/w1Ug8cUNg4I4eApzoybHlh3dYdw+H7gRis97kEnPeGh9ROnFcrWkXvvmq
nEwrT+Ih2TWR5WY3aHb2YmnJ+nGsMPzQbbT6zagYrnDD347cyCjJjdDiNDI38/3u
d1njAZKJy/o6ZJvCEDkmJSQ5dlzNormPYUcDBDGKZgifg6tOoyGNtan9kChFcKKC
tngwWLi44N+dSboYyCBJxt7DTXICWxLSGB4tRSIajlDs4yogNBcZS3i7/o5GzktX
63Zjdgj1+NAr2YzuY2s6tbKCR+63UifPqNV9MtuquwHOEBHoX+wQ2VJDWaddzyKc
q96hhU+cwnEBk7O6Sp+cj3qcscj2wpo6UUoarzgJfy4JZOxljf6ROaVR999pHap+
WYRtfoMb/3le324KgogTLiAid0kZZuWE0drwP6IgLMqxpVqIpBsWhNiGqpbF1sb8
lcOERcbvj1fU3TldxO0B/B6Mn67hOxJbyT9ZWhvuG+XFhfIChxCyA3Q4HB2fruHQ
0/WOr9LiuxJgh/Y2jVh2m5NMAxF6RgT3bTkVsIkP2DCGFml/HD62S7jvzRj3ZNzt
Td2T1ut10qTMV/oHtGLzbsvQRAmU/70zmW4IG6qbubZprg8kGP2cCcp+7iw2HsSw
tP0bHKMGLi7ZHdce2xTu1s6wsk63rRaebLfZjJ5OvbPjAzJLls7IErBZTbCJp/2A
x1mNM1VBVIDXh//WZn6FxlTGOWIf6RywY05j5NcrDk4bWnUchrxa8jW19vTckhum
4lJonzxS2B2jYn0z/PujvxpiKduZrk9U0OjJ5EtikJWpblChgsry8quY+WOn6slS
3AC3ONxyzS6SBT8kLqfr1RqsWmRLXfp+LiuOSjDEs873FRLSa/LR0PFRgaz3cfSp
jOkaK9ocsNgOqdlgZJF/5w85nBCC6wiUTsgx/LYsPm/MaL5up4U5ehhOTEGfa9F6
2MS3AOIjaRufdk8rxrTjLdHoHpH685zaA9pn0g3LirhdZECvBiGw6yf4LhpQF/8B
+3b9QgGJBCjl27zgFSGX2rae6M0De+n+IlXRT1zlvkHg/CktOnw51TR4T2syy5wt
5QjrLECrB79WKqh6a8HXOoNDxgkSpHpaPX4zCRJ5o3yDi3UCY/8kKZRsEskJMRe7
fTitqN20O+Je8HXZLjbaSnc39DOscOsjZy3YOWUwpi+CPVjGbXfS//2jscq0v9G+
3GHiRhF2YPGfQbx0pLCEChCi6FOdDbqLWfiM/ZmAzIQAAp84giBO8y3gt3WsGiuo
xS/NX8cBfMjlmUEm2AJ7d88JkB60CIvRcs+rEQf/2N7Se6CRrzsNpf/CixtU8rgg
K9BlvvdvOmt9j4EqNtGbgFBYOZjvrlBuTwAzgcCf5VaYLCbCDNSvE/RKc8mL2kLS
lazQz3hU6F5ZChBBlSKDmHHyIYuXNtZ3p0S2e1+o0Ha7l1+HedqOrw/UxPSxvLYi
1D0CKWc/BIb8L6vWnyVuyn2C69Jya+ViMvfh/CEt4XRYrJbhYdCBVo7txZ+mTCrW
XeNyBKhy1124pIXpgzDZYZtrgH22wEQ2MLurEkG7AKsQg6ofZV5V+Sd/Wza8hkAH
LOd4VDiJ/cKlBTeqoIUER28LgLdaYj9bChjIvOuVcUkyF+w6I+I4du6qt/UK/7+C
lUJElwOYwJn/PXbIDPEysG25Z0BYjz/Kwc+S2fRwwYE4cbrAe5c1qStjqgNsvd+h
tl3ACtvvS+K7pN6x8bPrAp4IcvwwJwKI9TQxk1Qglvv12+dAC+ahkRcv3ShYZK+7
rywbgv6l7P1TrEGphqsTySxE50a5IGuIJ0Mpf8IgWySCaekd4WPjiliTN2/+RVK+
//jGLxSL/vzhWhoTfIM3KbrP78mDdWWpgkaTmMLTWmNiPQFN499bb4pnXnLNRjHG
5yaN7BHXBNtt/wYV/rNa0ATPvWvjWV06G6W5WbmUyu7nkLVl0m/ln8nMajDfqg9G
Ef2bkF7RO8b+3mYFYdr9EO+OCw18W/8qCLfRiuS7TxDr61ttu52cfsHCaAMB9H31
K08tfFyewqzsD588EAE7ptN107w90d7hOqUvNnshqnk99qBQkYThiWEnWs44TpLO
xLr9rJ6ogIyBdl10SLdK1jpedeuNMYVsXN20L6P3J9yPywFCpd04j29OkoE224mz
u365i8vQVr0A2Kz2Rbf5dHQvYL0nuwTq9p8mERt+LSHwy2yUdoIXEO7fh8CacY9H
YBJACBTUedlwcucU+czlaa41/DaVl/NZg982Q7rwkil+lidEJ2D3lQfV8BTh1CYh
rVRuOf5JXXeZgp+whP+5/Nfym3f2K1c9R/Q498cYgEQDzRqSdgW05e/OmCD7fFhU
jcSgOWdlhN3sHLMVMd7IrTI0GvEqAAyplrMec/0QrnkcsVZPmleKzR+WUcLk3/Jf
KJtXmcA5d8SK99NXAhHddrzajWaO8jj805d0AgUeY8cJwp2auZDwn33bq/wsVl25
UPiy+lqKfgcc3IjhfPNRfBcRdJfrU8mezfNfk4/qrwcI9oYEBvba6kBt30drFrZP
77V1qR0Ao3wlstpV1JJCBP3sLnlRVty8L66rIKaKoUN1l3aYVI7PpH5Pslz0dwe+
40FWzMWA3LUKEGACj4Mp0IteEck70w4HNULIl62y870rSfTBM7p+IVbvfCmrEZ1r
zNLVzrPbLty0fV7cP5ReqXkPT0Tr6KSsnCkVd5zBLdXT4fr9zpFc8OkJ47gXAJWE
T7qbDLSFqhBLdVOOTd2lVC3LP3h3FYYnS7sBIxgUUyLRSbUZfLzyTBNRrFGGxjuU
NHbgZWzzEG1xBo9rl0fSYhJFPZWo4w7bGKrP+0NHhearF7XYewOKrfw3VfLOfR/x
eo/rdNMdwq9Ed4f8vPFB2h5TQNRTRQpmhbUXhAEbcmRR1lBUZ67mPQbdf8hz1nzZ
bv+x7VyN/ifXKWGYPrVOJyqR1pHAuq+bWGX/GSHglTuTawJOie1161/KVXZLCH2L
/mpBbIwFEJZwcOsbShAH0JTCkAp+yoWgpPLoGuFRMfNC+v9f8P+NlMQhKOAHCAvR
cnLaqih3E1CE7h3EwHJ+jsRUcwmrMpRi4JbFfkWTzl4M+WA5tsY1KudEfImJ+Kwy
Ni80V/TK8jbNOrpzOlX00P1P21LAJjypAc0ts37rgUp18KYmtjgnlwKm4YqVwYL0
LHVYeXgg8W7Hzxsce0bUIwaV3yf8ma/uX1GzfN/10ZKVNf0Z8cTi8H+weaASXQcL
zZJDis5VzqOBxYleNJQrrMhfJ4a2i2DUNNxMsIsSa9PGchJhVD39RK3npmLByQTg
dkGMaGdbANTsaO5KMpLvApk9Euwfx9zaNw9MivBfiBbZH+bzP5PBTwXi+vktGQlq
uy7oOfRBL8vWlCcnkb28Ivlsu8scqqnsXvyuB1d1dpSCKbipfWhOwhzzmoTnXGql
Fjd85ZX/MAhOL0+52kkX50CQPTKYc4LgPuoUXFTJQZ2DZpEbcPz2bFSqnD8UnIK8
ZTXpsMUInXcAlF+Y4zbsumivE9PVLBcjKpz4yae+W6hErrcs+Wh5/9oFIspTMW5w
YtWMAmEqOIPpZLYy709gxiyuY7/7ZEg9emwLTE2scQLcvHQ5vf4dQLIMEQGOsMLF
W7FYAzGMNl30XJdJSL2RaS8RIOjt5FIUvQzXFKC/sOPQeCVYW5mnh/R6T+oGRQM7
REoSqSCUDC2vnyWgtMo7xsoV0BYY6hxlgUFHSEFSmBc7hxz4+Mdb+T15SOPpJqe1
b92O+C0w9chpTVH9KlyravxpA9/odq6/e2TgAwM2XlR9MX4z4cg53BXCwmkQDR6M
Dq/5T4Rd8RjZMY2FraBBVaMAUrVKZt6tpQXnsUYYu4CqmBbdAiKdrY/H/WJu+Q/6
a8NS0RFnUdjmIXjkXaN7QsiFljc92CzqHKP3xcnTXEh/O/Jb13WCp1kMsP2cRxih
XyVtLhbXlFT8niBywSXc6cdGgfxvc4FYpEbw0atZtzPkULcD98LeAz8J/S1kw62s
3lQ7a0yaDinx140cfhJakpCvJkxqugFDiaxoH66h4v7xHh/+5SC41zCi+Gc68l37
myT2F6PJ3og7XEeaiwVRCcmwgMHHTnUXKUAlILrmXIZGhXhuX/wnMvrFPoZZt59L
2XNiynUuQuddaiL4Qb6CA1D25vqkPlTB+TZ+/qPihF8WvBjya3vIiIKZqumU/sJN
uAQMQ9YobTNx82mg6zGhHN2HZcfYPWut75/2ZBd4DTwV1FtqNRH2aJ5LTBR8w17M
x17M+giMOeT9XEZOx2HamzuuQcFE++xn5GdfdHIeLBH+XnFKJJPqBjkCujgaHx+y
smpXUvUZ4Y3lTpmvmiGpIW7gW52o9Km3o+PeAIL2iEdNl2ga4nWFfJleq838H7Ud
hWKrvSNwpgTyzoZLikJC0stJztFRWi+5cmViroIMBCPl5o1vB36XpHhHtEewyM8c
ds8JeAAYUTT6oNGtSW9bTkORv2mcS3sNh7wuokKLml6tf4dN2aA7c1swJ4SJSlfh
+d1OfgamsP7iKbes25UFKrtY3tNr20nLnjQTQ6B6lqg0YKlsoyM3O5BtkPS/D+di
CVVd2ynizcW5tU2V8QyxMy9TvWbxapdmnchClSc/9ZPuyMoGQrGOnT4pJeI5lpiN
HpBAxMAhh8856m8TO+wKMzYEuif6COURzBIiV1E8psWnSdiRYJEawcUnEmCr4xaG
3Tf5HdkYNaDIOVVgTxW6hE6zg3RlWmh1aYEZmPNK3D34t8+AfIcQ2cHigBHD8bzk
M9uWCAUbeJEfu6Dj2lMaGJWKn2KOON79jRPE7TIrJUoDOYbVrydy+ElpbckwRE1X
J7MS8vKlwRPov8wKcRgyQNNIOmbJQRfoKh0zMLn7spdz6cS3da2CYYw19Xq3MAm4
ldN7/+17qEU+2bNjY8fJVQVnqB4i+Tvi4eAAfaVeImcQwvSbGngoy3JIwWWEZqQa
pNcZL8ucS8KQbssOpnaGyyvrEX8Y9NAwQvs7s04uhUw8meGANdyh1p3TuzVJgAMy
ESfCBG5IrmHmsZGvkAdZAv5pfR68+AHq3FeqCr0Z8Ho5tx/uaLQiJNBU3wBSX865
xXlTtESr6e/evmdyxZAUXcHXwnH//M5/WLqpaccjZfgAfTYtceXxjvJe2AvvkeiB
Ddo720LJxJWfWYYk5ujGqdt/OZSSEahwqp3t4Id+JJq4F/ApB9mRZmD7RZP1A+Sq
kq96MoCxDNzS3xLnWk5rZUqT6auHSkI9XC1l6z6NJrPNXm3iac1ii1IeYi5D/BIl
waZ0nGdyf4ziJkyob0pE+4FuUNEO+fTM3sxJqDk/RMyyqmIQBIIWjzMFRL65Psq1
26M5eElwivQ8QhxSg6VErVtIUaxOZATm1ZMO8QgWetn9l+ku5MhvK0d7+GOoGV2Q
nIx7mo1fOqrJtjKEXsS+G2XQfbZkUPzFbrIdiNsqmdzEPEEUIewj5cxNW7hmmb0Q
pflhE8NpvOYuB3z0fuvfSTC6TDj/aXAcD8PhlqMfbUMhjSUTgtVYpNY/xX2Duik2
NWu7torZjTpbnZ1XwRCgDvRm6IcKuIs/PYlBH/lc8YXApNLMP+f+aV2gdvUYNMIK
kyFY6pLy8HvaefD1PKzxa/+hXyfah2lmfxocVliIgf7VAfunhBc8VXOLUpflH4Kx
LP2w8Lfg565r86TrL/zsDnbn1QJDzDLBC5NWNN1/GxDr8uLRSA4PylQXUS8YoO86
oaZwm3a3y5GJSktSt3DKN8EwS1smfJ5fdEEeyxLrzmZU76pKHMJp5YL2TEnGo/FJ
EecSS8n/M0jDPW/LjkpcxxkYqoW4xXnx1hdnyO8/pWyd7AITyhPeFJxlk8wz0f2Y
bOktCk2vO6jctifwSfebETu5t93j//mP6vtghfUY+oQxG7IEKbqGE5HAz1VbVmZP
XMxBBJGt/o9peKnpBEKXek88Pob1aNyj3ZrYCX8FSXxWNE/91SGYP7kOVvMNH8pC
x1oVb8/uMe8jAaAjXfN6QSeb6Z8UQIeDsrMkeEN8c4H4zcI4KjzqxwzwWTYkNbtU
sQIPKbIULO2RoP0ihGald5hkRhSc8UGCEYLr51SfspGA9JqCeXFWXqjHYghUDLSP
lD6NWV0I2PY18b/5UvKOrLZT9Uwh7Qk6agBFAdpC/DrVx0h196ksRzcaitpRRR/I
kmkZfERmlM7B/1Q+p878bHkHeDc2Tn3a5ifbTtWz/yLUDgcWyS47awsQny13KOj2
gtlyYfsNCfffgM7pV5JGK2KSfVyYowwM7YD4ZdPBxJX5ad+lF55IX2WPLLNxN5of
cBHhup7oBPPws8Xt5SUmQmjnSJi0WIF0gyDhEzA7XH3TybC4LjJ4/HWK7lv4ix7Q
Zt4xA3mKt5ueSinh54YQtTOx8N0qahylDZ1brCU8R+Ao/9yFqNh0cDBykseo9Y1u
vb5ZeBogIptPyGbvXmcVXGwxFHuXWaW0szcYKG5wdkbolVZgM81wQF7XWr6AkYmp
K2LFURbdrqSkTeyQ7RuPM1mckYciIvp9BnuysMTP88IpsZ/maUcaZ88cfRg9QBC1
RnYgsvJ3bfCmc57eNZ2lurfxMscdmjTPIp6RqSXlbsCfrleqW7q4+LcpbpNerHDN
/mjUr2EEvLqVgcG8842LJnjPZjVMaE0fxqhaQn04ijjE4DEoS4111LZ43T9p7diR
W5LMMHgWFY/1e3ITbwomaHcQGXv7+hyJKrTc/YwioRvwY6lonSKlb4Q99RoPe1tg
BmglJbsgad2FzHzoFqf6jJ/9Jv6fqssX6xNS+QV9BrmQ5XbsrSNhkGjBnrzCEdKV
YyACynqyNFRcMQDafSB8J3J8H6Ux4j+JUgzuMi5z7SiDqasVauMo3h8DI9wCPz8I
9l7NbIPMQLjYkK2rVbp6K1vbRZA1XcdNSp6XHqGBhsOa5y4g40xtVKNi4vyKOxwx
0uOMFldXIAwKBBYhKJHNpi56z9CP0EGM/DpyiC6oqnKf0PB60JRCwbXQ6F98PqyT
SqS2nEl3Fs8yck6GS5tQD3BScOLUafHygeChVj6K//8EE+nlQ/AMqbWdCAVhGMAw
Qjtzp9ZWscm8WgxwpzlWZPOiouK1QrLSO5PfXZJveMue90cO+lbrtkjhFBIz/huf
D8IQcVKNP+V60TYyXDZ81c0j80lmddoM7WlG9TJoBbidSkiNJBj83jyoBkfph8x/
wfyitBaDhvwp/YKhtqYFUwuwppMNw020dd5ar5ISID8w5RKPtR3o/1SOf476MAkQ
lh21iqcDWAvYG9bTOkDaUihuNqCmu/uTsz7GgtEQUAtYrOHUWv9QMSMh1nItSYuy
brXUJnKCKCJAHeyMmr+lNewV9aiMZHIthB1NZ3eNVT2s7rvic4xpXsOWvXcgQM9F
irdEg0TFjphTm37T8Y/zNQ96ou7OCIYcHxkTN2qc3MhrRivcTu1VZr9rAOl8MEMG
LUxRpW0lYWOR2foCd12klB/PKbYG8LGkriSPd0LRk+lOMwTZ+zkvbgfzQBYT3OaB
ww7Fa/a9nsak46ZqeTEkER9W0vzGRKNJoqkVRrDmw8dHe7+qgzPzxWLJZwziw1EF
WC0GnZovUVSFuGnmC4O3wtgDDKVyj0qOxzWgZaxG++zaTb7w1oXBv/KudTJw63mK
ysC7redSSEHpx7EcnlDFclwGw2px3IwAi8OZ/9UnqZFE8XlYXJkxGiUl7LFdPHYo
uNUqk4SjQwLy6TAE0nW2C2lCdfl8Ekg1cA6Zru4DyI92W4oF2svvQV4svHUTqvZ8
RQPVrSBcbHuqPEee3skMaANBYOBnvxnYA6D3AqTcjAO6rFbwzxVD9oL+d25exk2j
ob1MZu1TJ18kvhkIqNb4abp4+VPbGrihxE/UCBZnHBXiYgyNiHq/pQWYY1szIGKc
RbI+Jh73SfKJoLGte4/JEqZYIuUG5icDE7rXmvivPt/Ir03ghGeECwGpkSbxFna2
HhTl/ALaq4yvOpf6ItgbOqg6bT+uBFSufXgFH0QmLvbKis5EvRsN3rT0Y2aSovpZ
Lzph4TBMZRK0ol0N8yuH3j77soM3N/VClrIhQqXgEnWRq07fEKyfhh5pVviWHbSz
4rouK/uPfLdpQ0Xt4mqMfzlvaEAwBNc1re1rtOm8XbgxaVQL7GJieRgB2uMNH7dX
zUAu6Fbat30mesLStnTMaLd0UT510iBbmwFm/Pcv44nZbS3DfNfcfie4r9SiBMVJ
2EXcsuXwrqFlqvuRBMzEXBN5y4UxLrEYaTMeMX9e1eq+HlQrq7wIb9Za3wwx01po
/dfwMGVLYW7RR7fn+MOZnxK6q01+M+FpJAjIAbAbhIHZig+vpNV7EVsH0p8tc4HT
NDqoXCb7PWar484sCNtOerlPKOLkzCT0wjS5EEomjN6XP+OJ7cY0BknWcvjgv2mc
W/0Yunl9+tHaxchPibE8ZCPFoxdSM5mtxhWz+FkQszcyWXtEIs9SjXHbqVLQa9F4
eOlBQkPZxUf/qopcvYJgL99mCS5yXAf9R2P4WHlVpJrMfcShpmlOkC+BmP+VzwBv
Bv+37Q1GSle/PoHjpkUwW75x5jEntvdZD3Y8qK6APT2tttaf1JZIaEB/AdzIAxer
0YGz7L515UYXfos03dVXGjyWocOuf45Wb3THZyxfMy0vzTJKzOlS2SztiYdAaBTJ
TCEo9RhIXVQpsOehGzen1qKGS6ZmMXIknM8Bvo92ZUKP2QDBMXenuIuWzB6sfvKl
d3YVs60UZtIuwIp96TyGDE/Cs2Gg1LJ7Ic0rYKwzYNIaolxmOSRYYaYGohMimwwB
bHEU3LBIJ4WzM5lKOukjSSl/7xGIshqeYTA3gqZILvMYyvHqQm7CuI33MIfkfhZW
EYM16pRD4UdQkOieCwtCesVv3I06rFD9/e7bj0SxCcwgM6Qqcp+15SIlsKpfUijx
AN9Q38mdd+lTUxvCbCFRBsz1jAEbappqzN3IcOwIv5uhCivmbnsA/zs8dG4cxy/w
SrT3jCkHDetZqbXr69XeCe1c+Zq/9+zRn5yxZJgIzCQNTuLyPl1seFXyjfvWkl/A
oJ5dL+be0gwr7aenASGn3PWKKG3dZgjpg+PGSZE1g3xyDVEpbh19dEZtopw6W0xe
dhJAoa7spnK45IOALqcv483J3eHMd2QxIywZqp3KgQp/bsr0+X5qlWTebMcMzJNF
xxATl2qqO2je8vI+pf+MlM48iU0nHaunwvYJQ7JdfvfWoiCPtATW1mCQcYV/51Py
GEAJCALYYetXe6El4BiG0PexGwMm6eqTGWAHwkyNRwkqjh6WFhoNiO7uN+fkq1pO
TFq+WA/+tldC5Zqx3js0+HrtgrCiCndWTFzcfzOf1TkYNFodSuIyXlXz7S14Moor
xUggKrkUIbMzVv/ggy3RMW3IWmGmX2XkwQ0+iId4pyYvQb6fDi6pAd83pxquyjVx
Y6tWWFff2+jHWPYYcnN8hUxgDBYlJR66VxMMlQDHeUqNx+bLI9Fr08EGnzD8XYIm
P0P8YAuQulB6IbzgsawLxUjG4cbPGS5jeXw7mzx3XD35M83KQIkky42C3yMTgvtZ
r7NHEdL7UbOg1Fl16eReAqM/JzwPUmiDSH/qOrYdGDVO0HLqEGCvA/uK0svLAkUo
dCUKWs45It1HPLqnra2RlJxS9+KpBfh7WNmJSTQZhnZxnjUG7xUhelsLlT4JPXDg
5w1u9UnIfvAYJtNBTea53kbiABuqVgldtqblR2GJDb1gNrCOgCElF04lvdBU5Qh6
5/diRmhoNeEML9R0qdffg6xnav9o/PGoNwHCHjW+eioq/DX4/jJAeVr3gp1R2tdP
x1puPPhCJyeytVikpiFX8ljFZeMy8GsptTRi88xMydvqZ7LP1m1GoWNdmVyNnKou
ZSOyKWf7vodJB7lb6N2IqjGQgtDhMvWODAxhRbwYqbLeUQHjH7lly8MhlQiK3mWA
BEpYvQVHlMvKQJ4FqIl+oMFKzl0oUsrPsUKk/efselwc42khAOFPKj2AuLU0PerA
NoqrxgqW/vWgYduvybXaiEdLtsTRbos7zx3lzMViULHiQKk5jTSzctRd5AUWWOEo
iJ3cL2QXhaSCC0sUOqOhb/+Qd+/xuwH65n2/FiaApqmAqfTSx1riKEv2tPB+27mc
XILlZev6hcz+SRmD8fD3IUKt7zyRG4DwtnhT1Vuqb/ANB0Mh0OFqG6/r2Cdl0sS7
Xu2dllT9g8JOJo5yIz34aDO3dXC3inth1p98Q1Cba4RPfgPOVCWhuj5WxjyBW8bz
hqdx4aneblzhkvxhSufbwZc/kfGtOTj8olj87cnEQCeeCy9atNQklHD3yA+9xLyW
uPg2kdcS4pZ3XPnAgtQ8i5d2wvX/3jzywebYL1tdtKvJJHVpQM32lU6UQlcLAAq/
G01OLGt10iQCR1wFQ2lWjK8MzUQ1AhQA9bIuH5zcAoR6C6N4eWnuK3VqUU2Wq3cc
4EOA7ZbHY+yKIdibopa774IYsc74Lnf6koCc5bWq6Wz1KNZLZUQ4d9q9UU0VkyNx
9+QBg4/FZULwnLgd9iQjaikz00qzWmc/q4CYhvUvT4Ej71tLMdUzPBicFV5lWNm1
+wyKA45yZ71aaeP7DO1dc1o6M8zP9TK8frmsgHNy3STTV8rn64sTIB4R/bcjtoRe
/AnxM12RjPAvieG4oi+S6LsdXtz1AjLS2sx0wgcm6UgJbHFi4eKwyiTszZK0DPro
kwMotxSIr5yFA53Sd0KE4FQXwjpwbyeLUBveb0BDM1bD3EBMjc1xp+XaBJhQ9XD0
du3hUd7tehsbOM5TG5Z83jxSJ+yOc4gEjgWeCbtsggSHnq3oGvRFXiXqjawv8bNb
UyO7PbaHS2kE0TtsAYsdOpWOvkNR+0BVQpQTGwabyGpCg1lEgKvYm3RSM2wiMwZj
AWZUez4anA/ipQn0lCONiEe7iJDA5E2QYjv8jAdbrYwSZy46DgseQ7BU9Luf6s62
K0F0hT1huR8pN0c65GdlFbrxcgV9GaRahpTMQhAihyepSuC6PifmdwN89G0u9QCU
6OssPiezJFrCmgZZY84/daqwes/gpZP9xaZKRQeGnK5fUmtyMaUsWZQeUZeY5hbs
InU0139NTHtMqIyJff3Q9bj0c/GxjcIxaIVfSqvzqbX0m8GGQoCdepvNqv7QRtoE
wTVIofnbYpMQUKSCG/kEgX+MTONslHOXPEtyYjMAPx0YUA0bE+0lWg3jhF/cxKAh
drfGfh/ElV+gB0hTJ2J44zEOdKcXK1Yq61sqyVp0/9VtA4pQUgLBtwTGBnDzsYBU
kav1uNT6a8obR+3YrjXk9QHnUxokn3t2N4VJeiZqDcOPXBocsL6FXuJwQP6nvbaA
8X8FDm/FTBHiBtb8plywjN4c9ei2A33rLvyRlrx2HDOMDrKChY9JO7H4ZGwH/fpA
zq8mmmjH7BKH6XRahlZ2YJeImsPw/CBBSWLUUbg141bLXJBa35eDKzP8jatsIhF+
N/W00h6w/y2LSYXXM9W3kk/XwwKy/HyWuxIDbWp7awAh4D18pNkBNqxv/RWk5/BD
bprQrDoyWPH4XAPKtZI65pxSW3NMIkS6jnBDHHrgRS5WnpIFJlAmc3vZsnnd8NsG
dnh/fBgyuRbhiRxSqLC/mQsyjhyeTuE2Aew/BAMoNisby762nhiv3WL07kkRHFti
l9vCTxkGwxX+6nzsYSauxH7DRgqXCybfyYJeyNo++TnAlIOcquSnUIsuamXP3+JM
/a3GrKL4C6o2ZJ8uGQqWs+LahzNHKcf/ZvZqBs1ukIExFvaY4BGYHc7nzpbtRxmz
+axLkvfoBWlV7T1Ni6RuSjpVnT30Y4icfTvXyp3BNjgRF9Q+fvaS12WUrWpuH/w0
vK7+Ubfj46X9pqndzfYo9JIh3gJgaNqYl9WbatH1+O7V0vReqAJpxy+mN5b2nOkZ
LUQJRqLaQetVWeXvl4QBmKENp2/CN3htkW+hZiRxLtBORdosua8XoPKv0BQxFO1c
oA/j3J4Ljt8/5t92nANML8FyNQt83jpmIsXrSLIZEyLl5cvOxbOb7Kkg7UuG7c6a
QThwzgCCgTrBRojHMHBbapwsB/zzirsIKSa9vk0RW1pHQ5+kPhNAMga0wC4Aprkb
m0hbeOO8XccTY4jhAvstHBuRsfQRYvFs2Bbq9eAR8wuD4MBSJPj0NgdOsyClxsjH
kX6mBZF6b6wmQYCHqY2/zkGmdlkAWZPono2vUcf1RV4i2EO7JOWDIhAyFc3RCpof
0BwBUL9zYU/Ei2Oabd0XaZftGw3hDBCWYHEZDx26Q9zbO8Upk+QmcWtttFbeQtja
nV3/0+XDHExjIJqhTuKG2RttFsIOFkaxzMX0BVNhc7zeCJexTdom5bvswcnqSGMn
MfY+frOIYvas3mtiSLeSOW2vULK3mps1mUDhR1OiW9DzndEo4uCN/ojeUfTvUW4Y
kBeCPhfrGte0XeOMHw1SGU6XXkpKArisrgEdizamG9ADBax6EG8Vpp4fGLbm/89m
ursvS0nvHFWDtH+YkOhB98LqWTvbUx58B6X0YgXV4eK3UJ7HavIgWEnkSjLPB+Y8
0cdd/394R/p4vOe6EuptTHQ5dps0xi+XaROOUPGfOiTEnC6lq+KJj+iEyzY8QCD4
OemVZD4cTeQB13pi3V1cKhhQqLQUYD/oQ4DM9gh2deM/7DTU24XT3A5n2DYKAi6o
sNRfj3r1YelFloWh0HPb1TNld6OMZOb1TgDXVTZFgevJiEvPI475wKnGhR+F9mQU
gDusWhbRKLleGtGu+H7i4QYhuFEsOg8O7lX61IH27KcQjkJZguaVL7Uo7fU7lT6y
q53MljgQS/grn8LSE1kWv8AKXWgziPiravr0X0/ARL1bLDxeceS9CZi6w2pkXufL
JUsbXp4PsbSwrEMMxxYQlHiXTtaLhU75sn8tD/mo9f7dWinzRPFPi/HFsuBm4j5h
5JSOAYDNbowILSXUFx/6popHtXnKc9NdUTOXFXFyM7avTL6K1zUboCg3oij/qlKw
GB2BzimAWprojorqK3MsvY5VlEY3U17owkzGhmh8MdwKPq5TFMW0HQHfuu4DITEt
TCAXtEiKvBmhdN2SEoHNyIXEyhSKar6Z36oDeU/a7cSQVbRUk2T3GLMmTyUefR5o
SSrbUkddxY2B6r+mS8kPIrlRLH3421WNef/IMgx0/cJmPj4dSO1D/ws4tgBgLQqS
LWNvAfHd7UJeBOTLNDki8CNwU25IO7cH5kq8pGpJVAJZN07AkWlWZzAKAL5h42gz
D/Xq8IC2rXLMy+7FA3wXZvuA8UykCVXS/U7SLYkETFhkGfQbqGf090Ne41hBjsOK
gXT7w68/6M42lP/WaK4ZqZi3v0gw9JzDYyT52EO7zMjx8jQT/ty9s04WSMA1AaXE
M/HXQzew3NHxLraQ9byHKxx1DU4U5kGuuQi2b0GS/jNk6o9Hsf3ARN09Hyp3oZNo
zII86t79ZZfgtnG+0c80DjweFolFXa/O+/HL5pEQvHrhDTdzUxtVcB9y1ZsHy9n4
mZDW8hdpdNOCnxTIrcJ3htPhWdsS/z2UfPeuoxYRRnidyklVtFvaicIdF1/yM3fV
UWJAGIVLgrbORKSadkMw6Wp5wpL/80DsnQ2KChnGd1hmMqhqHTySF38JIDpndvw6
gvZ1Dea6z/9OkCqGkA6UGOWS8jYJQje2gqBCQWT1A/cvos6WR620HOvzZN63R6ip
nN3goxZTS+19RKV70epDzVP2RmAPxZPteXTwmY1kYdYp5GfVzGQ0IyctPerl3eDm
X01zby4AysRKuaaoNesDu5fQNBufiBcAJFoC/czmRQFhoE+9CMz2kuSfNiN0DUPS
iH24n30OYMKEb3bEbdoJSbT4KEmIk9lMJjRjPO59JvvfFHsBgZLSrYadX9Z8lVuh
lkTMHmhPtk9FeV1w7TxPdrnSLtM1ZSbu0f6E+4Bp74U9f6GEOasd0QUooVf+GL9b
fsEvfhDHdiiEQTaLsxh/5qKzP/crrE4gv7DfLho0LN4S8Ky4hMKwvIOA1+IvJaX3
lQxk/tNbf2EeU6Xk82G3yDvlB7Kv+zor1K/KeGEZUJo2SuvIOQd8bCH6s8XsOLcT
lFagemLGk0ALGZcpm7fZmmCKGnR/yqu//rMv1xTetE6XbdsElpzjRE91jJrVoKas
67NRlwz4PSAZ2e2HTuwwPNzQQ4fxuZZLoSJah3xismRepw/8ZhdakNLC0EtNFlmX
0UL8DN1VlNRh90uYFcMP021sJacUqTEVveiic4BqjnWVtIiW5j9vOGAXTX3EtiNq
8VrvG9d2ATWvVcxg4zCQ8A8CMge8QzD96IeO8i1jImIYxN1zc5xkcPUhckdwi/hV
1l+6wjBkZYz9Kn8wCQt/DX6lKW3BH7TBJyLE1GqVoQvJj75H/GnjkQlVI2RDivHS
dn5+CSZGA2QAK5QXOlWJ/BJoa+zLPeZsR7EqZ9vS0LB2BRc9aIHRdQKQk3dLb2K8
ceJc3giO/ChnYxhShZ+tsZPxwTuOi5Uoq3GQXUXjbB8dV/8alR/4MZMy2XtOplnV
g/4sOsAcsEBgxOLSax7kJo59b67fF5vzuXF2LBJeLGl7frarMY7keI/0KE4TRbPI
FppStOl6rK58G45IH8jqiQpLVYf2ycpJH27mdDLnomJudflZZTaXMlnNL1DJlkY7
L/bv6vs/Ny4HBud1DPcYTC0fRVxMANPcIFmgmIUtjcSzF/3dTM1nXRi6rouFTUsr
6taRW9gb1LzAwJXn2eRn6E7c55OfAFWApjC8rVwnlFs7Es0MyhZydX1eUs0CjV2Y
7+P3s9ypFs9Oi/JPkDDIteYIQlrdIXGw+QbeQs4PlZnots6pa4VGO9uTVZ+x/ACY
imilQb5ZUXR85YWqIqEXC91XuS65EkmMsMriHPmrEv3He2DoAx2RbkEVIwnECido
D50nuhlk2w4y1YRJpsDV7CbFkPxjlEuFMTLdn4o16wCJKaqF8SyR7OhVkTv0suAj
VemfgynH6XQFGwoIx8Y7upIu5fbNPxX5b55ePswvWPaDniTHGJXFfIF4HW7UmmcE
QeCpG/zA8GFizvB0l+LCKp4sXZA7ZrzeqWDIhHD3wopx8DoNvLmApsm5F7RObuIA
wy3FJN4XzT8uFRrSbyPevY0AuKo0lVWMIJEzA7+GXCY0CMYQnBU2aZlYNytKbtqk
IK0Sr5q2mjwbpCIQtRH8/wXx9meDG4Ea2iwutfiCXrThCnkuIfhR/WzbLk+Qgkd7
HZklq0jScpeqkZ+h5RIBv/bTAjNIduUszaSW9DkPNt8+gYF9gueuFcOYF0XKbwtk
v/u0xq5j6y47fZlom8GgUtqQ5/7ibnn57EBmr340HCjBqBBZhBM8sO4A/mIPire+
cd0/wTE6k3rxySrv9SFLUWlK1yG60xPECOx0DffxcSfnPUmwFKWpDEF79U0imZ1k
XkF79fs6sr0l3I5XS2kW5M9qbndRPZN+lLsZu1es7W9AulaqE3g2Z5+y5FsD6kGl
wtJUYvv2n/8a1kMKIdaG0EoRud0E9I/s6BAzSTD9BOLbyZ5ycosEXCF8QUqYfkK8
0LeY/uW6KAuZFfzNJKerYL9qIEK95GQQOqbJzklh3ywZpglB6z/akexlNCyNgHAJ
ER/IB5E90/0pwCN+tK1lQeJI2i56vtd8QBpOf/9LFaynHEz5ToN8jWFGuIk5oeST
sNIAM0QNy0RrS/p8+jQV01QTnLQShH84Q8Lq3p/FA5I2d5LrR1OxO1hm9j9XTEla
I+e3oTrZYA6CcjPItoKW/8U0e6QudQ4U9yyXmqDDuuynOwdrwlxJFSDDJevFpScG
QaRLPm2dhInuv2ozuqN2xS4/wYSuSb/XCARsBh2b5fnBaYZACSfnUtCwvhhOn4R+
Sqf8hbJ88sseA3+XVTMlMujxXjk8CuvqXrsaJKhjIPVqky5Aw16FbsVtkW+PEXFt
j0kxi7PJJifuqKvWL0E5xmFYpSeigRYsY4nVMBtRdAGZNF2xzYga4QfuHzyfRUSh
cPNn2PtDoMMPRJb8K41bg2CEf7bXqLOfQsdoD4wYHZ1ycpzzdPpQahomTM3yBUKa
j2t1Yj6MwC8abGBuPBq23BOQenWYLLY+j8LDuf4DwCU2bhQo5+uqSE6Qacvkyz9D
NSo0rnGobXTZRLeSXBENp1O17OQchjF/dQ9YEoJgp+kHLv4tiuJILv2JFgoFppjQ
1vTdmq4g7B5TkKyxYm9YDcXhzquKD8SDSKvuC7Pb54CVqMPyZXQbM58bKwdmn1mi
iL+ysRQsQNnQzKj2ktCa+cVNXgF01Z4mMIMdmQEQEvh2rLEKm1we+8tzWq+JwOnI
IoP09SjpjbMI4vlQU9O0nlyCCzWI9/mEVbF3/BGeGntyPgdwLJHic1bi2BtLUMzD
BicF7qmCWlOzoYVtv9eisv5c0UJFRi6yanx4wBatAGm+EAR4nixAHhDlyKtwhE6Y
QAX9o6rqoa1Q95Rnk7MQk1sblWWbJR+vO/jVK7p50IxbW11PYxXGTdPoIgdpLL3y
QILuMdVhUcCgohdQHLGhfrITxW4VprDQ4ZUC6nxKeJJ2yDVIk8wB0qVAumw2rtB/
6cMo8laO02S5eIeJ4Tpbo8XWbtCU1JxHsB1FcwupWMGBtiZQok8uKBAxItl9fpwE
cTimfPgdYWFivFOkatQu98jLnnxaP4dJO2Ls/l/5lS4ggdjQEsZ2r3Mqxnwmbz7T
yCpM//o/snpJhGXNz8r/6Y2eZw3NGUAwXDPO6XHW3p45EL/u8iFM6enZmVxGETl0
Gqm6mX53ya24ikSPKffPPHqleGr0m2RMWf8oi+XKnjjq6n+S6m5hD6lpsPdywuYS
A4k3PI/QOZBPkS5KmJ76uZiQ4w3jzwxGUhZFTW79ETk9/a+NLUQggbWmz49vqPsC
/Kx//XNYf2mvGZJwxiMWx0OIhXEAoOVW5LrY4+ZqvSbPulpGNqxLX61S9md9+ZGd
VbLOqqE3KREgwyw+/TCsjOIlNoYQ0Keo9lU7mmF6pm47BCvwkZGViv8Li51SRVum
H4QA2h4Uo5kow83+C8SconPAIypfUzFLwREoP7Izdu0HB+Do18nWikzaR47bdRvz
swlCx7f85k+wqE3qHRML5WlzCl0MajLVPve8uf9cCCfB94ykhrly0WnFnq26dDzg
Yt8YnG1vC0SJPUNQVHfh7c0/KUC516P7IoevdzjhQJmBn5l1NN1nMO0O5ZN3rCc1
r3uLgJPFUYASlXdwTzdN4pI1C74k5g+/FaxC8bXiRNMFHXkqibLZUxy40k2bDHt1
KV2c/y018mDh7D3wkeg7YhudIGbVx7Fqqs/fmowxnj985pQlqBz3EMW69qp5MYwS
UsVXzVMjBppo4PBUynZk+6PIfV53q/7c5iVNmmanJAb4vUAv80XNml6zI/90D3kL
zjJ/DQsLZ5D85LWTsFO5abIqiDb+c9N4iEZLHUXWoaAys5Uq6ktTFqNDwiSfhGmi
MxuOYRouZxZe7GqDUU0heTZUEaJSncCX+k5AfUtdWai0eduFDLkMTiacpkkO+4fS
dq2xtUvRxwBH+BU2Zf4c82B+ZAuPWpXrj8HuwVV0xWvFarRALqtkQlJHCaZm/j/R
hRRhhpcw34pftItHrE0BjRgPiUdEmmlejsLgn0nO4Z8Be6KDvfWBnmWK6H0SJMOo
H4sE/EvsiUQrj69DQVycZUCBOGuGDiegcOi8eb0aQrSBjdkEFQhnVlYvfkJgItrg
GZf3g0jHE5NMHm7J7W888wKvL2DJWKGjfzCjUW1VQiquvZNr8UZdJxEWKhq6ZRBD
ROFNeIlr4/lszMn5AUQ9gqorgQuR2C6oGu2CGY2Wi9Fjif2KdYSm1Ki0Tmjq8WkV
z5jA1rqd5NJDyacRirENSg7br6xMzg0FXckLBXZygnc74lgT0MxEqAbcj8FBzHR7
uxEoBNAb1YGEcnVJuJRiY4pxySGKvQMJvZ7IoG0oL/AeT1szxNywGKH5hYgbzqc7
JsjdsmzCtOGXdN1PrjFKvjJegdmGaB0YjAGasLBaXEXbStcxKq01pBRVM3vsroL7
GlSEvItI+UUuOgBsXZ2VsSKJXNl5xS7LptVNMEQJv5+P5atycAJ/3EXqKfKlwgx0
VcZB4TE8H+0+O3UhE5lBTgPA7W/pUkSTf46QKjOshkYIuwc3n3jt3JhRE4lsSMaV
BAEU3dahan7SynnziA2eyXllqWktI/MDSp+TdGNrloi4+VuNykPuPjN2wVAcwtJY
WkbjAHQu6NdYqfyRZWIlGdDonB5V0mCCQXmYOJnKCwaHEqS6QWdBwxbBX+ME5MXI
c9vIn5FNVJvGt5CiRtTCGQ+gwqOAZ9/AC8eXJkST9Rq1b37M4t7jUPuSbOTRtpxc
N+ZcdemYXisBnkHkXvvEh5mJCYkwWHNp9k8ykPA9RcjqvMosAze7P50gU0V8tEtA
jjK9ov3alWOjD0fjo1AfEE87ydkHx5uKhLUMSEVhsx6Hb6qFvDCbq980W4zV9o2E
9Qrxhsj1vswJUku0bvZI/JE/nt6YyJBDrJPjjxo5PI6lOg3SPJ2doPA86hekFhkR
vcDqv6UHIIP7TgE/JNSQ6odpDAMXDLnZvq1MglxA3fdMpJ9AorcqXuUcFKng3nEE
12y64JERAE6LJMYAtqBQB7IAjbbhoRCSaIzOYYw3G1dXQ3N3ADTHeMxmj7DMtDFL
0arzw1eg1p1+48XsrfuqPXYgVC0lVk2Lcw7c4+EQzEaGFd30WUHQ/UB4xPHoHo+I
Ta58YtDvj4ZNIdfeNWiDjyqlKd4Oq5XgjDtGj1BIotzdJl+9LET6rk46W9/kWDzj
lXlsZ0iQ+pTcJAvZveQ9tKDIz+S1Pvp88akhac14Rd6lRSUTSu/JSAt12vM/1jvD
AqZWPUUoQ23nkojx3Xu4vVrb+SKDV7mFY42I2ituA7P/t7s8ayaSPGo6DSbRmToi
GLF7y8hJvASQUKhT9RnTXBTwnKhqXhDTL0YxBCZN1+cD8dgIQl62HIPyFYfst8uz
DAUim3K2cmGwkwo/kdpuV0QIFXSJO5cnFORVTm7oYZViSZ/ZYoe4OTwP8rgKmdDb
NX4oXfAENOt4gCKq8SGrSWmNrQXINzBRBFtX2IrDDeRvwIvC3EgbX9ksZjua6Tv6
Rh5mcQvWtRLXbLAMUcdCgYaamXX2wotf4Q+rf8GM25grhqirGtfLldLSEiKW9D1Z
Q+2jwdTQ3GnO9RM5iF/LlUnZwhcgRprZoCQHnIFuj0cFfM+DKrZg17oVZ8U94LEU
7l2BY6FcGTQ8Sy9/NlE3A+KOBabvun1afJLaooNZSrs+JsGR4pmsW1KgaxgGpC86
sx/MtD8REGjyy7/qErlgnQ0F9XB8LkFnBxiSIMD8U0HdeenApfVscM7BDjI+z7+E
CtZJo7xHmdRMxSxS190DeQfGG0LfcSeigLGsTLFyc1XEt82wiZIoOcBZC2tgINp7
oI3fhNasV4bpsHWbnR502Y3p0bEsN1c07YF9IH80ofwoEGvoRF9m555j1DiP/Na+
/bWHi5qiH3SJd6YIBebOAPRIU5yYigjQ09wkOSy3wwi1WKFoBYeHl3X/iMKeKH31
B6VKP3rmibZJMx1UwnefNla2cw/037tYPZ21R9vhrikw34KsrBTJdHLJwwxNnDsL
6dnxA1HziOZOqKTgcUPcFTM2/Np269ysnOJf2uKPU2GHqbIYWhCycxviS22KVoHs
NUuTQOetV4FaFt1tpBCrvyKEu7vvhh5nWHIzw1Entkyq5tClS6Ik5RrXaS2LFKtn
B3SffviHYmrO9vQE4NpYqwiHbwHN+L4HfQofJevvvBUGGWfyIL/ctCqmoArYT285
8fAPk0K3F0/ZjxTxJ74qxoBT7gP+HYqDoiCyz6/tH1s2QGLJ+xqFKOXWJnFtzU9u
cgV4baFnZr7ElDBuCYT9F8Evb3jaqltKI1AObDURqP1Gtr+DjC4q0Jm+YSHOnOy6
SIS+ggEc1c82PvBvzm8vFwr7nwB6zuyE0Sudu+tCtlWC9ksf7hxGamF+YUNdI5PG
dS8MFqyk33efXAvSdPxMxJ34z4dw6b81wsC+QtP+f6HZiX7B66hCsRuP6Zm5izPi
TG3ZFGBiAlca0yPiY4RFftYLlIbkCGk1hNUXFWfTjhM3SqzrKCNV6k/MOEF7e+He
iMdbRR6KMOL0DEeOSSjKWc/093IQEWQ6Ln+oIfvIJHFzw7iJ9YPdRApyz2SVIg2r
xqgaKRSkUT0KGJ9DV0s9Fi53ZEaGbhL4HXt54XvlY+xgQRuVePyI6wsPkFRY8gG6
mgOT4bpRNRM+roCimwJAMsnq0/Y9ffa3dbfWCbNzXC8mIpCy4X+Q345PYKiNBzVq
omtrEewFBDvqD8uHlx4EfLesQsgt8SfILVX/iggBYqh6100YNlSSbQ2X6/JlnaD0
8xE/NIu66GOM6eQHKt1Sc0+gh2AONKz1/liWjbkY8V7hNK4aq8os6pG0Gg51CBTs
2RSnsznFf1enZtmeQcnI2hOtv23wZzir6phHCy7fiOTJ00XKZBMpJQrGXlu7k+0T
KIFBA29ydvyMBVK/0DqmQxFPetwNqPXtAWw27ZqcF9row2epVY1kUISzvaCwR0oL
Ga7tz1LXYUNkiBz1eMAVFng4i88P96m0THQ1lXXmI7wFOKfme98y3VIvWRMcuSkw
EP9TLzDFY8iCuq0f+vWI0h3A1AY3+Lk0w9mBqBk4Z44nNYxzQAJlmBhBzylBT3Uu
WSlL8DYrgfPatz1mioLJo8zzoU+l539UiC4+fc4LqD1uzV58rmmPgHPM89uJ13En
qAo8d2e8fr20xPMPHzCd0vxNVFpmNeZCZ18cROn8/8eg6ZyAbbMdeBgwHD3VYjzB
xpyZNksMFguMQa+TWJALVK+Y5h0r/jYexyvcSveYhrWnDUUZLP12KxYK3feTwi4o
RwTF+HDo1aXBknh6yZgO9zTbaIqZ6iIDZ4kbXTzzwFRoV8yq1zQZZeuc02WyTL+V
zTlDC7b0LNAp+8UnDt/wi59Y3TaGf8URUNkqpQhRuSm1vppeGbY7sDrt6reYVOK+
2xVAgAwdTD0KrO7i0cuIagCdmj3/jdHS+m+Pssjn2OG525IPgW6niJD2gT0Z0krL
wmHVGWATUhnIs/Sra9wxhyt21P7DSik7M/HltYrZgWk=
`pragma protect end_protected
