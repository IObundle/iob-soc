// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:00 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qV0kaU9f2imvyNqBJuGA2qC+2JDx9WRufqaaEOXfm1W86RWESY6as39lh4/14zqP
uI9QR+1A0lOnCkiC7KfKzrwD+ldKdEikU/vDuZ4kSlj8x55x+PAt8Qs8lJrhvKqI
BDoEJHoKSvjGvLTP1SMXyLs/bTJ2n48oeeS+SxRiRIM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42480)
mlz0fGkDQhXEj2vTjQw+cdYTfZ6XqBqWinKUtR3yTwuakbMUB1K8k8X6UB4q+/7c
tgOrVBHiXxYeX0hkm7DErYreCDUi5eNKVdUpePMZS/j5+1zOFHwcISdXd8sXvc0G
VKIretTR1PUEOWhHgTi8pmXVa/K041vN9KUF2/RGxMLRHQbwSOMjS54CKwh/Q8lb
bFvBmaA0+CVHPZ9RJIVDebdgFS/jY6urVaf+AOFvops4rEdpZ14yfteysywHmOBW
/WavDLcllhnkjXdKWRNxgGCtQuREtCG7GKfNhwj3kK9Ut/ioBNhchkvC09RPXJFe
+VLKDG0P7+4J+uS9uEHHsvp/7FimCxUSDsG1YtkMUAsaR1iBzXMjiB+qGQwMdOdZ
FnQi4eQYb63P7XHUAT4UzNtcvrjQzGWUNbRYIbQGgnjqjWcAy3aLe7K7fqMiM8D1
hrHGyJ6pq3/n8P0yyE7Vlx3wdUEo5EJNJxdLk8JgyQnUbwdGkUrnRYECRvCUkGeD
VLazAQ38alo+6BSpfnUWTD2xNCHk4V9mgYYmcwLhzchnF3aTkb43ccy6yvM8Fag/
Vwcm5CuTNniF2mIYKgc8jAE6wisY40EPcdLZczqyUuhGD8w5cZNhVRaq5W9D2Bek
xAFfTmzzSMrNFLkAO01rXOjr+q9AI4MpfMkoe7eepf2Xf+5YbpEhMj/SWQQcGmvM
hrPnO4v64wHiWOwkDZe258Uv2e1h2ApRPiDQbZ2vBFeNsmyu4wysVp90WH//x6LD
aK599yI2hwLcuDMpFqOHM0MQ6RFqoiLFoCLco47w9KUuf+GLtNCmVjnFaIs+P2ul
H2io6immste3O5Wo7nEZ1YgjmMLgEldV/4nVvTuYEtEH31+bgmbkK55uqLNjuh5O
fWSr10HvOYhppOUaatpFHwSrQisZ7BBb5mpClH2sNgAfJlHMHiUzA2glphv7RQlW
bRAHrNY+VS04j5FN/iIFNWX6sgRmUABerNkg/gpfJwmVflTvmAbiWuamf4j3qetR
+kSPF9R1rUosf0DeVltEzuZsLf8TCwhXXZGRPglFr2aff5IqMxnLqatocSy69kVe
Pf52sXxD37p8jZEK3+G/RB00pAWaTo2mTEr3sfUguBkRKNEkgnHVh72dqXNhSMh8
qGC6hdR216/lGALgwSWPJpeFKfXpLgQ7J1XucEy24lnBmnUSt7XpAEJMcN0LmfMV
jO3fnXLwyXYOkJYDjp33wxRuYcdhTRIwBZTfiinnTsnivwUFYqKtUVEriHJlkr9o
HeUsk+sdXCFJVS1NfzGSQiPkYuThU369AL+Att3qhYzDfeBS+qrNJCIOySYiaf2v
U/HUqhIGEUhR4tYFMXOtqiJpZuz6iILe5lIULFUjEhGn32xPRLTgRUZ12Kb6QwbV
2E8g3nPwFQr3P1BREkPabQXGrnZIuWF5ad0+2nWknPguc4dxdpni65nGVKTLwv12
zWf4BE2PzlFGMpxc2FhXSsbg/xq1KVxGnL3BJbTy0UveEd6IZ80p3FM26Y7A6fZs
jDsSgXgYo0DghXVy62r161skchs5H3KGKdIUnPHVhrj96Vsme49jawhVxW/Tc7qp
zxHh4ZNRNyF+NtpUvbcN3kh1UVyyqOrvMI+sMUqbIop97cADWaZKv7VIued81wWd
Dz00SOGJbTTrgOZoS60ZL8qkTuXWA96dZeJlfQOvxjcgSurL8eONgGIyvGIxkKIL
qgy9aKwyQWuF+YhuVazELbiocKIcAVO2mYCPn6FbMiRusHptfXapJk5NAQm5FiFP
OsMYD6iyZUwrCeex0pcTfTXS8TYRoZo6ZCtgXpLxqsOplRqeRzm278qCT/i9BDiz
CKaiMCyLfloe5hLmuJyB3bHRi53rGwbAlYfogOOwP3LcbgORx7+hAy6Nbft5d9QA
J2ZigAzFNM+NFcPAdRui9UMdQRxiLdGOANXEQQE7lWbWhpYXl7Tq2UKD4EkTNl2f
dJAfJmDXq2+kEZB/FlukAxHQ+qGUoywdkjm6pQJgpA6kXVljLwAWBFOeiI8XEjw5
gbmBER1YAQd2Xzj7EXI9yBd6A1LLCrRMc7bU6Yxilekgr9WbezDrXJ/TWs/CH7JW
OUSVC1UvaGt2/t3dwh5xn30QngVK2jl0V6+l1w3WmClWlg+UX5PMpvuxzZl2Ul2P
t5Xu/RteEqkN8VLqh+aijhNvStQX0Y4u3e4B8Rm2hTOiZ0L30B9iOPBjLXtK4BpF
gkZvnqdpdkU2k3EDrNF28bZDgkyHBHgf1c7nNBZxQfVbalzX9jib3/LAZkQLQ5RP
Namru/x8yQCV4mOj/pJ4+7NS/dSvKJneDxGo94Kf2hIlXKyzGeDETRiVz0Y87KF+
b/jBPdtij+X6TL4UzUu0iCAhyiS/BoXxsFDavYJFE/eM/TLTq2+x+/zvfjaiBPH3
PuMzoUeNrCm8M7Wopq1sT2/a9D3J3iGwZ247PZiaPEbzjYinESOlD2KoCxxRX23G
QS0umQehd8PNzUXg+vYuTADG2+uX0N5DJQT0JE2X/0524s2AyMiEsQXBNkxE4uEp
thwjy74BJOvbF3RO+BoK0BxvGdTL/QIJCuI4ByBxi5fZt8FYZXNLE8JiYvaAcqKN
ykdE35o/P0hPVJfl5yKqsmOaHzAeKPE5oqqHqEIoXIROO8mbWeN0Y1Pn/JbVm20z
7Jwl1sr3DA46/UY1VMODjOVrDF9dXkHYpBsz5pFSlyvijICPv9JFWTt2q/YNwdRt
vCmNdydK1lvEz+ETgSqKKw549sFC70vvVtnCeDWCxt6bCfGBf6HjKov6kPEvGi7s
dCW/KxR5YdHouAnZZbMECnWGXhgLIiSYMQNmhH/cXzp/mVAqdgGvDWYFLHmnIGk+
5r0NObuDhxYf07CZi/DN6DOSavdFSvBEYOQ/f90LD8QcoohNCF0UfZuw+yt0HZti
FaNHpiobegDMf+Tzd3EIY/ucDP8jffn4x/HTGmybqlofaGtci++3Z1cvwqjJDpGD
Y1u925NB5WkQ68wH5Y99Pth7eS47FcnIidy9Qwy2V+/rINLuHtUdOaiW9FG0vGvD
aAMYPmU+NejBcF29EM+Ycel7InOuPJEMF3KNfzTcF3AQk51wbquMfql86uJcbl4m
Octo3YZt74elfbLj5k5iPeIKHRVvy8uNxM7KWotaRAGZL2y0W7D+QFjxyZw0UvwP
ycikMdcy7az+TSwFjttLDe31p77o0xsvvuzLdcneCM+Kp/s7YGmNjfGrFu9np7bJ
YaLBKIQgBKcMwouUJlL/P7i5OUOKxAIH3zmabVFbVdQPPYXcI2FqGGlg5cHf6JCd
AYcmcu01aHxScFo4pOXH7TAXtt6LWv0ncJ4rpWjFGGku7guSjOgsgkbo5skcHo2u
U7CQ5HBTbUkclGJbWjNMfeDUdRdDi8c82en4jVdib4KhU5jZbVG44+anSjfTFGFj
1R5S9d9A3PiVcWunc/bac6XZC9tu4uMevi/OAjzTkXnkSXhWmb5Y4tS/09lwRZIZ
XYiZMdO6jZC5++e4AaYkqFrMrKtyfr5V6Xr5MckDjVN6jWIJRVcl8pxmpiQnr2oI
blmYEB0GJgLh2S8UeNL3uJjdr4jX6+rFG7d6WJ68/q87fOKASvrpzC/mChXEn6SE
fTDquNLr49J9zs2LO8BHcYBnFeBPftyGS5IntfDDkRsC1VeQ8QU+pO5aL7WD/u5H
jKc5Ck8ZDdCtzHpwex1i80GnB3F0MbQWQfqip3E2Sr4O7Afls992VRYIkLy7m2W1
QgfZM+abPas4NuS4BmpKFUxR0rRQROyiVESogH052IT6qifG3Ot944nzBq+ethbW
s4fA/m5j3wKubWPdgupjovnX0hxCByde5Mr8eHvvVx1W8+1jFIze0duRIMN9TqsP
dkuEQn/+MV95M1nWAr2myZpKhqSCEbhurqIJ7TDn5SAQZcSzxy7jWn9l5xA35ch5
zCly41qISAimYTZ7c1HUGQrnFhWtlY9DzozpX+gmq9DkYaV780ItSwLcHpS+FSez
kU3f3hEohjX0Dxn9qQgcz4xHPBn0dKPM6OGvaeLAFNB6zH77n/BsRQoVLcKcBXca
egVgEFAQ+HASSgwV3hWHhE4rREKTWshe3omfNNp+tSjDF7IQcch5OM2drpu82QGX
UgNNwBv9oOOciwT4v/Tvth4tA8K3zUrO18DmmFglek+27LzncbQzZFc7WrY5iABH
lVIgECD/oiN1rAEXAq0wlhXK6BRw1yiQFayNmWTTO/g0eQwbqKdP8pMk5flxJMbk
byBITsBFR+ioPEaEKi9zWqqL0+4pa7ekBazSL3SAnSjOCCOf6j3HN+Ay+saQc1AW
djayqZOFgzxVCsGE+RfWC3yTu3xgEFUDjnrpMhwSFecEudMHHVGMRM6/M0LDNiuo
iRhAqbqyy/guwfJejaC37BBlvWZUBcyt1toGnGeBBdqTG4s2ktylULDA8YHvDOFX
HT9xg8qQFlScHrwPvs9L3L/UbEGKATgmCNd5giADRrsaPfnNAAzIC7tl2REBTBEx
o1JK9BZdaavUpn8cxjk1gagY13buyxw/w0SRwnoUAwBIqmA0nypFJWv3n/EsFCv3
tkAOZgSOWBPKLk2MjPBt3g5xS7Arvol+xf+xXGJXegjNODCJKLrduMXzaJIAVReJ
gSU5LQWfDoP9EKeIjPxiQXtTyW+mZOWr4vfDhB8HuqQs/PxhCglkaVsupYEdPoVR
4576UnXa3GLmWisUS53hRJDEFVLqSynrsYukGXuTh2GvoMwcgMVC5ay7qdHyN2zS
MBvXy6xgO/e8MDssbOi7YE0IliiNhBeboTCZjQizIDnB3SFcgvQcKwUDywmqUcUT
91pcxHlG7Z3XU/OhNdJVVPagzQnvBkE4bVCHQTCg4Fc9jjnpKpf2njzN8uC+lZIz
8pS7u44ymZ8gxis+0deb9XDkMOkoXUFtDJKIU0+jXPwDNzTvMTpjfBK1RiiOhQPd
0bYw9DRim8Q41DwxcpQddHDBnHGrUP3WOshfhqP/VHu8AKgOJmFhw659yuNLPYIW
1PrHVGOt9WwY0+ivq1rB9IYcOnTPQRjlxBXvjaNuyyCzd73lL+hXq326oWZHpCx0
tySPBRFmwHUJcGoswEbEkDtliX2t2YEjmHsYGwV+hMHbKRXSdxclPan0UYto9wFI
I4RL/hZSkiDxIivom0VzO+alPR7mlBm1Krwhs8HauK1+yRpfjW0N5x0Saw8oUcay
Exy0QM+mNdyGVNoA2u/kChQ5PcUqnVRa1JX3FayUwDkrFa7GCDAHp8r5SHziYnpF
QB/X3ESAC8n5A+yzn2o2KkEthll+wQRYPEu8UL5DAQl/U2Xzy4Lxefuu/M6mDJ6i
YRT918hulQ7OlV6AsRBR8980hKVxpfdpAeXIC+OxZFZhF8qyptoPkA7SDFYZkovQ
PL6Y4f1LV6BxxtomEfbPY/HR3rxNYgJxu4LO/vcOVkEMggX523liXpYayHaof8sU
U9GYjQGsoy1DDRZ17HoQR7vvc2mo4ZjZYDEK4IPy/Vty4cX1uqd9mGHwFFmxs+V3
QSvxi5URpyGysMCgYvYVHCTYs2P+7FDYzCn1om/DaYiWAp6hJDUBD3XgYMUIUPwQ
v6AaQb27T32WgfKpAKi+MPnXiyTrpc0VnrLI+zPfMqUgcBgYvQzk87fvjSddc7o/
cs23uLR2ZxJ+mbW4LKdjcIJZdUPTJfpQz1ysKyqEc5PlhfkSAgISNFdaykLSmW4o
hcqUVreI/O2WpmvqaMpV4DMx/A+RvkwAsVYkjnjBLQC6HQLpZY0N23+Z7I4rlLQq
l75z1AYWV7Ii83Yu5TQIwCp4jqHXeZzeebMITjUKSfvNR9F6mWk98fNAG4CxsZEW
F1Wdpczr9oIA4T9kHtj/is4TsHb215i2pbuqktXeJWV59kN7g0QxoHMyLT8bc44E
/buq8sMnwNpl4FddyA10X15TY49iRYyRIonVMfQst2Nn2huBOAg6UtOf3w88GMZ7
VjvaWYcKJsyQOlsViVa+tXyroHDm+al0Rz0hn7VCWOmr57uPuCgYCjcClAC4Zevv
e8m3MLJZZR3hPgA50tKyCyRSPF9u8J2Rqo/GPtsFSMZs4qHSlnijjf8hY62xzfcb
zmdZJY/XhSILItXAbelnmdwVeALy2ivcthdCTD++1NelFgBq3yUx2JAay3fATX/L
C7Apse/jspeDj5XTdQtAT0DZ+Q7kHwD8a28cylKrH0SuZXEtpzO7Kg1pE32GKZbV
G7kDzv5ij75utcmrSqLoZe6jQMU3irGNNH+skmQI9J8bHRPO0KXYYueg3GBgjwQs
1MPq7cJLPxsf3iiR3PduP57OCob/OZBR1XzI7PtRtqq/iHxG1IhHhKF0BgTvaAx5
vkHWet6XnefLK3UkkMgh/aJs119Z5sNLbvcNV1PIlj1+rXQbMxIU07qd1IUZoEmF
I9x8el5RfQTXX4N1o/RwQ1tWLMBa6uEHeUGWn07FTcxQgPVNgn8wrpr24VJPjhmP
qod/TjHByQqpEZxg6tYpuAkTFX+H6FziwwtCWv+KlQ4o/ybXM1hJoF4Lzv06HHMM
YRULF4b8gGAjMbuzBOvE2hj7GpRQkYqgOV+zFT1OIcJYPmjrYZ2sjoPXq9vq7zQ2
uaLI8rVOLBoeQ103NAcadNjjVMcWzO8gBCkNOMdXrPdr7QSjus36s+vRFzDdPcs4
eCZgChJAGgGV0HITQAQrxFBZCymIMhYiBWe4elaF3LkNnNa6j4Canl4j49d7Bhlp
SKOGt0xDb7gE9Zy7iRGz0Lhx3QL2pz5CWAvUtd6nptXe//O7foL+mmqG+poFMAjm
pSSDVQ0HW8shKmZGFCnXmRbcFdVWG62Q/gP/P7/ppJ1TFYtjlFQq68JtMPnriFMY
zd6dWtdZuQf3uMLQgijMsI65jLJVp5QFY6s3nKSow7OG00BHDVB0U0a2aInaLi+1
fKC7YvbndM6X/cXDQBmCA18S2zodZkL958ugjeXljJ2bvKTvMwmzgtdJ4hit0kWR
ZhDLsahOUnuDNK57BYlLCtWCLB1/wwzeSELutDjwvbuq9DwJmSdYwIqneLf3DwNf
O5G3c9EghyAoZvIIdu4mvo4wa6FraVtQbqnSPTT1MNjJWn9raLRhwG3TXqLavX75
2LUvXxnvNKrYSDyyUThYIpLPHZwb5twTFHTjDLk4+YQuqdSjjX6Hvj7ILRyV65Gq
QOROQyUnEC4MPruYhi5KcG4AYTP1cJKoQrtXxeSiWYzZLSBdEbH+yxmBSkOQh1LP
CEDAvUY5qjOSR4OcmXgJ/kR8hSQYW7agNBRrGjy7gt9NG3ZDZWEq3kvnLDyqkcNe
/8tJFotAr8zCWa870fvhSiDBi68767WJRJF/kJda/ftJJVdP9hQxXmG7tgBCRkAX
c7xWAatvb7kU5SjakhzDlhEn0UTwbq52pKwsAOnLesW+MNwMdMyygCCw1bbPaQwM
cnoob+UWFwmsQ61e1xWbxA5wWNDatAo58qrmdtvJJQa7q+CfbJdZH3qzHl7QtKxG
WcYz2z2ZiSASIqAYHbcTyoUGhOcSPK9iLHEiUrka+gV/cv+nlViIeW0MA1KfmgnB
oRzz6e3xRHq4JxADPWai46kARWLsGfKwkFU2FU/xcIlMLCXKVHn7ZZ3d3fnBJXB9
c6wxvKJNTzuQvFXFrHeewD3dk5eEIs+3iTkDPLfLKMmz+02xu7uTqbOE6lFoTOdg
V3+nmmX9pDXGgkPr8TmJ/79ORajmyCOyfRXqKs+hO4jwsAOhCZxTM2pDzyCoym1S
oUKZDTEy/PS9ezUeSXYrIIgAv4mNZk0ZahgUoJVQj6RO8jMNGyGor8/RhCmdKqgU
ixXoztnSgHfgEU4UF7uIJxAxaHVzrFsKNUZoZytnAo4HEgnbYz0hnej+7FEdKkqj
GyZP0QEaO0kJv+d0uPyBcQrujpKA0JHbf2nWVMo43DGQmDapWnfsxwJJcSCVfYRZ
tSfm5z+6gasEsgAg2AG5Spn14UafOZxWVoc1eH5o70Z+tYg/d3QDRt9ZprsxBXCg
6S2pgwO9BeCPzBGlGhYE5jJHF6HaHCB6r1sfPxJQsvS1oofm3ffy+wmv8TA3B3Jc
Qs3gx8xxeyGW9VKpOC57g6LUEOK9A2VjBzxhit8x+iLj/zjENWuTqLoz3M61Oz6O
J9ZyifYy+7cCucnKnRFSXaX6lD93Hf7sE0ytb0hfjJbUoAhEit5yVRCuxH8nLeY3
qJMJljBwA+K9uGzcg8nnj9Il5WPZ99jnG7zrehYhrP8OLULuiZ+d1gBGHyEfcXrw
1qLkU/2U7S41EeIzuXYwMgeAWvQFibg5Ut7qNVq+E8cD+IbYSBPV7AaLKNc+Zf5s
pCYxEjoxuPI8Hq73WLWHcFPHzd9njT1vgqF/mbNwx9SuNn0xP37tFW5nuMMp9Wtk
mu9URgZew0f+HwqWH2EUwcc0e/EVtOyGVGmsNa8X74UTK2st16vBdJx1myq6+PKW
ktbnsxudRV2d2J/loevfCUNqNHHhYWXy7fxoG4+OUx3blu6U6AmiRpdIaRBzsKaK
TDbrAOQRGGX+XWpbain131wOWm9lmkaYjXbKYlOIlnFsVPM+y85ciIh+diamk563
W3Cn8a5VVvdYpM9zVjBSeWkdzwUtWtt+BjVuEunT+3Og45qLO/NCO8h0y8Gv/KM+
A8shqtjS7P/WiD7pMc3WbEJETTn3CSsPMw98lLbpcohQswXGE8iqnOcFvQSRc4l/
aY6XUoYm2kY5M4h3MhZ0t3ONj0uP9/0FpNypM1Prhgy+S2ASY3pZ237/65X5b6lo
1QJzq3bD0wAMGruYxCgGK7D16oHY4BJsxFmhbieP0jY2LE2fx8U44PrVe1tsqCxT
dVj9Qt7PgfUJTz36wGQQNv3F056xQJW1a6ZKa+jRi1g2EyvSVbZcf3KeAzww5qTN
toPzENwLQLaMtiv8DzqYf3mVbcmD2BnasUxxnU1ckUuR/CijZAHkkZFemu93huyF
htLzHK2wphUEUmFM7V6o0AZW98PTg+gWED3yv9qbbMf18Le0G03ICG5FQpEcVGM6
iSlmme6TEryYtthunEQc+6p6YekV9n/1+ttx4MrT5+kOEO9IWl3Glp+k5gW3UlFd
LyEbSivpCj4FmOHXBtP8ucV4IvX9tvoU0WOJlPfm1TP5qLHGHFYPEgPhjHKO+qAz
KoIr/OeD6n5hm+oLkfZRJD0wFqHBG/44ZMJHfl433RQy2CcSeGOudZ4T/OBh4XDQ
0p2u0OjxGnTkONCM2Xk2mCXOraksHaEWdbnzDowUMz1mp/F9nCSqzDNmypTZHS17
D80wkqZQQmRVLL8BzAB0rvYg9lQHz6W2Mvs+flZ8EfX46vMemTBXgGbiQ94M7mYA
vlyai4ob3O1RMbqPYqvnNTgqNMvHNO3S8IpZmxpVnU2EvZ875vSfNJ5s7nHKoIk0
HfrXjEush++mJCj9EfNdJQdehsggrRw6sLYutWxStnCKLJ7uyzVkxUmK63q1pnKh
n0VBPV01/WTkGWOBoVAj7/sAe26e9qhmXK2Z9heA5YvYrZ5LggjoxritwnDxPFPH
VMn2dS+ZPbAjWlzmjsrY7IKCI9LyjQaOmM6NSJKN6prDJd+eerx3tMlonFT5vTDe
iNiPOnAzlY6pzGKMy+09SGQnYnpd29MKD7n9NdjFhz1dZnNvs+GJGHvFe7gSBxKA
lORCllw9ujjT3++lwwqG4+NESBqsyqSly54Ie6sYb9uvkdb7cYliXg096dEEXDAT
DAkM5/hpOsh3XSwerq2rmvOFgnAORe/cEdLIt2nzqU4wS2oEkrob/n73/hC0ngKj
PxVIkB6Jm3OPJouDYILwua11BXkduC1l9QhlG4QRMWhX7evyG4H94G+kT5dVuD80
Or1CQjt57bxjwXEBc5UnpwnzdkzpzRPGuicTmTUQR2F6U4GkbwRZXmYxqsQNsjFX
d8tx5w4ikVioo3DZ+qlJZnUhVmNx9HWWsaQwB7dInlefztRIwkWGXNMtRsrexX0B
M14MAvb+09iZoz87i3ZfnnfdqZAAX2540r3apm51Nc8qK49Zk4M7b+hEvlImjugY
aApt5IqUn2VSYnoxMb2CBKOty+vrwutw+cFyhDW+7riJLCeWg0oYamcLRO9MEzUw
zYu/9AT3DquP1kAdhlehZgjMVkUFdqmvA+vuaDXe2NvVA610unsWrZEe76YyiyPC
dQ5uMFbKK7ZVtZCb20euGtLtwzjtErAx1KMpGJC8W/7QBtJlEMn11sWbDm+ptsFV
8l9mj66nZbOY86hu3ztxSHoDuHv16nqelELAki4ot2NCVeBzEuBOpfhX0032NB2V
/6l8eMX6LTQkYAbUKv+T5jhGjI9peMK4L2IMspSnEcwXZk4tUgfaHDEqsTVgreeb
1atbyXzmheUIjRKcB8+YRsbZmFAwg9dVia91+AZ0nhPzQkvuTQ4gd7fnW3ZNZzlc
xsZXYpnrP6kpD5cTGfph1j1Zr/6Kh1nCgZh4gI+5p0jcHhSu07HT6kzSTHQKrBQ5
TcsTSEMUQ1piC88B5kZex/ufRs9OXZeasLHwRfushIiSyAQjaE+wR3QtPxTs5Vh2
jpPozoCjtZ5ACqZTWvFLzTdEads+m0SfyiYAuD2a+0cjg2Zlz+kxx+oUTzeGeEVv
g/wiz946htu5a3eMk9ES0nRkLTfHwiykJJfPQZdfSAxeaz1Q/3tElxnX54sEUPWk
oqGZdBujZWmTKe1BbMCQihnbVVD4wDrHUCEbR+UHClOs1i9oREy9obOXgCLXgmBu
7BhQHC5RxvIFqSvSDoxqdSCqMMxsWGelZQDL5d/0JF/KVUnFKbS4P3e4GI1+TLUJ
2dFjeeft5aiXTc4kohCuY418RyFomzlOP6g/OtnwUNux411kcMLnLmsekHnN3kXV
pCNkZT51+nkUlA9klrWojW5e1H1RVpjE3vVuLV2FKDCa6pWiegfJxvW3Z95o5z/C
tdJWwlOtqN3hqZg/Ffg428M2OrEgsvj/d0zj6ndlXiNUXdWcMOwOZxMOtkvYTlqQ
uPZUl6v8abeZdWX5MQQ9gW/ny5qxS0mzkxZIfcTUmO0OztpBMEKGyWiDzYQjMTLd
Qyk5QI2whE3fkV/mG5rNxHMnRxYWJTBil4v1WagDg/X4MyEZuj76acM8lh0dBA+s
3UWWFcyaG2nfA5jfvxCTt9sV0YUJD0Ym6Qp9QCU8F8QD9kX5dB7/XZ+yi0KVJxGi
p8OMTOfAY2m2Rf021VO/lA2HhWhj991X8xAE+BHJySzyL5ifjMW71QxoW2Ay+1DO
UFbHM/r5OHIhCscM6DyobjAw+arHHkuvtVH/09YZhXfA4MZsYbYsjllin0G2RSRJ
nbmeDC4dcbe6xkQDcBCtRNkDaIgPJOQAZRHrQfzcK8o24dkoFjyK2eBoFmYYg15P
KFPRosZOZKi5ivFCC+Dh6Czx0Pid6H71d1iU5ZQLFn+b2jQ4UbNWFAiFCVg3WiNf
Agl8stfxvDxSaT47cpNSVySuIJXH1R2EWfToJad3me7nbDVpUKQNODKBljynADWT
zvo27Ob/0gJN6JzMmlsu0KkaInn+WizX2YsBpgr1Y2XZu7PiE7D/r3Uba2ZzqCUM
b2rNtEiUWjNMDk+kd8KLQk5mJyAE1PemMDu46KYj/9A37R3uhmf9fblSKKWcSsb3
hd5wOdr8ndu7Hjyki5xOInMWOYjh2rLF9mqh4IhYDNJJqlC5CCRs8cxrp/VPiRcW
ZkbalAJ8ZdR0gOSj6xWX0QqGR6LePOjODQr4nXPOGdsxGz836uMgpkDX02C7Tsd6
/EQNnukuLkAG8u2rfYVw/yl+Ch1SwOHWihvR6v8qmW8vKYxP74izi4HpeogLuUzj
Wyolxg1IC77EJlPy4mEZ7Hch+C5YPvqNpNDk4AEV2rfmf3gRRtCYgwTiYVOuzPvx
HAFMdligXW0GK+yO2sEeNiA6+XzV1Mk/aLGoU2YuyQNjxybNlODrZ7UUSUh1b+WJ
Je6AGro+ogoLr1W1ozWha+fqfHhuhU6Q4H+7ih9bhpv4xPEj4wBpqE5bPoYjYhv8
HuRS5GB/zvduIDoo9kMIs5PahnAaQizhUZYVCwv3MDQy3xhVkGSwUbe4VlCgKkE4
5jnhgpr//R0vBPTonsef/6oIqs8b+jRQ3JTZie1dyhUk2be3Vn4tYLEUwkrdCE9B
33C6yAa0HL1C5B6jhVL5FXXZ5HAzFEzI3HzT+gClHonXE4RLqnHaPfUoCdzTfb6C
rHMeryFrRpT6OTp+V1X6BF3AkSaGApzUXuHIN9haSsHhQTK0Ksm8gPAcNiyxh7Sg
sMD5gOqyX7mnKto8fOwygEDUHQY5DdYgnEErHgG9C5I9Prr7fcYK7O1Gxp6G9psR
AauZics8w5p20uL+Ge3tUXu6OKRNxeoYANfrDrpEhm9nWkYOV8AvAnZ5yi1/c1yy
DCrgj21PC3D3MainNZ3r2HZl/lxJ9eiQZXdBJnkxaALCfZjVXLG7C7rileHK99/3
1DjBuiJXXB6ZiJtQQDMDL1SDy1lFTm7Wz+mK+DSu6N57JmDcNSWSEDqbY9ikj3LC
zqavOymeXlv1jTyfJBP26W7Rd18ml7ENCPmUBg90yKAkyIf8hVJ5BIPwlL/vyAog
d7xKZC3niOwnL3VIvvrJezgPsH4NibT0QGF4o0SZSCXuTwuo3FkxT8L2Rz+cIxRX
0q3cYXsfDYf8qWjUTK/BanH7/LjT3+bHe+F/4oDEN5suawcOo+EAuPiXEEHhUzBv
EpK9+5f3Mqdc9Z+dYzxyGHK4S48xHrkinv7YrdPd30wVmoPQQCJ1FMn3dvKUiAq8
qOSG6Vtcvyaiugzl656iroBd/oylMLWBLcvcCIdE/VeAz6dcxuaE7vn+RoBInacx
tdUS8J1klTEYNAwNYxjQ7rk70DP3QylIVwSkX4O03PgWgp40Dk2dIo7hdzP2LRq5
WLBEBT6BT5VjQqz07wZKEgBX3knTGQtOdelv66KuQ8c4K/QDN8J8xijC9xc1uiY2
YKvbDxQwro2Gs+2XFAMrwPBL5DiqDm1+stO8naYRNl0WHzRPc0RYHFO99+9rYZ+X
Ima1xy+veC37fHZu/qPEYOFhVHlHr9tqx5HIX3MV70sBDutU9yzUtOJbP3JmOIVd
CN2MFFl1yYJ1sF13if2wLPLW3RYbEADZd+P+zgTsHuHUsHVwZvSRqeuCboq8SEzm
CMFJuPI/F9N8sx9idIEGd8Mx+ULONd1VxhiHOTAAdLqrspVukdNrWgbfbRga05eU
BcL/0H5WFpogFPQSELQr+WPGrtd+PqoSYWj230eYtElZ9Hfxu33qK+Et8BOUqv8u
xZjL99viq2CUFlO3Fhdg4M9SV2H0zQqOogJ4PyPabQO+rrlFzABtmDobdxiQS1zi
F5VxCmmDhNBpuLmBqV2rFXr4jwWoDCZGiV45w3/S2bwvIcg6LgzwyqYE4LRzO6WU
b2MDEXpTSqsDcP4Hg6v4uJHkKRndo96vVeobfnGnpJVyAOCsv4yFKMgBUqq03V3b
4yqyswKO4StqiozTrsEiqSKYYC+FYhFk4FgebxQfklgLhSyGdif1bgMVIj0AXn+a
M+JJ7ob3ShfgPoyD01dsPnDuqFHVaQ9kD3hT4W2NU82qniyeItFs7uO6yLQahXMt
74hT4qQm1Mc70uPVdHiHiFzK5psWsSMnFDI1AqYGyQVXIzc7YE+EKwOQutTMaG41
kUQc7uPqLLxYacbgpJT6jt55r6ZFsny4FZxZFaFWgYK2djmmLM8Sn28R6drS7XBj
GocVKWW0Gx2Z34MEN4UtgvL8/FXlgLnSIQABflgNa3RqxICgt7JXXoBVMsFCnyrH
KVZa90zoXQtl3SqHW4krgJENj6pv0pZG7FT3xt0uHYVdd+PGsLNExOSor9dHoihF
haeRu0JenJy+v+eVQHEEsm7GWYWWsf8vQXYoqz+Tdmr5G8cRDOH1VvrZrxGp3FXx
tRzg4WA2NbslmkTAf+Rvg2pjR38iXMxja3orZvYSNk2cVcD44dHIUV43g0IfylNC
ZSk+H6Z7YvTvn/6sSbuMMNRcJA+oK2nbof/0Tgf+gAfPgyXiooGnO/WuZDVZ8D9F
fdIx6yThsqy0DwrL+v1SlzyZBuzrtcRVzDIDtJWNL7fqmrL0D388wkvDjwdj5nGQ
Amhiwr6ahFwtlz5XU2QckfFPyojuKVBjXYPkqKdSEffQN1joXBzECfdiePqNbyZ3
Jbj+x2vgo/S80L0kCmxx26EZFlnyteZM1uiJyqKJdS+FlBNbkS5/zWr7CdtU97uY
ob0d1UtlS1YeYsrSeBsR768jZ07g0fLdHvKW6h3Zfa8eYFAtrTKtTYIsA01he96D
DuDVePtwETVNeLlpj6t2VjhX6ssc1Gl+AdhIZYRAymA5sjsfjAhtRl52g5Oy+n5P
bcf5khYfVuBpQ7Kzdvy+IS94o/30UyVMVr8cIPr7Sgpsfq92l97bDcT3+WEe6BF7
iT1a5EDLzkmBIfc4AIF489RN8/r6p8qoV4aCaQKDLuoer17grdKIIP3Cy95iZ6im
3jIuEww3m1mbj4NJVayPWE06qnAZye02xp16um7m1mFek+WXNDQYKYCdaOTXX362
zHkf5EcnGUrzPITWA6oHiNFR+LmG9q/uUKqajNcNJr6eGEP2uv7gRvrO9B5zYShG
FfLuOlyL9EsWuHVViXf+LNfYf7F7LOmYphWMZqEunV7tqeA00dAoRdNYEcB90THJ
8zyKDSHF6ITPfx0AJri3zBLTgDlJ8NUZ+jZj+rBlFxvUuNEoSB3kliPR4Kw/ic1F
hbW+2cql6QgCAHK60CNKm1prbiuPRAKvvY+kEVcdgGRV4b8jCPn/eEIksMeoxC7b
fln43R3UZX0rpz4kZvW/A7Z5jCmfuTL8wbYG1Jj5P9PvcCusgHzg54vo5PYKLoZE
ygXZxLRcn2ZrR8qeXuGlhY5MyCQ2abdCri9QHUN6ZgOwjJ1eekCsxMfW/tCZ4DKk
cAG8hM6zMONfy312xHeuC1DQppGGIJDBVAuRhPbMMAJ7yjjhFDUvIg3ABJfC0vrV
kXLj6cg8oTGOqxLgP9j9WojqJM9jxuDhI3NFcLkP3EdUm2hGZ+tZAmkoV4AlVlhy
Bqiv4umLNgtMiMDNV8Fexhthq902H7FL2LGeXWEakwkBOXzSCyrxUVl/v/1PYNqj
6qGFAX8zoWEfFmWneLS8Svt1KQIOqppPf1Kzf2ZE/72c2wge9vR37OQeaCXsxGSS
/yd2oJMqHlcpWjaY/ilj8sQxFgFvuBSvMt51rhDWrXhi4uSYiMVNJA2QfpGUU/Hh
9BJ2tGNNHeZnRIDCfNEGtQwMM2SjsX9Ip4FCyanS47Q0BTuXCQmJBw5miQ8f3Qvk
IP9edO32EiHpqObgA1uX+X8z56qC/kjIYj/4Ff6SWnd/pj8wlOOhfHlRrmFzq5sZ
KjPFGZDdwLhHbaPWbdSOmDU66iJJE8WDDiJbngzBAaNdTbB1kQCGuAnjMeH3VG+d
Kgml5fK8frk+xF5zqdEDK10ZrE4nq7kUh6geZLtxLPRBd2kfg0fb/fDg5jW/jWAT
JG7gskL+TMrmH/H/J56AN1AtqGtuklY+dC88O20t324o4F/5TdP/xefberjYOyY+
40OHPZcB/Ul0iSuJ3Rb8UjWkWX2AECH/mQ7rlKBZ6enzf2MYFDZ1wywegio9U8lY
vf65n3TjSmUN5p+qUQESWBj2W9LSBbcmwKYOsHcc/q5P+C1ohYWChzFpmuVwURcm
cdMBq/mDKX9I0HMQiLWCTidG5o2ql03Hi4TlNDsbVmq3x8WUZev8C9gflTkcR9NO
OCkOC9U/qNq7pWtsdrycdyXK1jsoU84eqPNQQxjcGzle8XmdJoMJYL6z9+C5JrhR
d/Fxfg7fnhPJ4+qLxCRyC33g9Zms7fvNYBf2Nfp2HN8C7/6c5abiZvIUTh3QNcDJ
XhH6Q1Y0kXauAoU4XfllDcS1aFn9ZuvXA+wW7V8rvzy1cyRI5lNVC8/H05mFz/gi
N/m6znxXM0EbJeQa5go34UCmTYs2lz0ObrkfYgX4JeB2e9YVyBjTCclnTy+zB5yf
DzNZ+EtJhxdDpH6Ux+8wGwJiy5ALZEGffZ/dibC0bDyNU9R2I0lkyihnUnDwi76/
ucH8gFdJ6KmphUkioez5iFjioW6iqUwwpS2RP5K2UheM4LIZkMjYrTIXVhiyaAgd
3lqd6rG/CfYhevCzhC8wHw7CKX57GmbQqIlsbD6LjzsvuDTMlw9UUCE7wjueaE1F
IK0L9oSZGbjRQtpPIMDUHvt+OsMBMqsYLfelH6ZeRQGlzZZdywLe/OMXUJVWxvrg
LyYXLFN4oj5P6M+/e/8yajFa8qAcbWOyVWnrsFjk9it8R5gqCjm0c51aoT+Kkuiy
OSZPZEFCKm7Hdtgpmbr9Lihy/Kn5hXJsGpvxKvWE12q0LK6NNmvSJi3oIm+1sLFE
3UM7LdjHQPSaXDog3w+VmLPq9hQmJlmbpgrnXaljXydagqLxAd0h/L/pp+A8u5xf
yR9qAOfphjjmS3xYLpNrZtIXXP4LFGLgpCBtY54Blm40CNaUfWIGvx6XPjRveOsI
d/Cb/YeEuDQ+5HY1HRuR2G909U2b/ipNRGtyEO7iYSNfi8eMabSi/OnuxBY9f2Dw
bD4Jbjy4gj7kwj/npVz0/CgK8GLLC0Gk6N3ixPINNQzEWIi3v1eFn9+SSvWyfIDY
NKunyNBIsAqZV4T+IkQwQ+lpempD4o40/osG12XCgfD6zEe45V58x17Lb+ng3Nxt
hvtY/J0NkPdqVPjouRRnJYaIRVekm3KiH+wOsmm8K76oHgh0FkABVB7aiRiQt80c
0aR6AVeW0VN5Y6lJrXCMPsmFhLb8g59i7lJXjk2Y07++pnP3Jgr/SK6oIhNtsIXm
91yp4UqIbSwZnER3pQWhfdwKMvnIV6xiF3TWcpGWPCKgvoQZ1oputIAjeEinnXXM
lwWMiWXpOJkaCiPYkql4Ih6c3jlRjjffj9jsk2Sc27ApcxDCK0P83rwox4C/kAOF
k81OjZ6KP/HCxhejBF+rlxNfgiiP5SsmS4ju8IE7Af3f9X9JtmreQ+C9k90rUtiA
I8RQF8MUy99A+UafG46ZmRHwt2IcysvoMDaYoGk/EXdkc8mHdrw0nqfQGwb7sjpN
/HKoQskN9O+HEdInoL+0u3RdTCBgISmOMWl6JF0ybbBL2w/U9SDTLOUSKWhuMRTq
vYQUkDBZ65TRobjpEpjsjxqIHHX9+W+gbwcYUzVA+iEzZRSM67zI+3BrUzUmxkDi
efCIC3hLkvkv5CaOOru1XTRoAkzCs+q2kiDidxETg9VEeJhNHM3GCQn40M6sb3Pt
DOiQPWgwOPAb8gQ35niacMBhw4K445sY2ISNJr74WZzOc9HLnihZ0gnx6L3KQ0Zi
iO7WBnA+GY/GlIFY0F9KAkctkthbwpwm1qZTT4F8Cg1tib/DdYzzvglIFubmRAKP
JP6ePJQ/G810FlDX/eIwHUMxCf1CjAWcNihPH9KenPzcVqZ/elAQf6B1U7Vh3NYq
OSIfhrMmzvZ6Z4CDetM8vv8+YdjXbCBlkRmJPsCQWGOxjx3+gBGlJnQv/I86K0qs
PHaGj/aqA9eUd+3yxTB83RTlm3vIfYYcMz41vRCb3M3ile5USgmLFGoU687oJ0DX
xuZzafg+OPyHQAiq1BjPeZzo8yvKuUx3mQhvMku3dasH7xg0Uhs7/HMJavToh4Gc
VjBPcJswMcAU0tryF9++DWuLTRvBZpbOs5+dzMYp+sBwXdE+yrELTm7JP5EpadKM
5scwCRMY1OUSlH5TWAbqzjcqKbHFI+2vGOHI8w7HE1+SaQRHqo/Y0IfSKgf04DPH
/4O62J9lZl5Zp5PQcAPog2hSSB7i7TNDBqSuPIpvJbrWa2QKYsjL5YP/vkmJ226k
lsP9hcSi19VyC6mOsRKOCY9iiAnV/uI+0yGUNfoAR9m532+i0r6nO/5jV3Nnhp5l
kabO2JdrbwaUkpGzepni28roQ0lSaUrEjzfcdrGDKs+GDEF8PIQpNgebM4pQ4AGX
XioqwBWXpSpXEV2ROIJwro1WdY6dgMS3vWYogctHtCoeEkVGpO+TYMM1acufZYd4
1IzNnrYbNxdNKVttDhguMp5M0/cgzjMpSHcNZ9IEcFR4b/H6EiPjy/21B0LTYyUq
nqABk21DAUnLWDqYHOy0opCTEAaoa/LA2MC/v0W8SzAGkmgasxR8c+I7P71hwpn0
866HAebAgpYuu4+IDVvMt68m3a6b8kYW2e5PO+HonApq+IHPrXw2vCj/cdhzlo2w
Sky0C4TjEw8uLhseADZMqJQi6ZiRhCtuioA/PSacjcVLvVmpc9EXxQo0Tm1kFI/3
7WVdhKMyiTVK7GuSBRkTn4BacaESY4eIZp4b6JfD2DErQn8qG3OuQoFvbFkAtMem
uedU+Z8ZCbDe2RXg5fYLTVLZtaCZdRkNOSZt9WWP6WlgnZSWFSl9MtruATdtlhNT
gTbAD/GDwuFfsS2FUb/BUyejiwaIj94d+SRo2ryNi6uebvoAjCFek+nRubdhlgoU
KS0lKwTMdyhBtkkE5dkHGruTufFHWKei+wIBW4LqCo9cf44Jt8MUDkt1hqiPXMym
OQHJPdE7P6rQqHSTKnYs/YezgrHodXNM4BgOhwUGZPEy3iPF0FwD8RSZXQ3l6o+J
Fxeg2CCH4fsn77fhBHLzqvfcKRbi+wX6EeB2yQcdi/egwOrns5CF675OCAWSZ9jr
NhhsDf+qtEn2qZP+IPEcNoLFh/w2dBVluIbYbDb7pobklw3CQey9VUpeM4ce9yGi
Zok8cNf4KjhNL6MfzWE09BNC9U5RdndSnbTEY5tYMbriAPxjfGpY2lzWtbPvnCNO
e0eJRW1haw/bVr/1MhLFchA3JuMJplhtmbZ5dIAHzC7tRPP/kXt/+l87xk1w9oO7
vJCGo4XCu9ZuK7bxkX2qnVXxJWjOr9r74so+fFekCsbIsgpdA72KXfkHmgf8jxm/
82QBCJjMm5lFMwmI1nkBo+AL6+t7MXBB0bJ4YbYISoGEFKetcTDdrdWFoG0ef2kv
8fbqZsRnigY6Zu3vJbbNaHXVOP3JpNy+cLrvjUtIQP4PYMHrxdItK9obJSY0nsFF
hIB1Mjun06QZ5E9MphVtUCAJAHl+Ykrz1PsgW+wQReDO7zvbfvGYgAb+m64BFxFP
UZmwl6NuczFVL6GTnO+G/A01oxFeuExgnTLWrqnTsv8/+pUDKbzlJB32RxRlsxeW
eRKTxix4qUu6jc8nXrDbX/J9FNbv8RPCReW99bB8TNzd5SfBZGzItxGWuwS3sn1f
SdrLRK16Mw896MykC3TdxmN5n4t0surClIPbf2EhFH26tSHxXdZOjd7/pkG5EWlF
aLk53Kf6ywLJWAP030HObL5quCaelc9l6rDQvdS0VzlYoOHZxGpZaIsd+y+tHnjg
1W5QWMte855Nkd1sZSyq1qUOOjbVJgAafThFxuycFgy8uzG7hFEvNnIfw+XmI4I6
xuR71139O+cgq5w9JO/QwsVDX+EAkSMVHrb7Wt1NjHialxn+e+fkTmqOg1PCP/xl
XEyRzrWcGnFy230xH44lTCL5x78bx7HZvlbu90A97WSgdmgcsMjPdtAWQNJXyLgq
D9VpmaJNMf90lLoLtgVsFCMTjmi3NImE2ZcMPaA1ZLDTg7q9sUVhTGyruluCR36K
AYWRF1rwykuMgQYnJZHHKD8r3ypmok1wh02QSvtq8Y5nIDXptv3SLnnPUipIwG0/
x0/elmcSz362AJixFjuazQCi2+S8Z4z6LtZx59kvkNQdsxFdsOXC2SjjumTsDvRx
w4jI9xLZ5dhzGRE0Ctr9DXLR2c5S7oTSfjYdU2Fzldb2+MwlGOs2JVKvBnocArfi
37PhIzI9jqz8dCfmmGNWocWHPEMLXUpfY4OPbm7dt/mTQXUTT/jPlYrpJfNfY1A6
JNvVDoFrMS+1yXKLB3VJpKHAK80iSN4vAqxOpRLZ1kdcfCjihmfkER92elGChNwW
4AMtzzO5i2fawaOUs5o6ienIxKy8O/TuDYEm2W/56fgieg3LnRbAec7+3oK475cE
e/2Acp5fYy4n/pjKlIDpvGNtoui8dFq6/2BlThEx40h5VHoWWGejZxn0oifGR8R8
wxQ0OaOQPzBmDWapLqNFWWNH3LdzjAH3VRMWE+isgAwC4z1Q4g400N5BhdhaRDiM
/761ZD6bNTdOh/YNsp+BOvK2WXr+oXNmRVJd+nooKS10jHgV5rImJkWkXu4K7F21
zBXqq+d5kLkhV5+JtXevQu0cYIBFGFDdwtzATOgCajBKEQaKv+4kLOWjaa+31mrO
VHNV+ziDX5t+eX5zdnVx0j5FOiTH/0X769Waauu4iuXwMhINgZ7k1CK8V4vYSi9B
TzQNG+sM0/qGipir3hfYvBi0iYnQ4YxN16xlKmRZnO64/EAiZGl/hL+TVnzOP+b8
XcXw3jmGIijwIPqocezIVOWGI+gOOQE4q3rWV1ZMf8uRu6fI3X11UNRwPKph5tVQ
3/TV+0L5OmT9d2oCIYr/PZKsb9UxdIR3AKNr8/pGHVjp1BrsWHDc6RJrMeNRIDma
+5LUSGKtleqWpvCarxBgmcXrYpEtUbXeyAsf4bf9PJ0Y1O982YnJoCt6FOqJo0Qf
GjYgoTGCdylzsYfq/+Kx3P0OFnZONkO8hpB/CXj0NavkhH/2HDxF0NrV5vimavzW
dRaYHE/loLefzR4a8c0m/oCKHH1ap/TjMR93c9gDi8w0X7CqVPRW+i2fT7v47s+l
nMoX6pkQecOcH/6moK0rxJYPaJdKLb5UEhJ9dQFupbCYfHaZb4/4Fo9pqJBf4FhF
pqNa9TQSlp/HZl4SfqWiMuzjwTUKieqU8zr/YBFkU95Dw39h8tI8/UhQ4BdEViTv
0aomZqQdBC0HJelw+lvZJktiK/bFH+Wwg6DeAGvHRl526kB3qzG/GHBGW/u0Py7o
lA3WZRx0XrgMg5G3Ttl+Mo+f9hqy9DRWBgbnNtgD2m03t1aQszycQDdmXYYdi/QA
1jROJLBV4C3BWNqqcNu55dI/MBuvyaqPKbhLJr4XEZ8kn5lk1HSKn4dxLkPD9PWi
hKIERk9FVH/aM3tmqE5JVc0I5hyRK/3ROVS77kMNORmqNYW/8Lo2GPvOgi+i4fUx
vapCIONUGUizP4yZj4/ZmrrWgpwSXh/cElH39deqvt1vC8QSNQnRz48g7OcwvFaa
stbZkhI5+Ge1VpXvdYO4X8OHk/owkHDB3GX+CanToczBMxfwhM/AuAwqreqy9DK6
/YUCFIUS4LBd3NygxkjSGwrLaRyyHk9V9bf85y+d7ZX5l+HZ0JbZ82T1TtbHmQDi
HfzvRi06t1mjWwTB6wBrmUPt5ahHroT1ara0vDjy8APzAVp6EiVEA8eM/O6+sbxH
ughKw2REquHn0Ev6CqsehEGAQIWedMSjicgCutndVRgig7kynxfN2JzArxChUlQk
gBvrkuF9SWBC25oqv0ApngtIBcK+KPguJwL85QOJ5y0bhsv7kITuAJrelG9/3eP6
BRUcpIt8YqjtnkIbsloCUsEUGnR2bdYoOxnfGAdnpR0Xm77Uagu0kZbAztoaNrl/
IGHFYWGJcv+/RSEa+nYpnUXV+L4QgT5PXc9d2yDxfY86KtUEsmQ/tUFqm7kPFJ6P
jUzOMTnK/kapoXV65LrxxasbDM+wvoLy3w1fn8HnTmgerSWgBf02fb4eWRot1T1f
lmpYvCi6wGnAaoUxzKxZMoVKU7+7vsm0iaHwOFDm5kqPOuBBAp46O5oY/Z6qM0A0
T8zYKoi3gLIs1F3bMtTLgFyJ+HsttOVMdirOf6CVJu8mTLX24+WrVqqnUGtVo/Tw
K47fvJ+UEplav5wmB/ET0btG+R8g4HUUOkCc7p3HRFKuwjNKLCYa8u/tEWUi2dN8
NpfAZa2jVH2nxkRI5GUZh27MVwb/52lYvPDA+MYUHSVDXAb0YsIudbU2yELH9qFx
Xr1eo1xXeZA2D40IdL2mPh8GGUbHcKk1b8XEPbOmZKelh1MKLH9tkm++W7Nlm3EZ
sjS4giMxyWNPj1vYF128ldZyS25B36ZSk5QNPhCG5B29DA3qeU1/UNbVwIdUtnVV
UQbE8LpKEwbyzIZ3/JdSJr4J/+CLmgQcjNnWradGzhgYgToVA2jx+/Wo7rej7hir
Ym5NCIPez9NYFg4TUSQmtgknOoRNOo/F4PW9H7nLZQ5mNE7dj9nDhnrUvDqZcvxm
Wx+WnKB9Z1iXr0ochITR5M0T04C75iiat0EUbd96FwslMIKPWgNnchHShLwQTbN1
Z2vMR/Q2psxW1HnthhB4Q7Xou/NlPS6yC7eV1XuBzH5QMETBsgvSNNbDF4d0MdEQ
OKfVjtz+3Z58oFgzJjACG26q6l1Kt3Fau0RfDf/r4YKLVOt8n9TKV4lAi7SCOXZ9
YqoXAPrKhmORYzEt1kGbVj5siusrO4kMOzEQQENBgGyBq/Cx8ONOL6lgg/UqOyu8
uNJQ8Z45NvDfrk0bVe2vLJKacOzTjd6GssAr3CeT3kmecui7JaovICZqvfOAGP4o
betJTHPumgeTdsV8iqpSfCVnFUYV8TnZL9SzPlUXpwY2PUDlpW5peRiKf0Hmib8j
2USRHrj/IJPfC8N6CQgh2nv2otZiErYaopcIfw+6Xh41W3p4pf0U87FEGQKVDH0Q
wmaqErgl+4EcXFSLw+EA9RHxZHgsGFjqRbRmX1M+U9djvyIdTuGSCKyV09yFu4Bd
eRePt8ribho39akExz3GfcT+hbQgy64fAOtxGDSEUypa/LqD6ZlpI3S7EC+/iKwK
IHOR2s/HvtmDSe6VRfEixZYt9d1N/DSuM3LSY0B1ILgwvFAEB8dVmhdHuNh/bxaN
1L+xITPwPSYYqR17BcpDnAhH0D0HCA0MlPnaLCVAigokoGQlKCkixdiqoZPvykK9
2HIoGh9qWGuEH8ha7Ybf+6mqOpw6/f+g/tAWYhiij/gA15E9/P0Gfzmeu0PJmDlH
64mgD8BZjmxb4WnMtSIEjFzhCWjTasv6jacQp6MHKwNBnX3GyidbrN3KolC+Bllb
DtTjEXDnNVqX7NFrw9aoPnQkA8HFKd7I5UAahewvMz1geUQQVLWpm3h3FBRQzkel
dQgMast5ff1ZKMtjeNyOhce1+P70hOPd33vBPITWO1roHZyzv4mjHLH0ilNISYbC
sE6ULyXh9qRT6ixLstj8kQs1kfoAmxr0gTokByxpZfaU9B+geNKX7HseaJyBRX2b
QD4OrZyWhqPWTcSAbdMWyBmJDORkIRPTYprR4dASyqNWTPK/h0PPPpQUbJXrtZWr
oAlXgSPMfM5fj1BMA/G6dL+9i/W1SomyzIzmsVcLO34ufnuUFnTYRFkq8Sk2Zse2
703MdJQvbqmEhLDdary1g9gqnv/CWRo/LDLmX/lxPXcPLc9j+DQl8Y3pci0R0oU2
YuyjbeDmLtRtfOfcpISln6NEC36q+3ymBP+TLGtSTX9RBQLvRkSDHuX5HytFjaCw
8IaaZVGhJR8ZmldJCUyxhj/9QHndg9TqwWKY5vCUzMbZVxyXO19AhIvByuBxj24B
fEQbllcUiYn6lCYgS182UITZDhOZ325Io4lZiN1x59YdY3Q8OrIj+XUbRCfnwvCI
xc8pjEB1tjFoDtTFO6ro2niR0Rb+Oj+gGAXCUnEUzBEujS5rtpJkJTEUN9gtNTM4
o4kORKIcKlRFwV+n1XDzx1P+PdFKTaceST/YVxqwYbbyqQrHYe/RxnuGN8E+pbxp
/fwngUFWbsNt46SzxlTJAUIMe6qHfDjfw8JsjvVi5Sv5ckmLfx0iHxRRVUS0Vavs
K2/sGZbHzCRLDUoH5oII+gnfZ72rXymcqmQoIZR7j7WJ+5F8RIYyDAJ4QPuOtSJg
oQFdqFOMPuB185jTjXYexZBgp+ZJ50509t9bOju5CBoF2ptItjFSkx8G6MgkoFeN
M/Tg/+jr6CgrgGRCPqihBmZySQ44sdNjY2erziH4gWqUSfjIaIIDauKrRtqNaAdK
5vbAx5FWZAftc67Ey5O077OXgD+cCyE3gyFEQfVXHl4e3kjnunb0xITRUm8hLYzk
2Yw9PqMk8dZWH5/C2IUEz93WJTONR1MlaQ6LRuOupyIEfdyd0oaOZcf8pDvb4rHq
BRKOSgff1GZUe0hRF2T8dykWehaRaGGCzGUIwwWOUZXzqV8eCWVpGpn2ZV3SIrtH
sICg1567a8HuA4tqukarPdG6V9otVLA1+SDQ9jrn37PzpKer9oOCGRTrbEM5TGhc
lGnXVFWp0tfzhYgiaJSa2w80oDDRnQxTi8bIjkhnKM6Iwi3KmT+HWSZPHwe6uCw2
EJhOiMkMl1y3L3cNwYTt3FlHQRKjFMKtJAnyOt42i5txC+IWKJzEHpf54motw7pV
HY6jchqZDGy//KdWKFKqDCu4m/QqUU9Ng0YnYjlDYLcVcqLUw1T1wyt0uzftKT0Z
CgwYXKadIIhcAuFFLKg7Yc1YmGBYIKi4Np/0IHj6ZmTuKPnMUeFGPyyiEraGlWzr
o6zxY+b0heEhlTODXNj5mduf5TNBy994nI2f3uhp1xX4AX5RPa+7/HYp9QzxHlCI
sTYL5qZWlJSmqIwkBYH2bMZIuN1iOHvomzKZWSKR8smFZW/lM+eAn28lTQfrSGLJ
YUMGI2SqQ561ul/Atd7XuRcvvHS3VOY1eNSTQAomEA/t/UylVpXbWCXiQRj6DEy6
m+VEx5HtExnYCsXJarFNcSjOqUTdp3IAZXqCSQ7YLCkB7VjmVGk01nunCUx2U1fy
HsNe3v13/wo3v/YLohJwKZTjEXorVEY0hP+FNgUDWcm7RwkrR/WuZLoMW3rly6F8
Owy4XLYqt0ZguqoLKNKwg0AfI9qsFoUGL2v9aSAr9HvH4tvUbY2mdaD0dNkKewZy
GX6W5WfjO+pQDgdbLlzP6/SRUwHxgAtlgMPxjqQiyGz3AxluaYJcT/pJpSp0C8st
CqBxLncAftfZMUisMnrB6FegPatsX1AgarVued5Tx72hH/hc/fUaEkn1Q6OrKZUQ
aexJl88uLxJGIAiIr/xxfoD1DcCjzzYs9petzLUyiUW0gZUBasklm+tNogXxnUb9
ImCl92RHNxO5F/CLouDqZcNPcpNnUGWhkMQDdqeKqkY/ixRJ/OpyM1DY4FIMVSE4
ZcRtAlB0YpIVrVnY+LjqqfwEFRw2o2x5h04x4z/ooLt/2NH44x/iZDToQHjeqE7T
K0NVuPRgHBYC87yCuI3kwG5fQiiOmkvl9FisFNTk1jq5IW6YFKeo4XZyfFhakwQM
j5XmnVMBsXhc589yU1+BqCvfuklHfCXHbq82T4IWJxQX7pfNAyHavriNC4V/MVj7
8+aLr5oKrCqYVghD8shd43A0TKii+PMT1UPV/wuF32mhUj35H2gi6Izo9n+jhcOi
7NzhB1tzz31Bf6ugxGRN+U6uEfnvbM3Y+V8h4NV/r/N0zvgwVMDS59N9dZM4fnas
LQIKVHod9zxUlf2zsRlsvx7oAi6/tL0tk09eoHDwsn/9jiEczQyGcjNqdx/V+xSV
FQZIzB/vNt5mRUOyroVPod7mXIaj6WqYgq5YgLgDL7JX3tsXM74CfTwOjrgjpD+w
LhEMZakz52fJ31PYachL+BENZV2GJtVmpDmqhPL2q01fNA4q2vt8eEi7GRf+h/rK
SJXCVMwxtUlA3kZcuiaBsfHSopwdBkY3k8oxOnADlex81vYhshlJbyRBIriu9/8n
KJ1cDKok7quJo5sAlvDRWvGe27nqjbm1/PszSUBNmq9L9X1evdedW3TpZsrlVqRW
OnpubgUEGpUZEW71AbMrg8evfX0lUCO6i0z2160Gc53hja0zFsj9WO2GPNxZgB1s
VyhA1m+8BSXzTWVukblUHTlPL2Vb6nTfVwy94mSAjwts4r+zAuW/CUsHphpXsafS
tlQ7HEuvXUOZEC2K2RSze9xz1rAQX2G9YobJjcbbln/lpC9s7khppdL1DtrE+nQv
0ww0zGjFSWzjBOxqr4ukOvlrzAL/IACaaH/sKlMGIJJOYps8k+urJgykQL8CDbbm
UvD1yp41YQED7r4xjpxJdsZq4Axz6DuyNE+CHokvZCvGcPI/gY/1/7Udgj6B6ZOZ
sbcW1pyGeze2yEyA+jRetHfbQ4c/pwFza77ZmHD22dS6J8wsPu+HxgELeiZskAni
fPly1U/Uo/ulbQfz6t9v+MWCBqmBYVjIapmcEuxoL54kEiVM6dlzBFuKcbOu23rj
I8vNLfzDOfgR8aK8Ms/pk2GITl0sTAoi9vTxtE46Kt3sDWxZOyo9td2sHLNZBhW2
yTL2io5sMUZyX8HTXkArIckyBCu/v+aqh7Wz0IfujxbueIlCryovg9DB0XiMEVjh
v7IbYKcpdJKmwJQLeeNsWpowtsQVVE/br8Cz2hk4MrKBxALK9o+41MOKNT3HUbRO
K6DQF8Wo2REcUUOQQtMLUqC6p49z9tbaCvXvx3RpQ1bVae7KpC7avC45FKlddPVC
2byWvjV/HmQcz/RXJNEe0uizxwH7o3lfl6PXGG0XMN0lwOQDK9rp7rz/TIudsSSB
Z1zH5QvUkEiPRtaFgcGtHVzMiRTzxz+vR1gRBQYkm4ZfMhzrOvSQMHf7NU3y7NcL
Cny1VAMz/9rVskak5FEXXZYF5yo3uscKsxXAZ4LiKupGkikMdyQRUKFwrP4vhyLC
Ek+jX42xeEEm6YhPG4mUv3TjPoCakkYRUtU9tq7pxolHXkIbrpoQO/Pe5vyvi+Et
1j0QlwC+qt4ypj6eqd7FqAfjTutJ5uhRY41myauYWgDMduiPBI71OwT7OV1B4qob
ewchCrK8f9Nr9+XwdMOJWC5jgLEttJxqyfid+TYiWc2rym74loHl2ms2yHPBkPFw
+FW7gHUIPPTah5h+xR6BQJ9ZOcHftOoBd4vlnMJe2WZ+NtXRsH7buKlmTDFJai0m
nB6RSDK1DhEV+nWNkrsawboryG+bfrdU5brNZxZ7RO04u063uRXTj3hM5CJTWvaT
XJJp8+OjPrLTG5VA+l7wTanKO4t7qEn+G9aejjQ9XCYBfedp9NGYpRkzrlcjKJlC
5QZzEWnOyPJLZrXh/xkTjg1tiW6EuMRvhk3o0PDIL0EIzRNnCeEnoKaGxqY9XdFk
3qWF+NlJwLQQoyfvBVkRdTI4Fhx6e5qfq6bIwUhsgSRpb9WjtdqCN3DkkKwKQA4X
XEoIhEXmRgbWE3eoFMnkNyodW0eUSChmEQPVqhsODMy32OEcVG0/+Q7rrqRpAE+9
d06exJ2VVi44ZSu58fK42JLHvzkZF8eBIWWNSHhk8Qwr6DMn9U/Mx7DzNGhUd2Gy
Nh5Vyw3ZW6vkdiBbYwC1Whf8OoKAz95NynFTacpssIsfDOP9Gpwsw3aPr24IeK0Y
yHJnAm1S8w2OmxwTcfHSXR6Z7KLvtuKMtVJ8zZLgc6lOKA/g/JqKw150Wkv6kgSX
tQX64Yd90aRKzRco6Zq74Uom8U85jKfhTej5BIXDVhFFlOFqcf1TF3LTPIuaaczM
VpG7RSkWx+P70w9481a1YzKOR+pyQ/hjB7Ep5ZxUnsRNKsDNl6BQjZf8ZDS8p2eF
kMzyBNXJzFXgXbUpqxuxp4gA/UuFfJwdr32UfzCIGu1vtn4bXhgX9x5hPbOqCtcI
BwjZtQUw09SoGxi42Lx7p7Tj+V1CjBL2w3PE2r/g+gxp42FF+mmjjG0LZb0WIZW+
ZeeFJM8vepVCB356d3O2xw1ASHdxIVscINpr6GKTrpOvJABBgeyDY/GiypfFCdkf
lun+FjFtuR9nIRpkjXRqBTyIKHg5VdXltEp5xeq1VvfYxY1WgSy/BpSelNM3+YWt
7J7bgxCNqSPjcIsUfukHniUvDXb3tGTllC/KJeeKG2Lq/ZTftKEv7EdBYcUQpmLR
LSW1V2fmQnquE4cxU/Rd4f41nJ+6TkKY1llX+83Fa3b5kwdqIrHkmwfyAY5h5Y9A
Y7AjXcItX26uoC+M1YcgRJLYQyLlKbhVfYTbLhbYIt0ONRyyRuUgGWLHK+JIwPFw
V1GUAxUfnA8O2tAkabq+lmMS/TCM8zPn/plJvXV2DtSwH2oDWE2XF+CKakCYdfan
oWZig02b3Y7fuDpsKllRDZDvmegZDZuUAFNTcepr2GWfxvj2LT70pTNZb+MRWJy9
wNA/63jcnHsQ9jyenpRBbuaas0hohOmQgXl3q5ReUThxIU1O1HbegDWvoeKEKmiY
72/9bbQJL6/J3Kqaj3zv7rWGKQGV/wR83wzdGH48ahnbF8kv7ByP5nZjdbw3QBW7
JpV2KvI4gpGLcjAmx8m3Pz2IbC9xav3i3yVzXmGW2CdhRMS9YPNbZI+QuVRJSF3w
8hFI0SPAIkBScY+OzFAWOmOZGIODKt/Ll8BxdkfL0GkqFjanqvY/iDZxCi4tw24d
+0ysYFm9osd/0RWkRPND/qBt969DUk1Ec+/GoLg0hXaWzHbnk2ZaGIEt+nywJ12d
f5ADBBl+/Fnbr7uO8+np2DVk5CwA0ntO1fcVOENejWjCo2lsqYJoC+DixlMYGwUD
eys7Kr3lAryZC/l4dwaj9813IcC0xuBnukQ/BToqHzdktdYy0Z8qyjePSVhnQ4ME
17YCcPpZs4XeZsG/qSmhmbKABFCGTjf6hGx9mdl3w1US7a5TYcnm1nhKJRbt2eZ1
zgSTkX1n0knqH11oHVR+GLH7j/mrCpuKFGzYuITMnZZlZJ+cRSYEF06Fd5WNB1Zc
bzwxDmH37PH21JN/Egal/lSBW7mXvVF06sm2tLCsk0sSbVzn7bcBu6tWMNPoGkg7
RzW6noug6pHrwC1sHC8uegDAgbA1hHtJod0sg9BbFQ20OzGGh9PaE0gbNtJuIODF
tg6OxJmjJ6P0yRXH2EaNfcDUCZqarvIB1Gy3atR+mgq/uYggw+5vhDDcUTppaEgA
n70qy2rDzJqdcYHzdkZaf7ffEHi9LKTi5WXOlXi/fq/VTfzwq3eMA+P+paAp2gnY
+KEBbjLp48iENe16CySfdHssAWNFruU3cKNBUcSKzL4HhPF2KSFA2GUQlAJCuSzF
M3QOWsRa5mAQvbIEY8E1v7bVyyluCTvaWfzjGEASWRDbLrQE+lpMRSJOPklkwdYj
Iv2KAfhnHpeqkUap7G1i14Ds6rP3L9PqEh5m0WoJLB1rywvx6AzFtvzIC2EwRJTC
bv65rMunHG0gbJuz0wM7CJa6sMCjV/UMaLwv+BfK3uU9acTW7X+tXqppx8HoMItY
T5lN9CVUJu7mLsF/2+mjeHgfS4Wz4QbxVRAYcQ5qVLZfT6XPRubX//rjia4zah/N
hZDagfRJKFDdTbqL9sNks9K2q1ZP6xA5Y772ibkZRDSwq49BnMi8nTvbTpS0lzbX
TP5hx4ALJdpmSWDXNJiXR8dCbXxADnVvWpv2ltGgUl27a7sAomXy0Yivo9wz0B1e
hjOElcyZtORc64D0IpYeOu/blFegCtabnqQGtx6BxeiH7slj9YhwQ80BkWkeiqM+
8tGZKRceMEyPo2dvprJjsSqoTeJqun4EhFTramCZ/zWEAt75UOUOo9OVbfFEXltE
QQJe1sXbfL8FwagMEpHxPjwWaXOtx+cs/5ePj1A2Ay71ZCkO5v1tkXy73DspqCJr
faPTzeI99PAr7S9WRixMYJb1J7YeFEgmoqqLJtESXenCUDZvDkfQ4dge3sVEMe++
AKd6iO8G2tmA14b8gx3biGngVLLTJg7if1mJx7HX+srkQCPRnNJDNC7lEbu57nhO
/OyjcYrhq5Hg/nzzsxgzVOdDwxN8WJmlYv/wWHjvVP54B7fT87pI9FKaB+DAKbFT
R3brEFFuOmA2XapEv45Wi0JTOX8o4EyjYIq7+iH0+es4SmAAqgdsCyVlzwUQqHEC
LkSU/+iAync7urRNN7zGpqvCldCmtfMfgbvYruWxuxu1r5s4p8N667F/kyFj08Aw
1m6mpBhGosXev2fOR6fLVnLFW0ohsERwjo5tFFLGodk4v40ROdFnQjsetDc5EXuI
XUNrulvhKs14MyH4izvZqHeTxqns6dKN/Ls8iD8qTC3jNsti/pSACSIFy74BD4AN
lttYZdIdR7WBkynrVIsq6g/7CVo2AOy7dNeF4i7SdhpHXqa94kP83+bqRq/t332n
lyjmhQ0/VnGdcXkDmMgVbZjYZVE7awrMk0FzNpez3bLsOJu33FgyR9EKrK6UA9yR
a/SLFlaRBByn8b4h2oNgmxSLrhHz9u1aMuVnbJwLPSVPd3oX0yyGdnKUn6FHStFn
igUGDaPSboQqnTO/DjsH/BDzKNBUmyRHo2ly9/fP5lJZz/bJ0Wf5+Mg0dHytuyIj
3CtwLMy9ldL9YW6Goqb0y4H2igwrUqRj0nL/MYSnQ4TIWDzMkAKIkHs7tSX3dK51
AEgqg68aD4tXxZdgd0XQ35mX3dsE/J+NM1LMGZM1sfIR8pZerw7jtAhlmlw71tSr
7qH6tLLkSFo0qNw6+ljhOIUTNiL+NtoypznbnuGDrYvwqFkzG5uLM2u+P0knnqOM
ysmq7IxbdEYnoLNYTI1rN5jixpQJQvc2Dvc8YW8ltealUkiFtrj76zawaXGCq3xi
C+p/hz7RUFYmhKqNS0U4YjKmWy9THaAdkBDCnh5fVCHxed4w2sbCbUWykKCZyIbl
JnGMHbEuPZ6SJrDeqhvDVdvBkFJ6gXyQ46tZHqOgZp1v/4WmnDLrR0jtacolNPcC
35por9+fHoXsdJcYYz/eAew+V/U96wGkvONnGByCbSENwqcCOPKSQs6JPz0M45Cp
BtB7bMe/W8sKoRXZ121LcC8TOdlkJ8tbq0V+pthdXWj6+DtWC5qc4EIPCIslRqvB
/19FQRBt5N6T6c82hSe+HGEd7nBAio+EhVN6WNH7u5IbFs4NzQjWsv31rGERajIE
Ns8Kq/kY3E45pw1vsTIwQeC+jk4sScfwQpjr45onwqzy5XB6mQgovo63uK2quvNd
88JQ7ZjkwD30hL3DGRULvyLuSQaBiTQLybS3Sx1tCuZiIXpsBzE6z2yqTBfs8RY+
S2xKzaQRMK8xq9i4Sv0pExkzu1LuDrheq2wP2891B0koCGOvqTN6C1ToUpGtqqVd
MDIZQ1zfifMVX/U1VGvh/RhwvviiZ/WhH4B0HHCDM8wHFMuNT8mNhUFfUZXMF8YC
U5S9jkyxTuGy1trdtM/5Lrhjp4+dps0mVZTyx8WtDe41CY2QNAxEUSQFPugp0tDN
qDYWeg11phLbWUmuWTQNut6pWLHhoT+Yvn2GHTRgb4GYiQcQnXNlPZ4Q3L2PV+kw
8AiDUDqLrtLxLKfKTIPC0zTrYwfXEi5uMx6hqczsjEvD4p2M6VyU8U3z06bZNYDm
y50d4dKMoV6okrwzc0Gi/Dd6u2C7S4OxpZWdxTmMwmKREAnmzRONhA2p6S4FB0lP
ROZ7nh5QOXhoy3yYt/J4Vxthl1YH/VbRWaTjkZ3ycP5j3mIrEUgQj8Ca8yoYwQ9I
AEpgt/1HypuO2irvbe9hLK3YlVcErjRrkGllMe8Fk0eVLs8JQyjyqsjmUh059L0L
GSISLklf/borj4pr0RvvHfBeFBXrly135PuS21ifPLnvc//4Y79Waknc0cA7UdNo
BMc9sMRR2K6ixisOblfN4Rxhuzxbl/gZM4R1lIOSc5Va8FKXiPQN5UZm0P1+N6tR
OTUTUr2myuLsF7PMKSRO7XreSZ7BWhEWnp7a+HTJYXe4sBGdjqrD2R0mGB9kdJMw
2ttMlURsARBYOPwX8sfI1UBi4sKMSrPryv//vKj340FSFXB6w5rM+DL5gIw/00/C
S30PK0wyt9aDzL9gUo1ZFKEEILYTW7F14hZg0J8fNnODvtcbz+ZtNqzMMv9T3OjG
6mg1SytLZd3Rv9vlWAX2cuBwYu1F9eDnbKgHaNsAtkzmMbPwOvtek7GAqb84R6mt
tQbLnafyPaw1q7Vj6NqCpPwaZ29BhmaK7sNfYldTdcz7TjvECvzksKzZnFZ9+YM/
RKyFui6tqnpqhi7HTlBAOFIYyt7hM5VeNhQSiAER03vj8AQ6IKNEaC14gUEmp0jN
NtXz96303+oZeBky/1xUQ6BQpiN+s5nKS5A0BTw0UPaKW4ELEkN25a/TSS8sHgbm
4ndn9lVL0wn3djPywYR00wJ4XOONn0d6t3U0h2ksSGeZBN7WasBk/jJK3xabdJNv
iML9lGDDflqWcdUCQhA7t2pbsQiiQEhL4ESKYxO5aOpQexyl25Xw81EMTyXZJkpH
zpNpxsGGGnwJe3uTVdxUvHolS/opsR0TgwaGIrtPU4SBcnHFZUwbqeOE59EgUUzf
Rz71ZuzX1tl2N1Q5hNEBRX2Vo47fhprrvmSNnvdUKO6EsBFt4KXFHHZCGPK650If
avxklMF/yDWnKMhnIlZoZFr75Zs8fvDUYOFOj/I8JBB5sHJQ84uSGHBJOwj38/GT
puG59M+RRqrVmbN6WS/KNq8fJ8VFcUAWjwNPYzpbyXIizUykFUJO9vqYWJxRecRg
Zt+aQKUokKIdI1WWxE0iy9Jrq+6rfcFyU+XioNJoSy6OLGp3jMoOd9phjBHhM8MG
YmqPzUsQX9cTorxQ7Gtxg/ITtTu6k+Al1732sD+odiypsjDIgEZRkJg3AuQ/k0yK
94D5oc1RvG4EtDrnjQSbtCtQf5Rhp5SsXCY7rCZeraNdQrPOOGUoM7a6wl0+bB2m
7lfMHCN2gNAmP2t4JPeB+grRmDGRaFE/zZxLHEXWUzbVCOQp0osNopJJ3nmjScls
HA6ePdgcEtAqRftw8CKTCAAO2yJPaw11AXE7q6o1Mb1b84sl2DiV1H/sVDmpaCoQ
rJsa+Xm2zTiwCP3Y+P8pkGig6qMRuhSQ2/vkQ1BQFloCj7zOBX5VpTQ1Z3tnqRTX
DFt2EIjYeSeuso0lhvWGG9eMizEIioOpcRHiAPpmS4QL1BMrB3Fj9zZgIkkIpBfa
SXpfMLP6BhuHQp4ElUhe/aalfPBb4BfVlWoGDOlSwbIHXpK7DHaGNCNiFnaOENI2
9ObEzdhOsm35BEqVgqnW2da0vaUUOcQz8j/cSewpRxXEldQRKhz3J6b6vdggSj9z
kwIWZhYQQKZ4NGTo6rIByKr5P5LBapMlTAaRgDO7350IN30CAH1RghqmAV6Z6Del
jiPQ2LUcdQrWNd+yeKVwbi+9Q6lFthcem7D1DigjoGJSx6EOMGNVinmcLbYNpmrZ
pUoWVSRI/hCyDnT5uO+JVcrAOc9//rbglXp1CmaqaKE8Md1NfTtN3uvsK9lS5TxI
hFWMUjVpoMJqgnYQa2fhQdw/bMSB6Guk83VLq/f+siPgjj/x/UprWaLRTyt8sTht
g6EcbViQ5RXQlVCUs+Wc5DZ8HRGBuRdq0bEtAz1WeES2ZpQ6a+vyl02F9Ge1n4WG
mvy/LXsamJynBsHZJv8LHcDGyLASyfdDHuNhIzh+rHJHQhKU63E4EQxcWLA9eSE5
jXV3ulDxntkVHz11b74uwZQdWaaD3aWC/8DAaAvKZMD81hssmutmK4gyNKadOi3y
9DBT11BpAOWqIA5wAKqcmUmyNCjWE240SaqXYCDJ7gPtFpdGF6VSukSSm5rGSelE
drDGHYxOnepTAKSAUx1Q1GQ5vhKRgc6leUqj6s3vC7Ah//sgaynb2BqbN59M6fl+
cf1pcFCODozPseL51kwXiEfg/gO8V6o8Z8utP+HRhnwY8oDeUUxso4tHyjBSrFvO
wg5JZ6J6A4dYABxot3RBsTZjBARdkEYnMMhCn85W4R3/egzzK+0QIEQh9aNHlSul
ZWRRqdMMGAiak40FrXfvo2zWPdE8hiUIMR3zpWDmdMxlZh9lepgllxYb94x98Iu7
iuV54YmYabiDj2UX1z99LDUn4ZPMuxqNHRlYj1NB+iQrOpg4MgA39U0rTKZoM7oP
pceiMB0leRlHXr+3DbPUapgbXB1ytfZjyyaNUd+fdBcwKcWGrO8zUplmQMGFzcFD
Ed851IoFuU0q5N/YiQAWo+1/KjbfFg8vISUA4LxAfeP/JjxoKGg8wp5JUtD2hVk3
h6oZrwj3EydUJ7UxppL4cnRCzEVc+taiw6+7Kwo4tfO7HhHa+R1jHIq/Q8Slm3fY
CpB1dIAVWvgZ2Mr5Zg6c9Vv7NlfSxLPh/+yjNInJABI3OGBvAUO0btFbdMUJ5k2Q
TiNdVDoAoltFV3Bkd94F2y/O+hnQMvKv0neHt5CHNa4//l0Jky0WCuWe1ZlV2koF
5fANZNrqTU9+MZLmXICVKgSj2SS+vLI3LG+YveneZZoQmsAvI4JpgQFyybX5ZdXl
QtSqIrA4Xd7yfGT/62L3vxXkNwFxF049AJ+zGSuqXivNHCOulFzqIpN7Dl/M4ZlA
Wx0DO6gTy6tbwenae8CSVxtii6EZGJlC1EasdKRTHc0qFJY+reqmyop+bYOZlAq3
HGZ2IUJ6BqQ0mProRpBoudzeXyAtTmbJA5g/KyNjve7MUHtSlf0ow7nSaIbXtKEb
b6nggXiHAIBKYQUx1ozO74jZcYkZiRa5NlGmEdpPepkASYqWVBEi8Xbbml/fMY5N
MfPFG/GbT7EX0tWAfbPZ+LP6dJr0CN7yEprR3+/QlkqIaggc83rxJ6LwmINmYcon
LbTuB8SktM04TyEW7bsTcoU7ultoGlGG6RCucOnOnoqaeLk3NF8ppAnsJOBP1ZLe
i4M6QTRXWo1XxgsGyN82y9hsQK41ASv3nPJkiU86AW7xpwr8m7qIheJ9B5hZ29ZN
yq26c/Lr0cCvYpCGZ3hme+9o2wYmZhE1zXG09CogJTIWL3ZvmqYqL785cIC2Sp+L
bK5QTrDBIGFzXl3lg0+cO1k4o++0pyI7tEa4E7OI5eoEokMfv7l9Z9z1cSu2gkL1
1hRZpfKnrCY5+5BCe2x99Mr5ucEhPndO5U55y7y4G5svLujJuwa+eqJGIBDh2Ydz
Vq9vyFo2mNjQLfJKee2s9SlEJ575//4Dz+InZnj77+NtRcsRArC+o7hU2w4qwdnA
4+dSSW/osgQ/mawZH2lOFwH51gvRb4Klwt2ye76DBZ7WMjLscmZnArpuf+/ugCyn
6RFzmpCA5VyGh/pIeDGFm9WDh2goPa/q0k0z9eGI1wr708q3g5baY4fNpZvK97QG
4yGUDTWjW+QSDFL1xE44TGia2l41zqBYk/6ffg0bJs02u3vukd9aJfh11vA3Wx9m
EZhBoP09f2aYZqQcMa0lMtsAi4VeJU0bbLylMMkTxcFDiijv+vwBUJjyx0HkhG1C
aNZ7bSaH3mJ2Ch1q3JZvAsuvxBrxiOOYSxy9TzKUtgth4nTaVM0XPuyGqh6iXxeO
eWUDhPVV4BXep88FMxL1Fg7wObkn3g6CL2bmt41Uen6Z26lEG0epyGXEHUkn59FO
P0odvcnDERr1lvZEK7097bHl6p/XLQXBkd31NbccQlwSc2iZ+CzzcuY5ZNWbN+AU
SEdlpi9NQaK6D9SV6NBiTqzkHRW2AHdFaS4/r989FUhGLEi1lyzEa6VC9Q9UGpaP
b1LCq59JwFhlzjUdpoDqjeDSdK8zFWRpjkARLScrRB66J/Rmk6uTJHBOEPW27eKC
zTvJMJL5FsalZ86p1dJ70eIA0HCVTjRjb9x0T7X15MlhEzxULeRfq7swnjXaoJ8I
RU4daGDWtGSalc5s6SCVwu1DjAeWOpexbiHAuoewqcfwVPs9tk82MVhrXF0/Njgi
A8xwGXcRXkBnKPYoFlojh8C6/seDG3gX8M5Lb0CGOOmiAt8X9cavGGK480gNEjaG
UFtl0QKTRc1O5pkMDGK9PyRdN+urxcQrp2SeGvN8ebK3y4Xlhj9OReMvyzDESK6j
Yy6k2ciPZip5xkHZM+ONQGzVrl9jqN0F8+0S9eTzrFf0PS6VLuxfyRmipGWvkdBt
KU09tAc7ChAiN1hoFvvOsRV1A6r/wZ8Rd7nJOBJF+8uXIawS6wbdquKBfp9Lflw0
BYr/qtQ3yDYMpxjCDzF1xWATbEGI/UHs6HtlJcxAetnWuHqyCTV7h7Q5TpXage4z
gsbvSPOyfiDryCPygvec4I/vbaJkfhMCZkxC95S8DvCwkmDxkh9a4nJtPFVeNtCc
dsbt3Psirn+8vqUvbc3k0HJJsQHQ2FF6L5HWgWcKHb/R1wqgKEvGzK6RgRMzegTp
mfF7+ZuHdb5hhwA4UyRFtcoypWm4yxc2P8MmVf+Vuwr8dluSVm2vXdOCqWXKRKKq
vLfbZYVNyW0/LQVSVsMFXXQW7EiIHH60+/4mhWVV5LN1WCJJelTERo8QoPXTcfV7
A64a5JtNdeHFxmjFg1sd1QfI8XbPefAyZttUrnQ/mbxGpnu1/irj7vWj3OpI+TL0
w5U3p6tFrVopyCw62VMMvaaD7v2DSIKubQK4nY4bmCPk2feUDH258BMfSmDQqJGK
sQjoIvCeUaHgg+IXYB5M+6I2N9ruKmjH06eUlthkQZ2TejBv0RWorp/J8L7x03TN
84H8g2klueQNlXpI5TMbdCBjmUxwUNq3ihlbdI8NJCtiNZ1PkNqqTvAWHZbdi0J3
oYk2IRk0DC8ksXB42XVRetzgGeeSgr7BNnjHCLzxMKZWIb4oVDoffFP5YkaUjr1q
xIRkUA2fnFK22L60FlAuZQLB1DMJvISMSRuKjse9DWubxw7auXD/bxH4fYMyta5J
3pb5YZ5kN+GkITbbSBHz0P+gDOQYaqV+mzJ0A5J13kPo+PhH4HKWi6323rZMVWh0
/BeSx9OLmCzzKe4r09gyw8x/6EsLpyRVKr2Ry8uruBytlorQaLvBl6Orpg0OB2l7
7dRW//JwkkdreR3WCiDLl+oOe7AsXsSKIraGhH9MO2MRf/WTUakI2mpi2OAZ0Gt9
f/aFsmJV2kRF5Kd6/y0ZIOZPq76C213h+3o+YN6lT2mANPirRJQeIPBA5xll9g34
GbGP5T0FVq4WI5alWZxbaZGVjUgIj0CY0khT9VrLA1pJieyrZhccmwe41LQof/is
T5wzOrBA5VitLbIrwE9gL7Az79H/DMgkHd1rZLlLF+KMCthiQzeMQMMe5wadlRZj
bdN3zXXDOBUt6WAONdcPK48RvfJAZc0QEakQ+wvYNM8lln6N0PIZ/Ceyhk1bcv13
MoFswwLlo7tPiRqAX/fVmBBDVwhEy/Gt55imeduspgbyjyPb8nQ7KQLMl/1T77CA
wbSrvnk+0fI/US67Y03TzMOVPf2JV5piw8h+OF8Fd1XHg+W8BBaVgqy1ORlGSsni
pMX2U9jsx3xl7J9mikpmK3+6xRYjJSTapV8Iv0Gz55B+Ihdb5taPkFqjxo2rvPgL
KIzz+k3Y8eNvm/sP4oueqZHtjbzbSTjxxdspj23rRDHLv8tjQvhjRlzD6C6ftzMT
s/aGuZgURiMc+c5qtgA4ExjijgzmzPMBOC0urTML9nZnSkGeUBcEup7ieKH8DYis
UKgyzexoB7www0p4DCbk32LbI1C+MralxX77YQPLu7aasPcathOFGNp+cW8AfBVu
H/r5Ka3v7hMsR9Iw1LzmIC9/BbTTfQXh5LuO9Z3m9ZKXqm2yspHmHaX0NPll2Rar
JOd9sFYHGUc5A1eqr7djtdjoxC4Hl4Viv1w8StxltnE1wIYXDt/kCn7iX/N55M0t
UXpLP6pmt3IoIFm8EoYuTSSaK1mVtylSmGwlgcY63/Ku4HQzH0HDhOBoW1HMkL8q
2OrAzfKJtx9Aq/IzGzoBZKqTK9lFtlsx5p3H15gjAk3rLpr5+CxVyGsoXlg2vCRK
q+KyAixx2kh82unW0Sv/bM7tGqpaVxGtYM+GZOrqgiDSuW/Bp4+8LsvYRdcVNsnJ
FqF96fGNMYfohcxXkfUdLA1tfs7Z8NhCZ0nZtjephKLbN/oLixUmPn0VUGAMmiTK
sgzDDapupvFeqGlsx7Gg6vbQEcmG/uFEuYhncVEGDftlcT2QWmqT7DWoUxNI5a2t
DtaAITN2H/GLNSVFdL/TOzUwTOx+2scRehKB78bu0u4L+Dmt/mwL/EE2K/UPGNpr
ENznS+WRN0OS3URH45Dxu2UAppErQZodD9f5xlKJCSAvaWdNaORK4Y8DwrMpbXdo
CAxu0Y1rHnYJEoquZbNl2a4WTCQeYsWY0e+9Dpgz+8FsIgUfVG6tSGdTDbGdgyMP
vO/2SGYlOH5sMA+XQhAx9/R1SbL4oMRbgcuJ76CfoKe9yVl2Jei0jHsL1sU7v0Do
NbfUornZkKw2OACbbALPU6l84zSlBJJSY2ymwRe20pNqyxszRIhT6HG8E/DBlGGh
rdQF3nKFnsrPBZsy3OGABWB+gGNGWXSzh5cs2drv+XRj+oZu248NfuX5XwzBpWsj
q8hnv89woly/IDAcG8OVA0Z9NKhAk6Y5QljDP1E2F+ajjyDI83ixVjxQq9q3/CDY
j33bMFHChPZUIjMutS8jvrcdSG4yUFVv0muD0ig0kdCHn0Ua2Dzfp+87FoLffJ90
FSJ0n9KGT4IxD5Qd5/wMddPxy5KH8XhOMa1AXiUj/VRxnOyivfAJyQypzpRYQD/C
oBSgxjVdzjDjK5OmTkizMzQVed6CWth8E7p01QRSNebixaGkq31lcfOVIkhOCQ5i
qlnuL5sHfvwxJDoQZl18ijysjy+jNlmddRTL71Ea/QrAmKG63d+TFtzOoU0RHjjh
8YLaJJFTWtuqEZbplGMrWnMoZpcfVKBgAnuGzt/w4U38Fe3m/Rh/v5McRaWCJhv7
iwsv+BxpPIYQeXUFJHhWsq+bHt1193F6L6NwNRSglZmN8k4a5QFN7vaWxAsb3F0d
/+GA5paTPoQDH0g58K2Ak+2Gkxrid/e4D3WMpkjHMuseTjvQgv9HphflaMRZ1eHz
vREisGHyEDcEdg1JFdTqYFFBmThvQPUjKDwu1RgylrdIYkrooVV1WgAxfjTDLC6g
dPD+YYM4FGRY6vSgqa93Hu2O08yo54tTfxln9R1kozgcJUuKv6/8rh38sVShJ88a
w/LTpvdlbcsY3Hnu0uBVYE0RksGnok9zzCB15Nag1X1mzXfdw7jyOd97Vzj6fLuI
qcmQyqQcS5D/imWrBJxYYX0ZzDGNC4ukYIBtqAwveMk/XdI8aA74GZ7YIG1VN/7M
K0rKjRCLAMwh/6Yqs0BFSiLagXzRDdGyu6RYM0pD9x49bz7K2YZZnQ5iKGwVBxgy
lMM56uRZtMdyxLZ4xjq4lrqYsox6K5uMM/bXfma6+NTEdEkdu4XOlAfcA7+NDHIk
k6iUnGcZI/SGKhPVPMV/J+ulh8GlZIuBce7khps2Sl9ktbSDqaNeFuGxHyhbQsgL
S8MKSPocOBpdmSqYbv5AJaJJVoiS9/2qFu4hbJqPB75arAq7zN44/svebKZwTeO8
UhHaUOQh0xlrGKOB0dP0mkIq9r1WpV+aYvdsUDL73CBKcaYwGPzDAek3xThLiXxq
5mabuHz34+2ljSxWwBwUaS3ymof4etl8M9yaC+2qO5ZDo3UIKTp5+riQWY7A8yr3
6o3/XnxizU0DhvOrLsjtzBZjVUS8mdH7YNu7WP8d3dx3c5V/gHG9qXOXxZp9MUTY
kEevhv6A/RtLZF+cnXxW7O5NMqSNi4oo9sIM2Foov+Gta4Le4RERYqm+kVQgyjnq
4Q/egLDK5+ZWNAMofykbNLqodjfTWlU9+cWKTM+RPrSZBjBoR3Y/NIF7dJ5NF/OU
6ql0BydI/5Nu8hBp/vA07uNBi+BzJj0Fq4QFrMKuSkrx0shRrBz605kzkDHaEiA2
Qd5KA3u0YMMyX/EFYMjAEaQFFNqSNWUTnq6Kr7ECI+8M6Mtd68HsBKy8gly9rTNA
/V0QOuEYUyYC3N8jQw1rlZ4wmYSXELkBQnxLs1MAnWnw7V5JAaYN2d/hf4x9iJ1D
SQlvT3LMw+LnAquPMRSoS5gGPk3/f5zScAZv3Rp6kw0efEzkZRHWI0yOyj4BuzUm
kra0+4CmxtWQpdOCDWIM7sHq4pNPE82JjmJh53/MXzyJuz7vSzJ0PZhUC9HZU1Bw
pTpqaCoJDj7yamZWpWqwWZEcvlaF/sItS1hBPm0rCTVxHcQYRe5XOd1KRV9bb5VW
GhwiWA3ZS55iwgJVBD1n2V4PAdZrkbiKDR/MQlhC0eoEZ7ysUgmtnuix4D0PV4Oh
PuQhWDKoYy6nhOSM3bQUXUuzQfefVN1rqVKVFbq/o/Q6DAbt9RBGzo8YDh9Li50X
0bmPIoqCx5q6ro5g5xAq4V0P4iVMjFrR5DKPQjkExeKtWS7KOuPSX95LeEJkyY8X
M8xsoMX4W3ba7mj802sVdmZaVjDz9u1bxR8CrjoUnwtbdvkPnk192OmbcLQXgWW4
0b2zDLRVjmyIXvzmTdiPvP9KJbHLvTphHX7TgHvxkL83gvT0ULaNrdYJjXPwsYeX
o8tcoUDObUPb+z9qINbetr5eXAF1wdRgjesTJeI3APNxD7nQtg9rDJTMSQ9k22aY
JXTpwwt0Y+0RSH89bB20Tw7UQQoNGzZaWU3XsrThEcnvSDDzf0RjrMM7IzXdUaHo
AYRd7gcjk7HCmjj3ZRUJda1eh0NWjBQ0K+c/VzRyCA8R50CzfmskRf8wc1la2oj+
ng4SKnVsSEo6VY9MU9uK89SGIx44lcIs0Df1usa66R4ncSv10z4mwBYl9loO/Cbf
BpCmQ/k+6ZkOmYW7uXgosKaSd3wLyDERNrjTtchE3nKa5I+s/CMTgQPLy5yRiSfZ
2ikQonxdRt64yonEAc6gFn0MSavbORCMyR08D8vk+9q2Wsd/bUCvjda79S22Ewvd
uafdUus9Hmw6zlT5zduamktp5jmv4cZq4YrPZVm/IhdCTfgF0MmvPYtPkp07SS15
LZlY4Ko9N9YC1aLu7IJCa++rmBfVpE9LPjOFOrw1Vh/GDSha6jrEBtksq/SoNfIM
HtR5UlYisovDqZFat+M12Y9nUc039mgzgIFLEOvx28TrwmSIx+OXBpmY/Zm/AXHx
yAXFpYvJDVmjtOKoCZ0P4wrKILyp9LSt1WiCbfYV40VuwG81EfuCajH0NebSjFLy
ebkuaO4X2SwsLMxHbl63MMCiJfyh0wOdHQwcx1qI54cQQQkA0aGoKcszeQUO0ULC
NQS/YIKFDgoxLRIhUkLYg9WOjckrv6NalCERGUwuBZv4lu5jAig+D5wXBe9HGr2O
sdcRdESkQiiE3jRAAT+pS2B857Iv1kUQaVBWWcd+IVcbTVN4gofOIOC58V+SD5II
9tRSDBu3D6Z6UUOL80dQclR8JzHUodpCEu/mktMEYVduwhccdstQce2lPsKPuHId
opFd2OyqXjNC9CReJdatAkOtV6/hdPMRI4KTWS8KWucKX9fbd1fuoEDpq56laGME
6KW8MhmwsMGiiFnLweW1rNYbGfn+gg/qzixRIu/RQ1tmgFlcfZ28r0pyuBpePO/K
iHcEyS4XU72f/Mr5xZI7jL0yMUpPGscJEUrxSDaRxmrDMjplcXBi34+VbyHafe3l
jADfjYPL0lS7foGomrAZSZBNUeS0DXWMfg5US9qAHnn85wuxKz48MT0ODZQqAh+G
8YfAZS0KOFpnRP0azAUqSOgd6wMIHWex2zMKYooaQC7AHWAZNy2/pYI+HaTd89dk
B0S1LIXKdnWAhOD+uPPkkgbBW0E9RnlvakDZbbmxw3tN39xRg1lqdtJUKeDK3kbo
pzC3CU7Qc29Sn+jDeB87iLxmSL6NnHg05s4PUT9QwrnaEim+4zqkplsKhlMsmfIc
RCFYwH1p7owUL8GI3nebImykPHfSKEEvtx3rRaQo7fSlLRR5nxT1GXRS3pjZ+TM9
a2h0Q2qRIoLPU9kppZi+qmM5p23zLUtdQusdz6jr6DeUj1++t95+NvFuYk4sDCMY
m6uwRhdemOi2NAc+9OWTx2D3ah+/471+eDIsloE//m8bg+0ErpbIWjiaiFLQ5gZ8
dRPZWbhHdessujrzs+DXVDKPhaXxmFqR13rupXx8ogp8bJHWley4gu8743Kycsyg
1Wpo/5Pyf2ppIl1iO3vszMa41By36E6fmub+wFju/XDsgmo96ys55BL7gFfwb2UC
j1wYskyj1+uz4EPoosVkpanuBqAHEtfLxPT+afbUhAfLJqk7/qo0WxM+LARH2CdE
01rf5Srw3vKBkElJN697+lye0DnJWPkxmG7ExpBbXXD7/n+/K6ZxPGxb2Tn6VThf
tqBOVuvkTePSgBfhnM2Zzt1A/jFCmO5ZpQ25mfCnzXg/q4mIEdlbw0LTFtEv/aQJ
i9v6k3Ro7tWaIeX3mg9QvOoD+6J8ZVnv3sa5pTciG3CLfiIC3MValK8PeMYpgVzA
3efZrk6qCeRrn7HpOvvI+QJuMMW8aGutq7yzfzmqY28YgfnuqFNM+06e62u/FPTu
mMllkpTmPClOuw5ACvXCnTFpqMf7GVWxK52tZZnZ42v/5tYbaiUgVkP+E62v10g5
YEoRwa+6yo1psfk6BgaJQwGRc4+FUxncrcHg6U8EiGD4EUr3/mDTVO8AluKuPWFT
ZnlM+gnEVymtd9A+4eY2/KESdqzzACJiJUCTh6r/iw5YMh77/JV+PIWNMmJw7zFX
8gSrdYdZwJbdto3pPZ+3Tm1kB4UNCDZFY9Mc0gyVkouoZiIeEq20/19fNJxVVo1B
qQQKudJ2Lmj9k/OIwkVQp5Xzb70VqRHCkWn5OeRd4J/qHSyQnoyYaelJUOJbK0JY
+WWK1GyX1ABTyeoU6Z5ZG+2iZcXTZuEW74+9IkmmaADDwx04P6fdhUne2pJm+KvA
5IT7upJQxdSSbzEQ4+aYzM32mJwPkwFskDG9Nx97JJ5H11x0A6O0juPngq8grsf/
sbgP77ugdI56UL3yfIZAHw8sEuKodzXrYwBNuLllp+aqqe/I/VFjWPMWb/GFw5l5
cSrXf9/nUqkPpw/nwgDHef3bfUJ8X1I7Ck5uuBf9iSwWAqZHbx/geIVqki+whh9B
ao3HgKM+IJ20Udvmbl/sXkVwuJUXtzrbCXHtTpHQqXY81AvfRFlTm+7c1JF2h2Zl
hSJbalU5NgRuoRqmGCc1HoznytGvbztbrdbAFzRBvCYp7B5VMth1UNmS7dyW0F1E
ifMSAZ9ISF68NfQ7WhTkPisKBN1WBEddnyR/e1Zbzwh4Hp8G+MOPWe9U8BeJLJlM
MdzKCpo1SVYcyzyW8ydME6WRCwL322xbzUg8WJVDZvkqScndrZNwr+wrAjVr9pAi
h+BTtE16u1KRdG0xO/h56MHFD7sYeW7PCbnEEp/99hEuLhvCZY4lwwt+hw6jCPRW
ayHIukpe835xOTrvNFTpg7cOLUKME3RmWWnvx6HR8LI3D3KbOYfE1FWx6NwIc+ry
fcip3Jji6hxR/rpD3OSmAOs6zu5yLXSvBtLm/xUB9nT3FFegpcIJp0Dl3zb/KQpG
K8VpvqBTA6enU5Jfb/O7nBB9j0w+cyIM96sdDujSrd08489bVyF4vK+Po9Cbe83p
sSOu/+o0svBkDtkoHb7D8n8o1aQ6E1P0bFR9piz8aMNW42D9KRUybJMJt1XfO7FR
oa0uRhXwiVIexZkfxQhIJ6MfrjS+rkjIeBx9To9fZunf5k9H91Ri2IWtrnZF66XP
U9TN9oOV8UVEVOffQEYLQEqkSWO7SjXNqfzkjfpu+n3GWUz9NcDkEd13QW2QEJQO
0V/Dt3Nu8bm0/nngqxpJtawPybLNtO9UhAdCXjmM9ZCBPVaXn/9X7h6YvxkzfJDr
eAAXN+LdxyBO3lbjh7OFA5uXcsPL3xzRV4bC4GnBFAIaDWmu1YskkNOP8f6M1In3
fdljMJ+voQU1ZVYrMzeDh8VTegDy2I9kI4x5ZMpbMx3o3XMCv0pDwPvmDs8mCXOM
ahXkIHtWQ0xXhGwS2AAITeh0d8HbyE4n7cn6mtJs6Z+rMdpj5LH/+2E9PumCtbbH
03c1808L6AE97RGx0ly5T0pXkNX/VHa1GH2934Awzmnw/QpyYVYL85p4WqtEo2iA
L/hEx/5dX64TQ7Tzm0YCXOLyAhWjTAeJ+pJErXiq4elsunHOqYao1bDFDJmJZ+r/
Yl+Ky+lfLA6j1uLQW1cSyUGycZb6nN0XogstXyr5QIUbmONy+W8Wt3jN4JBPy/Gf
P7wbm47BTN6SjXqBa3X56f6u+8oEdz5ga80G4ujD5Uy4ldJ1iyzEhdZiO5IBiBZv
aWOeCQV1yw6A+UnCT6npm4AA1Ni0eyH2JtSDmWdcNYz4+cg2AibGybl/HYoZ5fzA
EGdT+zVgZk9/RGSEl5gDgDDXUZ6uftybflbKf/ajRVUJDDYtM0Bo9AZOQTmn/W7y
ZvAQtN/76smMhWbJAm+eE7suMrM8x8Ib7UUEDcluAFjsO5KwGanfegqe3LoxLUJr
p082D4oTUxPk0X/K9YahqF3hW04kv8Qpkfdz2YddUcfSmOkhd8khKIIip5CqXuam
UFo30gvPEI6HouU66Ezwu0h1Ve8eAlv01M+YC5Nd7YRQ6g5QIEqsFnBFSctqqtiF
1DcLIvebGWwdZPpcvpAEFRDf8j6cq+5txtp+CEzE4JJPgnQMzD66BVu+ycBE1xhd
aS9xAOStL2y0KHUm9TktcWxNjgLt/2oFjEDyxuYLcTwY3UlqsD0KxIRyD9tEjBY+
ZGVVJIXQmrCturx6/DidpO2Jbpy8+zjzVD5tW1uCGFsE610Q4yv/lcl3famLe/eF
h+KfKZexmrPzwGMRvdSnuV9bCtlR4d825/TpOH1lr38J9CzWSlDq/9Oj4eNKDT1g
/+4MNtQj4SVwo4qPQbH+ZD6WctTBOFt/9mKatm6MkqjmdkS1I8L+gkhLSzfCMG0t
0hX05F93kdKpHDO/yyoDnuvky1JRh7gwvj4/hltevNeVje9BHy3LK4zFu0NDLpPp
Sc58g+i0Taff6+w38JrRXt5zyvyookPNAUC1HtNnS/lUWGz4xqPO/hZfEZ0EEidK
R0LJ4kcEIIGwiUoX92+sFqN+D1WBH1eLOlPxSZthpQhgKLaFLqhHqpg0T8citiD/
9s2vK0wui1rXXZrDCgyCjWkLAJh92V4LDjkYjcV4xYcZk1KQMY/nREL9yV1VEyyD
wJv05hYNpbkL2UyJmcqZT9aK5RkcMcK/lypWhI1ckqbfyISEUrsbeuNMt0pCSPLa
yrxQ41isBvuclWzc7I5Ex+wJK4hNK4JWR/U/Wgy4An1JFQ/xnbOVvDVPYdLVBGRz
BOZCJflHW9azP55EXomG6sCLbGtbdYCXUkL+ZZBO7X6CR5A5afnmzZSpOgH+rSjg
3zhGAPvQ0ujqgxBltj09TE17Qn1VWU2wD1E3xw4QFcLTvqBVzlc6C7j4wgg5Kwp1
HCx6vdgqp6ldbfjn1UQ/MqlPMEzwpWs+aHv34P3KOI3FMEzH+tkyrZVvr0IwU3sr
riS8ZmOCZPhQEci+4X+dcweTu2fQTY+f6alXHOfsrLzv8WRrbydnduGSoJzAq/km
WBUGnD3awztD8jO+orEg+Pqh9bljLFyrERpeLCoL7GllTdOcTu3QN9jtZcqd6Gyg
bVCqLF4gCnhsiXD6CAbtpGQdUR4xkqaJqwqvqfFv4ARIsPUPTqHBUSFu0/wg47Qm
BBdvvizeEjwqezFRkgkGFX3OQVOxeZ2xmbACo1Q4TNfrDya2T746xhoWCO8PTNkl
R2Cxr7B4/p5PDKNJ/phePbMk53acqPp/H0picGYCRcOrJ7T+ICkbiT1SF0eZ5yor
DgHuKbdpFSj4NP4qvJP3CJr8ww0SPAVM07cfBZHetboVSduroAsP/r7729vxDDTG
WrVAkuQOuzpOLoJeuPHGRNqtz0Ihevii1aeGf8aZ3/HmwRq8ijBrw6gL0qaTLvq2
budF1NocAMyYfQwWQ5/fHraUb8+oxu76gUFV4hBv+0DZmAZePJXFf+Nbrc6SOJbj
2fDyJI5U1U+p33T/A6BNAIrCMkAySM/pouGDasnNrl2Fvw3bYn8k+vwuNpT3UL69
WN7TpWqLZmW6nwz/YneJ0rP+DH7+Q1Zk3RW4rx8c14SUeFCWC6dRC02wL+9GOHgY
ZqnG/t6QcdKeyuPWw27AqKpv8aZU+nA9AR/3lCoYtk3lJvPx9R8jMlKg/D06JMyd
GV9F469cS9od4s8X5h+Lrq2/+OG2cGTIPUWINSJuX3AR1HNl0c/piQl4KoA8oCom
A15S9Cdz7MKlJ/XyYZ5uq0B3PRsce0I5azqE143HPBdsRAfyClhH7STN3ZIeYh74
pPE3e6PDvyRIYJKxiaYoqbNdoxK5/qkwPBFr2zAFa7yOjtHv2ALzgdEMEmNcgxg2
sOhu2kIjaPHoDnRCGqEFxr5qWrTSwIKBXriay/upSrboDZTJNLSdyQas0MqbvJpn
+dHzP/ZQG9/Cgb23Uy1kjZQLLIH3oZPrUq/a9gdLCOnEdJPNw8/V8n8pd7m0AhE7
uwut345F+sYAIcCwXTQMqKbgoe2uz1PJf9BDqxdWCr09SBiZUD0QFUXlWXoS41gc
mm2XZ3dutfHsm3HAeJbvKgNwJCSG97hjRj1HDzAkZOLXtOGtFtVNiDd7OrxIZ5m3
JY+V2r3Rq2GChz9RCBb6HHAkiTW5t5oghyyf9toBfNIrLeg0qTrhWEBA3xcSakgo
gmTthc4wLoiR43/1VmrKPeXDxzMsrRxd4tLoY7zfIScJsdizLnGvc3JL+ddy3ni5
QgT1caJZjhd4PMs4WWCflAYXKKXJ6hYpmG/AKnTL/VdnZ8ZaW3dxjP/YMs4+5+Fo
ZbtgG/v643fIqNbOptEn+xkJSPhzeMwlDnnkpjPGSvzWu0gyc/LqB0GxBFQHRgc5
pZ++C6D5C41H4hqKK6is1//5zsEQs05ztpgbk9rys05W5fO8Ip+SefZK18s8/mKo
HvMGwGpPbucxP7r7kGQ2SeXKlrN3IfpHn1hF26yxe7j9E4Xp1o7RnAlZviRQ8jfJ
hitBsshQ+v1NXf9Nj5xPpxDxjrtSmcq4GuRUBJrsz5UQeEflzjWZsRsj2sK9r6U+
ZbEZOOazp52aOWmG9T1RvN8yf9r1dS7X8WJ56XFQ/L52HL65XRLiy1uHpsa+X0ge
Wzv61btM01CtuF85gWKwr46i0N3w4NIPiXJ+mF3RMpE1jjAmA3PBF7f4U8njW64s
xxVGmSrQmLR98o5MQwMNd8WWoFPTEshZpKirJoe4H6bHdTEOXTZ+igT1aKJxbjx2
/TR2ylnCcIZsqi6ly0Vx8A1gawqfcCkojxFrJET1PBukyAdGlXWmPws+12AONVGq
JAUpxOb44yiHCX7ZiKgajU6+kJvhne93DCT8TuTobkWAA2/OVRsq9ENGR6sjwZYA
hC2f409WYgxrsPct9PL2DcLuAlEynlRzqqnN+RIQuaGeYmGbeuhQGTQWO4knEJbJ
1tBjpbdHMZVOJFJBfbgiqcS9L5/L8DE6qTkJuUOrrU2eiXzHjdG3L0tb1PK+bqZV
92DGY1QDSlcs8x45LETavcfLqvJLaSiBkXJQVOvjkm+LFS8yEqUhWTq9rvvTyF8m
RGjjJdHuyK978gFORkmBLoChXVJRufWMno7w4bfvbMJW+Z9ARjGvp4Ggf8et7pdQ
bKHNuwlBt5r7L4qNH7dv83+LajxLzuWi6hz+zTVv4oHcxsdevfw56Omj7qdVXyNG
bcMH0U2yMivihGOK68i5kZx4hYrys+zLuB+1hYynnLW4vyRbV76PcBCRaSr+xQFG
HsawmF39SmBfAxBDBiMgYCG5kS93t36xS5vBhEyFW3JloJMcFtfG7+OKIQJK695v
V813Asc+FnN7D+xuKcv76ARj6D2evnjb0p8nvZ0k2fSLE905NrmcGg/GQVBs4LcE
vcyVoj/0HhIQbEVLh+NHhCsxAmQIcUiDSJlW3BJcn+Efi2I+FbWZPVv66j11qpw2
DK+B4nvJkDWhK1jrewK0+m6LCHHJ6vjR8QyD2ArSGVP8qqdmjjqqMbLtVSWBghth
sy2csCeCet/LcKhVzKaDPNlxXyCTNew7v4gPa2V3yDl8E/R6fQ/CrkrMW3HYMnVV
htw0CJvIoDYEHcQIazN8OBi6H1fwiUpSzPA5/07fbGCDFRSGhv1BGglIw3z1vX8/
xeY1nZZNI7xzBFawEzfMSMcJJ1Q2vePQgCP59x55sJxn9vIlYs4Gh6u8TFlqdlHW
5IMC1/2fHhZ9W1O5GBJHXZFdV7+lU3xaKE8buuU7vdhGJrZavzGoQZpw5yNUBBws
Fszx6PkPjDu/WPy41BIS98CRFT8hFg/U/ZIIg+++FvF9H4l1OED4PQf5VEiK/8SG
Y8Jnr+wR59RnIcnHzmfvrJpdE3rI5UhA16Kt64ORBB9syP/UdRyyY5pfMh+GplZy
EtPb03L6tPiFtTuko2daGPuWSqe6MfeRQi7kBJo0QA0d1M837G5+/Q3yjlcQCvDV
KtaQkP2ABq4yJ49vp1rO6PV5/mT27MIoq/vDV7Qa4p/dDxXuhE6baxmoCfowl4zm
Fri+pd42yCEtu2kcTNUhkekWsxHz+URZEEeAe86oyAQl4jJskGgRdD1FfITfgd9R
7rvN/9ER07ntAQpwlMsiRcoX7FZipBEMJBj6mn2ftk2IsaZUdOVynCTxgJS/bxTS
35UgKzau8Q6YLUWumHKMrBtghtirpAf/xw+kjImCIsoIvCbhfKWrenxkYovs3FgS
7/i1GtP1CwMSBsu+Fv3QD7EOnRQ0TshYrJeQgnScUXGba5V1H8aIAsjsvRvV1UNC
WbI0O793J9dXr1UuVlrd/C/cMXIgIyxmgHlYDcBxpr+iSJIFyEwePWeQo2ZQBD8O
CmfZYm14lgZ45tsWj+q/EzB17X89j3ZFZZaZO6oVAkLiMxBZFfbOs7TwEi8DfnJc
gtbPRtH54rI1l7ycNkCupTXqcH13ay4jU0sPnXT9pUwLH2gcrZrJvdep7VhZ0gTk
32tvsQoII5dKGD6P3JfOYiMkuMhXIOd60QrTJiFT8L9U+B6c25ywOrrONoUBSs+Z
9POcECJ1I9tOMySsHAqhkD7Eu9m+R3eddyblxycKoXg6Rhoj2BGTP6HtwMEMGCcs
xxIEDaNy2Nndp8qCt4lOyVnwYylB1wIip1/NkCHQymSk3rZDmX5nt0hvUIqCkWbV
HivQR0CYD1KhXfg+iNAWoJ/O+BXJu6ndetISjRj3V1LkmGPf8Ospzn6uKeEmei5T
ndppJqHfk1OSFh6uXCxtmeuNUvJj3hksf6uOve5Gra29GC8pWL+c5b4BWKOtu06s
lTi1AZkqI+PYCijuHt+W7ZFxDJEpc/olzDiLA3V4aqW6Huw3583RMIT7G0aL666d
f8YWzsbGUi3j/l6WWqZk2kRgKHSUSnoD1XrfFJ5KwIQEIlEne5S9/auA3qUu8iuo
ZuOhbCUkdg5Z2YYXdNbfmbkRg7SYcHfMJN5v8cHI659fcnXSLrvj//x348+L7kf7
mAWy0K2yH0BigEb4nI+JTSSQY/1iIlZEfqJPqRwGoRtH9NhKYgOawtUR7ZUdq7rs
fcTQsiLlZwLQp/KtVBAXuy1Gi9Y/1D0d4lLlgEVrtqYhlGY/bNYd4JdmFDTyT+Xo
w/my09fG+mN3o4I/reiQ5rUpmwR2/7S4cWGeigFNzc2nQvzocrBKDWOOVfX/FnY4
rGMdMHIL7Lp4vQTnPvNHr6iFeWFuzUHlbPIPcV3Vn9ymqb7yc002sfSEmoxA8ZHS
FDsXEIG5s7h5NJtrzTQxVWu2fDmmmLCi4CqHjyqV2nGhPcPuUDMt0p9ewRHQWtmv
6cYpqnag6xzToGq9a91fnLbBjh3zwG8NYkgR0PBFCDRvwi5Psza8t5+Tv84Ur2mC
HDrDu5+qlPZNGUpwyeBDDz0EDLTMHZu3yReEklqyhcmaJR9p58h79twLkahXY/Pn
cDc9y7cBUjZhnKA7gUiGOCsz0DWs/uFjUr9fxJwfUvnQt979k5T4At9ESdBBhDp2
n+ArvcFwQzTYxtgTBALp/Z+qcDOX6iTVXTxXmbdwuC7duyaXqRLYfTSW9JoeyEuz
mZ/z6LViSU7YdYMLcaJcQXkGn9YM2tLXuBiHS56SzVPyLPPH+YciMhjoH5UhQgEq
iL/S4ie6bCc7CeOoXby6b7eOoxR28uZNh14v+5O7i6LVdlXOzP9nV2QvztGFxnir
94wELeOIFfErI7D3so1iDKzJWpqDtNcap1Z2HCSDWe/35vNlK4wY/vrZ4y3pHmfq
VvLadJKigfeq2q8qAWFZv7grTvoit93Oy4GIm/N55SXSa6k66EKESwJvPiiKeiAJ
7RmAWWoJiVCCtmSbgn4MD8Tb1Z+m91xvfM7c6kEKQOVy3qMP9MXr7AggyCf38Yf7
Y0aJfbzLLg2nJ+4RtOH0IYeml0auLYpfRJk0UtX0Y2dLI41FtIoiXkuCl7cpoHyN
MbIppOdvGf7PIWkcg6WG7BY0+HnXN9ZW/+2TjeDcrWsvfbzxy1heEoHpVsZHllwX
7t1lwXKdTbtxNZfy26O3arAz2H5HN2jUAB3RYmmkpYiK71XeNCaC64qWnmIcy610
hqp1muK6odcpCgINv7sayV4c7SoOyZUk0HP46+fMUlNoq9Gjw697UIMiK7Qq7a3+
NMn129xnFfa/u/ZMdo5mMdGG0FUZtOmuyDQdtxdLMclrmc3T245cdiflZOSfa624
s90r6XhpE/r1FuB0zbiT5A+OZPvaKBHUe7CFzFidQlm7jtDIW1nVMfsjkDg7EHoa
KdS1hjmB98ycQCRKk86cGzUyAljMlhtdnuXLsF9aNjss3LMumC1fLT22QK5jtZLD
Q/VrmjeVYJue6QetJF1Rt6M3qmhvagNhLS5Y08ZUpKfKFLTQi3BJIxWq7vttSqzi
193UBEY0hIou7C7okdRSIP/0da0mwbhgqvkzX7tRM6DhPF8QJq3kZyuFv6gWLoAn
XS5ZI0Lr/qwgZEwsOw1I0dXanxaRob/w1+07H998JtPTXzHmhroVAlAxQE/MPag4
4mlUkQPFHTL6BgvfzTQiX5RNXRCd8ycqbF8vmO6SRenmt8u8JRMSnl5Am5ht80Wa
x86t7eizerYKTuXYcOzET1ZP4qaJlv3jbAuMLXZcIrKhLo7StiU941qFDLaOMq0s
yzMe0JeKoJbbCSz+VMKPNfuhfkS/wdJYgvmL54hhGtoH4e/++rFxj1OuKFa7Wx3q
JROn5NsjDaNPP/7KzzYATiaIwIh7bfiK9W2i2bSIMtT6ufj2ZiXNGobTzPDXg2uC
bpTFGVLhBxX0x/xYZ8m1TRhh6fx7EWBxwwRMxNKr6HPqLDwjg4HVWGLPxcD4g+oA
HIhSDi/A6jNoKeIjER39VCOSw8DnSoR9tFjR7tsAWzWK7v9VL+gv/49Sz5jpaaTE
NvW0OkZXi4Z6qcYCwkUveSc0ilTl+gxC27mwxDJmWcOUpv5lfKuzAIWYiGEjVOSC
MtiLdnWzpMwCgLtbIScxbt2VVrJ9IqWDg4UB9f7oaKol/XjjE1+KxsO6vIyI6V+f
ZoURnQATI71ULGQEZCflhdnIspu2bI1jgSAhb41lV8X/Y/mWviEl3MH9Lpp2UwFL
V5qlDleG1HooALYQYfXN1PlI4nQeMrMF6kRHSUZM3MHl+TrMnKBEmuBLorBsZ5wb
o5ceRKrodTWHAWQ+YrnluXZ9t27vuic9YOs4txPE0gqwksQ/4SyBtdATgMLCAvtM
3YwKMsLp8W8JbLImzTS+2DawG7DKxsdtCe8XmQAA4mzj64arrzMt5mJKfbqGaRjB
IxdNbSb0HtvrG6OwcKVmR1QH+L9IN8wj7h9HNvAXAyGufgmjr0+SS8n5M8gZkscG
06wYy+9hl8FstLylh99i8eqkCD2u2P/3g9zTib0xPkef5pbR52lxTyQCV4b+4+gu
K7rLgm1M5/hUbBfOQspXDujsNFBr4SqXJII+fcr5jCxYBE2rHZdfAvrbZJ1T3+E/
HOuLeKn+jxlVQ7+Oehjka9WQwW3WklDGg9hUueeNk42vZbUCLj0fFCpM87X21JIG
wtTgcSpzCISS9BN8fMt9wtRROKalBRHWEVKp1kflHlbrDwFMb7YUaysjWoN/Y5df
Pub+ZQITRkZ2fDWZXbNsbA9S2D38pq99c0r3FAPlLaGHEBQfy0zvNq5b5YXwWgoQ
QWB0xf5IGykK77yor5gQ3rQI8noNmtq/8mw+Nj0bDkHLaO1GErXPjSo60jrdG8uj
auA8rDPd4wJmsjwEPaQdNFXrshflifwxBYDkJ3Q4pbk08gO5xuYNAn6h0oXZfKF1
gm83PtIZ/qxXMffOPgJpp760YcTBT1ty8mTkivjZnvIgnIB8xBNmXJ9yzZvBx+O+
FYVC8Jo5Z3KpTLlVBNg9hgu9Y2uKQmTe1sc3ka4tGq0MpMjzNUnnZ+47zkLdlOJk
aH3kTAHRdnQPDFeyjhkMmvBTN5HpcoLMRtoHz82uTWwZT856KmcnzqncOrqVShSD
hKUtsh0A/hrP+ryWepwPWPRfTyEyIaFxjVPCyvqaA8k2NmGRvOzy6c9NdqWuX1Wi
8vy93Yu9uYYB48G13PpFRx3SMgZprz0Chcmkoai22iXZ4JmlXeTi0V6rSopt28OV
4fm/QbRQLQhz3w8qLjwoRZH3DeHXj9qmaj0+tssTOAPxN7WANQM6XyDXbFyO5qB4
sqfXjEmTHB8KNuL/ZGEdRQKMZnn1vV6C/W0AdGrdtGhHuCPp3wh5WHSeCrGZBbsp
M87g9d/JjLUwrjgc/5Oyil6g3P/5QR2LsgjuG0E+9iDPBOVbAQV7qPwWi61z7jvf
wgMDtHHq+SsuCQKrB8M6j/z2gPyeE2Pc9lGXPkS8lx0hY3spQ4eB6dcDOUJ+iHx4
ddpIQxPEYuYlRNlw5g4uWY3Eu7XBTeI2rIqczSgly2XY45evTRvE/ujF/q5zFSZZ
DcWy+eKuMi2+rhfU4SyZc9obEqLTeS20QZVHSxaMUsFRkYtzL+3MzjEbhap2Rwk8
h0I+kdixQPL/VgDaocmHuYGAMssw2aGBcEwOaZwbAaNZ7jU8Sm3ycm9zSt8WkdQ4
CHM03Ps2eTaNs8xJFhmdUcjOHVmH9OcSSxQmmAs7MVG0zwf59M0ZQBFh7Cg9cL+5
Mb1pNgpoUEWU7GIzGGDvOZ6kI9YseohwNyldoOTrM8RWD6AzKVcJWPPip6uLSRjJ
gWSa0KgAXsxXGRsj2TUIQNw/un4h60Sp1jMUfs2WfwvHoKHAoNxwBC/dT1pt6Eno
Nigl/2JI1kqAftCQAACw1mu2ONpysZoP2Qn/+HkFySRksXSQvEfnRV8s/41etfH9
zZcSX5EfCaIyH/73lc9r8kyE3hf1teMuzS6n8v5tr2d7sbufvCZODp2DE2Y4j6vT
1ouB6QYTPDSUiD4HUgTjbM5DvqoeUUjiNNhYx34xGTFNCy2HkXGfsSOYvwMOQD8C
ig8UXMyqeGWgO+1X7g6aTDWoJX4hqWtO2dPRCYOOBUYqSIX91ZInf3ZlhnEKNP3g
SBY9MqT3wYYhAL2YmSYiuTJ2F0ewmNT3McIMvxSDDRSuAVkBf7SS+uA0D75qVgZY
pOjnhg3DFV09PWldHybgUqhIeOlXxRtpwR47QBLnXBUmOIuBXyf3bgXjdcnNr0d9
5Z/8viejBhanmn/hk0tehj/LTwutEwMAjEIm4y/G6ymMNPXtCZ5ciI0wl5lTCndV
QzZw7Pu7RHma6j+jkq/KBRuJzJYRliTf7C7lRZDYi5a0RPK5Rhv27YahJU06txPH
H04wTS4BabLoCAEfmLekHnZJYuWAZKkOXz0JeZpp0O3BRh3iDP898SdAq0l7V5ta
+DAXHsPREodK4poj1SyT1Sh1zAOdjuIM4Xeu9o/fR6uEHkleynUYB/9XuH4O9Qlu
EUPDcNS8NzxwmdSL2lCpJYYfM80154XSQVvS59EMM5zEfS3CwC6+4jgZd1uB6M0D
CcsscEM/bjxNWN+kIBAnX9YwNmACrEHZzG3LOX+UsQH08eGWMYx2XgtGnL/NreTW
x10KUGa5xuulSQArjTC86kgHMXi91xRZOdG/NW7uji3l0x60RsIpOVBCTfMOnD+L
AO5Bg1TSQUEQ8YZG0mw403bsN2psjjAipApRuFX/xtVwFQPrCUIt2A1YlPt+2Quk
QtI5M3WJg7eIrOSmiIIHD097Hnu/US8ybPYlEMcIDRv8NxcFPUCFef5CQbcTK66b
zGgqJq7RxJt756IK564kn+te8HfLlsHbNL6N5wNaZiO4DjcTp0BsiNzkOL4xA5Kr
CQ2FL3WBHBOzwfuOjJZ/tgHuU6HYwXYqHMB/TOW+uOqYg6fDVu4V9RYLl+VOzQae
Vcl+zzMC4HEjyDv9kBx24eAkdRlA7l2TYOhgP4eaX4boAA5GhaPu6gskLscybcmJ
zI/NCpxFn7n9xzJ7BWxcjpJtUG12wJeJLljEAJOPtJ2O/5xSl4KNaYc1XXcjtt9X
oeCLpDsW0gDQZFHm/Nd77Cvjy4akoyiJFho1pUH13w4mxvRr7HHZKGRh7pJ3ybGo
TYjztbTfXm5gLYJidplDpQ6mYQ89pjSP1jbCzXEGjzBWhT1fNs6fbUktI52VF3eN
fTaXfNMlu+QnUaWh2nfwgAd2w8S1KO6sfnnwjA0Tidmdd3GeD6wHlbv+PuOMawgI
BzJnc2biI9OzVRvUK38Nko27IwZd7PJLGupsj543oWSt0TAlIWsr6Nv2zn6b3zZV
4QZmzsLnGaA6xTuAsxqsWvjStimODxQFEeBtMQYKWRLdYdTKqXMR/ik24EO9iy9q
U/5tz21Fz+ETR8mRsyrpjvRhmy+/Wq4HtsOArsssaktMNotj8lvL5tuZj9F0UCWz
Tfi08tifIBF35vR/L46uEU/6wQtlIAix7BBrhnNL0AxN7tUkDoHaIQumjAxQ0Vll
jwOafq1KL21ONcMrDrI+ogDWth/YjYj4JdXQUkHX2ud+Yo3VKs6QgIrivHGEJu0t
iWIGiWph++ICA/Ln6fLTP54cXsWU9nDNKOLevb+CcmMHqQ8K/HXWgohwbj7poMNO
P/UzrMubGjwSD0PDUAMlpTvpfCK3M24caMO/F27SXPk4euVSEbrTwdG4k7hxko8B
8TMtFRXIR+GLOCfsmEOgQnjAI0PghguVJ3AyFw+Wzzswwfsyuc27PyM5AI7pOFyl
r5OhTHmzzfy1i1Yx7hZagWKn1kCQwLEJd2pHqB4uZE9gSgkDEwr3R9OORslSWMJa
zwlcY6/jnWMKtK7CrhLkgR1ZGOujIZOJhxs2615CZK2CN6o9frDG7BAMjYvLUd8W
Ctq0tepJuWLZ/KnLkv8+mLq+RxVGPRaU1U+MrWyIkUQ1Q+4lK4c/Zi0bq8AtY853
TMtfQMyqm1aPAQzmF2pZq0cMsc81A8EWMfWGmpvU1r5lbAgq+mJJFePj8T0Wszoq
pMzk7WQ0+VBS4ypZwA1sP/aDlejZuqnjM9w9ijvM3Z3ItDsBrMf93hkq05e9TKAD
yNf3lZgMURgvQQ3qoDO9A1Ifwyq2neeRHpcgq0PKUKac+EmlzxhXikre12S5yr7e
aqGOSd6HxhCXzse2tActkDc9sR7DyCLoWNXHWf8Qc7aD1Cij4U3OyEjGiuV1wx1U
HQj+XWRamLfvQP5hVU9YiFuA7CtbnRbTxCHndm3+a+cAA66QbGjEN6/IPHy7tH83
2cTCRRzijkbOFipIv9oamFimxUHgo2fA4tRKZhw1vd/BhybpIbzsPiE7uo48qr77
0hd+5pFksljLWzt9NWIvtvoeBgHYmYASWsC38Xa0aKG8t2sUBXxRcajGsCTrUnSj
JS6x9Hs64r8Glht4y8GnRdUukXU8ou3v14G3pq/VYKoc0VqHxnntn0sk7Jb4aZKR
PpC41igU30Tw3ECCQlrM7i8jnX12aY5hR+ig4AykMkOM/Mr7k9zAJtJZsJQD9Viv
OvjHsvtQPI0FizJVok4b/l/qdacJQkEJl0RKPXSUmZer4ebYa1xWDeh4FvUN1hK4
IaKu6Blr2C0Pd48Lq+Uv6I1AwNiQKid509zieU3jF+UL1PhyNqtk7Tbp9Ike5FFa
ypJMdKIAJGuSoNRRaSBvhUliba1bsOW3Tqzbcltg4Xxn5/ja61JQtImtgTmQiqNL
RicDrpKHNRC2kPSYE8fqExHSJabCUlual5GdvCs/6Pf84q0wot4MWFmPNzXVXUjT
v9w52Ljn3rbURLroSIYZ4t7zvYqO9/AuEnNjwl98GDU8ssZsOq5ObVcGI+uNbKkS
uCWQDB1UklP5P8SyGvfQ+tKtBxamyymJR3ZwL+J24WBu2zXftVtivXsphp1pcM/K
9Sja7jvervmAPszyTswYvWBJ/Eh84SsKLx3zl8mADeF6UL46tKBDfJqzmnmji6zE
RREItu/i0TgVVJT362bh/QmOdu4/YaGRgZGOu5nTQd8KOjVcM5gBd5o/FV396u9y
1hV3tNlWlKQ+fhP1tsqGcjxvC1CmwY/UaaV81iaqFn5+DIx0wQie9YxfHCxo3ifu
oOud4LsLHrZeNOF9NnfLM1vp0vk1klnM1bDpLXm0Zp7sTRQUTB/vLC45I5SuNiTE
`pragma protect end_protected
