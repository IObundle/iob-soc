// S5_PFL.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module S5_PFL (
		input  wire [1:0]  button_external_connection_export,               //      button_external_connection.export
		output wire [27:0] cfi_flash_atb_bridge_0_out_tcm_address_out,      //      cfi_flash_atb_bridge_0_out.tcm_address_out
		output wire [0:0]  cfi_flash_atb_bridge_0_out_tcm_read_n_out,       //                                .tcm_read_n_out
		output wire [0:0]  cfi_flash_atb_bridge_0_out_tcm_write_n_out,      //                                .tcm_write_n_out
		inout  wire [31:0] cfi_flash_atb_bridge_0_out_tcm_data_out,         //                                .tcm_data_out
		output wire [0:0]  cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out, //                                .tcm_chipselect_n_out
		output wire [7:0]  hex0_external_connection_export,                 //        hex0_external_connection.export
		output wire [7:0]  hex1_external_connection_export,                 //        hex1_external_connection.export
		output wire [3:0]  led_bracket_external_connection_export,          // led_bracket_external_connection.export
		output wire [3:0]  led_external_connection_export,                  //         led_external_connection.export
		output wire [1:0]  led_rj45_external_connection_export,             //    led_rj45_external_connection.export
		input  wire        merged_resets_in_reset_reset_n,                  //          merged_resets_in_reset.reset_n
		input  wire        sys_clk_clk,                                     //                         sys_clk.clk
		output wire        temp_scl_external_connection_export,             //    temp_scl_external_connection.export
		inout  wire        temp_sda_external_connection_export              //    temp_sda_external_connection.export
	);

	wire         ext_flash_tcm_data_outen;                                  // ext_flash:tcm_data_outen -> cfi_flash_atb_bridge_0:tcs_tcm_data_outen
	wire         ext_flash_tcm_request;                                     // ext_flash:tcm_request -> cfi_flash_atb_bridge_0:request
	wire         ext_flash_tcm_write_n_out;                                 // ext_flash:tcm_write_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_write_n_out
	wire         ext_flash_tcm_read_n_out;                                  // ext_flash:tcm_read_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_read_n_out
	wire         ext_flash_tcm_grant;                                       // cfi_flash_atb_bridge_0:grant -> ext_flash:tcm_grant
	wire         ext_flash_tcm_chipselect_n_out;                            // ext_flash:tcm_chipselect_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_chipselect_n_out
	wire  [27:0] ext_flash_tcm_address_out;                                 // ext_flash:tcm_address_out -> cfi_flash_atb_bridge_0:tcs_tcm_address_out
	wire  [31:0] ext_flash_tcm_data_out;                                    // ext_flash:tcm_data_out -> cfi_flash_atb_bridge_0:tcs_tcm_data_out
	wire  [31:0] ext_flash_tcm_data_in;                                     // cfi_flash_atb_bridge_0:tcs_tcm_data_in -> ext_flash:tcm_data_in
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [28:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [28:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pb_cpu_to_io_s0_readdata;                // pb_cpu_to_io:s0_readdata -> mm_interconnect_0:pb_cpu_to_io_s0_readdata
	wire         mm_interconnect_0_pb_cpu_to_io_s0_waitrequest;             // pb_cpu_to_io:s0_waitrequest -> mm_interconnect_0:pb_cpu_to_io_s0_waitrequest
	wire         mm_interconnect_0_pb_cpu_to_io_s0_debugaccess;             // mm_interconnect_0:pb_cpu_to_io_s0_debugaccess -> pb_cpu_to_io:s0_debugaccess
	wire  [10:0] mm_interconnect_0_pb_cpu_to_io_s0_address;                 // mm_interconnect_0:pb_cpu_to_io_s0_address -> pb_cpu_to_io:s0_address
	wire         mm_interconnect_0_pb_cpu_to_io_s0_read;                    // mm_interconnect_0:pb_cpu_to_io_s0_read -> pb_cpu_to_io:s0_read
	wire   [3:0] mm_interconnect_0_pb_cpu_to_io_s0_byteenable;              // mm_interconnect_0:pb_cpu_to_io_s0_byteenable -> pb_cpu_to_io:s0_byteenable
	wire         mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid;           // pb_cpu_to_io:s0_readdatavalid -> mm_interconnect_0:pb_cpu_to_io_s0_readdatavalid
	wire         mm_interconnect_0_pb_cpu_to_io_s0_write;                   // mm_interconnect_0:pb_cpu_to_io_s0_write -> pb_cpu_to_io:s0_write
	wire  [31:0] mm_interconnect_0_pb_cpu_to_io_s0_writedata;               // mm_interconnect_0:pb_cpu_to_io_s0_writedata -> pb_cpu_to_io:s0_writedata
	wire   [0:0] mm_interconnect_0_pb_cpu_to_io_s0_burstcount;              // mm_interconnect_0:pb_cpu_to_io_s0_burstcount -> pb_cpu_to_io:s0_burstcount
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;             // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;               // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [18:0] mm_interconnect_0_onchip_memory_s1_address;                // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;             // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                  // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;              // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                  // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire  [31:0] mm_interconnect_0_ext_flash_uas_readdata;                  // ext_flash:uas_readdata -> mm_interconnect_0:ext_flash_uas_readdata
	wire         mm_interconnect_0_ext_flash_uas_waitrequest;               // ext_flash:uas_waitrequest -> mm_interconnect_0:ext_flash_uas_waitrequest
	wire         mm_interconnect_0_ext_flash_uas_debugaccess;               // mm_interconnect_0:ext_flash_uas_debugaccess -> ext_flash:uas_debugaccess
	wire  [27:0] mm_interconnect_0_ext_flash_uas_address;                   // mm_interconnect_0:ext_flash_uas_address -> ext_flash:uas_address
	wire         mm_interconnect_0_ext_flash_uas_read;                      // mm_interconnect_0:ext_flash_uas_read -> ext_flash:uas_read
	wire   [3:0] mm_interconnect_0_ext_flash_uas_byteenable;                // mm_interconnect_0:ext_flash_uas_byteenable -> ext_flash:uas_byteenable
	wire         mm_interconnect_0_ext_flash_uas_readdatavalid;             // ext_flash:uas_readdatavalid -> mm_interconnect_0:ext_flash_uas_readdatavalid
	wire         mm_interconnect_0_ext_flash_uas_lock;                      // mm_interconnect_0:ext_flash_uas_lock -> ext_flash:uas_lock
	wire         mm_interconnect_0_ext_flash_uas_write;                     // mm_interconnect_0:ext_flash_uas_write -> ext_flash:uas_write
	wire  [31:0] mm_interconnect_0_ext_flash_uas_writedata;                 // mm_interconnect_0:ext_flash_uas_writedata -> ext_flash:uas_writedata
	wire   [2:0] mm_interconnect_0_ext_flash_uas_burstcount;                // mm_interconnect_0:ext_flash_uas_burstcount -> ext_flash:uas_burstcount
	wire         pb_cpu_to_io_m0_waitrequest;                               // mm_interconnect_1:pb_cpu_to_io_m0_waitrequest -> pb_cpu_to_io:m0_waitrequest
	wire  [31:0] pb_cpu_to_io_m0_readdata;                                  // mm_interconnect_1:pb_cpu_to_io_m0_readdata -> pb_cpu_to_io:m0_readdata
	wire         pb_cpu_to_io_m0_debugaccess;                               // pb_cpu_to_io:m0_debugaccess -> mm_interconnect_1:pb_cpu_to_io_m0_debugaccess
	wire  [10:0] pb_cpu_to_io_m0_address;                                   // pb_cpu_to_io:m0_address -> mm_interconnect_1:pb_cpu_to_io_m0_address
	wire         pb_cpu_to_io_m0_read;                                      // pb_cpu_to_io:m0_read -> mm_interconnect_1:pb_cpu_to_io_m0_read
	wire   [3:0] pb_cpu_to_io_m0_byteenable;                                // pb_cpu_to_io:m0_byteenable -> mm_interconnect_1:pb_cpu_to_io_m0_byteenable
	wire         pb_cpu_to_io_m0_readdatavalid;                             // mm_interconnect_1:pb_cpu_to_io_m0_readdatavalid -> pb_cpu_to_io:m0_readdatavalid
	wire  [31:0] pb_cpu_to_io_m0_writedata;                                 // pb_cpu_to_io:m0_writedata -> mm_interconnect_1:pb_cpu_to_io_m0_writedata
	wire         pb_cpu_to_io_m0_write;                                     // pb_cpu_to_io:m0_write -> mm_interconnect_1:pb_cpu_to_io_m0_write
	wire   [0:0] pb_cpu_to_io_m0_burstcount;                                // pb_cpu_to_io:m0_burstcount -> mm_interconnect_1:pb_cpu_to_io_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;             // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_timer_s1_chipselect;                     // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                        // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_write;                          // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                      // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire  [31:0] mm_interconnect_1_button_s1_readdata;                      // button:readdata -> mm_interconnect_1:button_s1_readdata
	wire   [1:0] mm_interconnect_1_button_s1_address;                       // mm_interconnect_1:button_s1_address -> button:address
	wire         mm_interconnect_1_led_s1_chipselect;                       // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                         // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                          // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_write;                            // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                        // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire         mm_interconnect_1_temp_sda_s1_chipselect;                  // mm_interconnect_1:temp_sda_s1_chipselect -> temp_sda:chipselect
	wire  [31:0] mm_interconnect_1_temp_sda_s1_readdata;                    // temp_sda:readdata -> mm_interconnect_1:temp_sda_s1_readdata
	wire   [1:0] mm_interconnect_1_temp_sda_s1_address;                     // mm_interconnect_1:temp_sda_s1_address -> temp_sda:address
	wire         mm_interconnect_1_temp_sda_s1_write;                       // mm_interconnect_1:temp_sda_s1_write -> temp_sda:write_n
	wire  [31:0] mm_interconnect_1_temp_sda_s1_writedata;                   // mm_interconnect_1:temp_sda_s1_writedata -> temp_sda:writedata
	wire         mm_interconnect_1_temp_scl_s1_chipselect;                  // mm_interconnect_1:temp_scl_s1_chipselect -> temp_scl:chipselect
	wire  [31:0] mm_interconnect_1_temp_scl_s1_readdata;                    // temp_scl:readdata -> mm_interconnect_1:temp_scl_s1_readdata
	wire   [1:0] mm_interconnect_1_temp_scl_s1_address;                     // mm_interconnect_1:temp_scl_s1_address -> temp_scl:address
	wire         mm_interconnect_1_temp_scl_s1_write;                       // mm_interconnect_1:temp_scl_s1_write -> temp_scl:write_n
	wire  [31:0] mm_interconnect_1_temp_scl_s1_writedata;                   // mm_interconnect_1:temp_scl_s1_writedata -> temp_scl:writedata
	wire         mm_interconnect_1_hex0_s1_chipselect;                      // mm_interconnect_1:hex0_s1_chipselect -> hex0:chipselect
	wire  [31:0] mm_interconnect_1_hex0_s1_readdata;                        // hex0:readdata -> mm_interconnect_1:hex0_s1_readdata
	wire   [1:0] mm_interconnect_1_hex0_s1_address;                         // mm_interconnect_1:hex0_s1_address -> hex0:address
	wire         mm_interconnect_1_hex0_s1_write;                           // mm_interconnect_1:hex0_s1_write -> hex0:write_n
	wire  [31:0] mm_interconnect_1_hex0_s1_writedata;                       // mm_interconnect_1:hex0_s1_writedata -> hex0:writedata
	wire         mm_interconnect_1_hex1_s1_chipselect;                      // mm_interconnect_1:hex1_s1_chipselect -> hex1:chipselect
	wire  [31:0] mm_interconnect_1_hex1_s1_readdata;                        // hex1:readdata -> mm_interconnect_1:hex1_s1_readdata
	wire   [1:0] mm_interconnect_1_hex1_s1_address;                         // mm_interconnect_1:hex1_s1_address -> hex1:address
	wire         mm_interconnect_1_hex1_s1_write;                           // mm_interconnect_1:hex1_s1_write -> hex1:write_n
	wire  [31:0] mm_interconnect_1_hex1_s1_writedata;                       // mm_interconnect_1:hex1_s1_writedata -> hex1:writedata
	wire         mm_interconnect_1_led_rj45_s1_chipselect;                  // mm_interconnect_1:led_rj45_s1_chipselect -> led_rj45:chipselect
	wire  [31:0] mm_interconnect_1_led_rj45_s1_readdata;                    // led_rj45:readdata -> mm_interconnect_1:led_rj45_s1_readdata
	wire   [1:0] mm_interconnect_1_led_rj45_s1_address;                     // mm_interconnect_1:led_rj45_s1_address -> led_rj45:address
	wire         mm_interconnect_1_led_rj45_s1_write;                       // mm_interconnect_1:led_rj45_s1_write -> led_rj45:write_n
	wire  [31:0] mm_interconnect_1_led_rj45_s1_writedata;                   // mm_interconnect_1:led_rj45_s1_writedata -> led_rj45:writedata
	wire         mm_interconnect_1_led_bracket_s1_chipselect;               // mm_interconnect_1:led_bracket_s1_chipselect -> led_bracket:chipselect
	wire  [31:0] mm_interconnect_1_led_bracket_s1_readdata;                 // led_bracket:readdata -> mm_interconnect_1:led_bracket_s1_readdata
	wire   [1:0] mm_interconnect_1_led_bracket_s1_address;                  // mm_interconnect_1:led_bracket_s1_address -> led_bracket:address
	wire         mm_interconnect_1_led_bracket_s1_write;                    // mm_interconnect_1:led_bracket_s1_write -> led_bracket:write_n
	wire  [31:0] mm_interconnect_1_led_bracket_s1_writedata;                // mm_interconnect_1:led_bracket_s1_writedata -> led_bracket:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [button:reset_n, cfi_flash_atb_bridge_0:reset, cpu:reset_n, ext_flash:reset_reset, irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pb_cpu_to_io_reset_reset_bridge_in_reset_reset, onchip_memory:reset, pb_cpu_to_io:reset, rst_translator:in_reset, sysid:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in0]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [hex0:reset_n, hex1:reset_n, led_bracket:reset_n, led_rj45:reset_n, mm_interconnect_1:temp_sda_reset_reset_bridge_in_reset_reset, temp_scl:reset_n, temp_sda:reset_n]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [rst_controller:reset_in0, rst_controller_001:reset_in0]

	S5_PFL_button button (
		.clk      (sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_1_button_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_button_s1_readdata), //                    .readdata
		.in_port  (button_external_connection_export)     // external_connection.export
	);

	S5_PFL_cfi_flash_atb_bridge_0 cfi_flash_atb_bridge_0 (
		.clk                      (sys_clk_clk),                                     //   clk.clk
		.reset                    (rst_controller_reset_out_reset),                  // reset.reset
		.request                  (ext_flash_tcm_request),                           //   tcs.request
		.grant                    (ext_flash_tcm_grant),                             //      .grant
		.tcs_tcm_address_out      (ext_flash_tcm_address_out),                       //      .address_out
		.tcs_tcm_read_n_out       (ext_flash_tcm_read_n_out),                        //      .read_n_out
		.tcs_tcm_write_n_out      (ext_flash_tcm_write_n_out),                       //      .write_n_out
		.tcs_tcm_data_out         (ext_flash_tcm_data_out),                          //      .data_out
		.tcs_tcm_data_outen       (ext_flash_tcm_data_outen),                        //      .data_outen
		.tcs_tcm_data_in          (ext_flash_tcm_data_in),                           //      .data_in
		.tcs_tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                  //      .chipselect_n_out
		.tcm_address_out          (cfi_flash_atb_bridge_0_out_tcm_address_out),      //   out.tcm_address_out
		.tcm_read_n_out           (cfi_flash_atb_bridge_0_out_tcm_read_n_out),       //      .tcm_read_n_out
		.tcm_write_n_out          (cfi_flash_atb_bridge_0_out_tcm_write_n_out),      //      .tcm_write_n_out
		.tcm_data_out             (cfi_flash_atb_bridge_0_out_tcm_data_out),         //      .tcm_data_out
		.tcm_chipselect_n_out     (cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out)  //      .tcm_chipselect_n_out
	);

	S5_PFL_cpu cpu (
		.clk                                 (sys_clk_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	S5_PFL_ext_flash #(
		.TCM_ADDRESS_W                  (28),
		.TCM_DATA_W                     (32),
		.TCM_BYTEENABLE_W               (4),
		.TCM_READ_WAIT                  (144),
		.TCM_WRITE_WAIT                 (144),
		.TCM_SETUP_WAIT                 (33),
		.TCM_DATA_HOLD                  (33),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (4),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) ext_flash (
		.clk_clk              (sys_clk_clk),                                   //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                // reset.reset
		.uas_address          (mm_interconnect_0_ext_flash_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_ext_flash_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_ext_flash_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_ext_flash_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_ext_flash_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_ext_flash_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_ext_flash_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_ext_flash_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_ext_flash_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_ext_flash_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_ext_flash_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (ext_flash_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (ext_flash_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (ext_flash_tcm_request),                         //      .request
		.tcm_grant            (ext_flash_tcm_grant),                           //      .grant
		.tcm_address_out      (ext_flash_tcm_address_out),                     //      .address_out
		.tcm_data_out         (ext_flash_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (ext_flash_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (ext_flash_tcm_data_in)                          //      .data_in
	);

	S5_PFL_hex0 hex0 (
		.clk        (sys_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex0_external_connection_export)       // external_connection.export
	);

	S5_PFL_hex0 hex1 (
		.clk        (sys_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_hex1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_hex1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_hex1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_hex1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_hex1_s1_readdata),   //                    .readdata
		.out_port   (hex1_external_connection_export)       // external_connection.export
	);

	S5_PFL_jtag_uart jtag_uart (
		.clk            (sys_clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	S5_PFL_led led (
		.clk        (sys_clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	S5_PFL_led_bracket led_bracket (
		.clk        (sys_clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_led_bracket_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_bracket_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_bracket_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_bracket_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_bracket_s1_readdata),   //                    .readdata
		.out_port   (led_bracket_external_connection_export)       // external_connection.export
	);

	S5_PFL_led_rj45 led_rj45 (
		.clk        (sys_clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_led_rj45_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_rj45_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_rj45_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_rj45_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_rj45_s1_readdata),   //                    .readdata
		.out_port   (led_rj45_external_connection_export)       // external_connection.export
	);

	S5_PFL_onchip_memory onchip_memory (
		.clk        (sys_clk_clk),                                   //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (11),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pb_cpu_to_io (
		.clk              (sys_clk_clk),                                     //   clk.clk
		.reset            (rst_controller_reset_out_reset),                  // reset.reset
		.s0_waitrequest   (mm_interconnect_0_pb_cpu_to_io_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_pb_cpu_to_io_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_pb_cpu_to_io_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_pb_cpu_to_io_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_pb_cpu_to_io_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_pb_cpu_to_io_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_pb_cpu_to_io_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_pb_cpu_to_io_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_pb_cpu_to_io_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pb_cpu_to_io_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pb_cpu_to_io_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pb_cpu_to_io_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pb_cpu_to_io_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pb_cpu_to_io_m0_writedata),                       //      .writedata
		.m0_address       (pb_cpu_to_io_m0_address),                         //      .address
		.m0_write         (pb_cpu_to_io_m0_write),                           //      .write
		.m0_read          (pb_cpu_to_io_m0_read),                            //      .read
		.m0_byteenable    (pb_cpu_to_io_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pb_cpu_to_io_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                // (terminated)
		.m0_response      (2'b00)                                            // (terminated)
	);

	S5_PFL_sysid sysid (
		.clock    (sys_clk_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	S5_PFL_temp_scl temp_scl (
		.clk        (sys_clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_temp_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_temp_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_temp_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_temp_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_temp_scl_s1_readdata),   //                    .readdata
		.out_port   (temp_scl_external_connection_export)       // external_connection.export
	);

	S5_PFL_temp_sda temp_sda (
		.clk        (sys_clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_temp_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_temp_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_temp_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_temp_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_temp_sda_s1_readdata),   //                    .readdata
		.bidir_port (temp_sda_external_connection_export)       // external_connection.export
	);

	S5_PFL_timer timer (
		.clk        (sys_clk_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	S5_PFL_mm_interconnect_0 mm_interconnect_0 (
		.sys_clk_clk_clk                       (sys_clk_clk),                                       //                     sys_clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address               (cpu_data_master_address),                           //                 cpu_data_master.address
		.cpu_data_master_waitrequest           (cpu_data_master_waitrequest),                       //                                .waitrequest
		.cpu_data_master_byteenable            (cpu_data_master_byteenable),                        //                                .byteenable
		.cpu_data_master_read                  (cpu_data_master_read),                              //                                .read
		.cpu_data_master_readdata              (cpu_data_master_readdata),                          //                                .readdata
		.cpu_data_master_readdatavalid         (cpu_data_master_readdatavalid),                     //                                .readdatavalid
		.cpu_data_master_write                 (cpu_data_master_write),                             //                                .write
		.cpu_data_master_writedata             (cpu_data_master_writedata),                         //                                .writedata
		.cpu_data_master_debugaccess           (cpu_data_master_debugaccess),                       //                                .debugaccess
		.cpu_instruction_master_address        (cpu_instruction_master_address),                    //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                //                                .waitrequest
		.cpu_instruction_master_read           (cpu_instruction_master_read),                       //                                .read
		.cpu_instruction_master_readdata       (cpu_instruction_master_readdata),                   //                                .readdata
		.cpu_instruction_master_readdatavalid  (cpu_instruction_master_readdatavalid),              //                                .readdatavalid
		.cpu_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),     //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),       //                                .write
		.cpu_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),        //                                .read
		.cpu_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                                .readdata
		.cpu_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                                .writedata
		.cpu_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                                .byteenable
		.cpu_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                                .debugaccess
		.ext_flash_uas_address                 (mm_interconnect_0_ext_flash_uas_address),           //                   ext_flash_uas.address
		.ext_flash_uas_write                   (mm_interconnect_0_ext_flash_uas_write),             //                                .write
		.ext_flash_uas_read                    (mm_interconnect_0_ext_flash_uas_read),              //                                .read
		.ext_flash_uas_readdata                (mm_interconnect_0_ext_flash_uas_readdata),          //                                .readdata
		.ext_flash_uas_writedata               (mm_interconnect_0_ext_flash_uas_writedata),         //                                .writedata
		.ext_flash_uas_burstcount              (mm_interconnect_0_ext_flash_uas_burstcount),        //                                .burstcount
		.ext_flash_uas_byteenable              (mm_interconnect_0_ext_flash_uas_byteenable),        //                                .byteenable
		.ext_flash_uas_readdatavalid           (mm_interconnect_0_ext_flash_uas_readdatavalid),     //                                .readdatavalid
		.ext_flash_uas_waitrequest             (mm_interconnect_0_ext_flash_uas_waitrequest),       //                                .waitrequest
		.ext_flash_uas_lock                    (mm_interconnect_0_ext_flash_uas_lock),              //                                .lock
		.ext_flash_uas_debugaccess             (mm_interconnect_0_ext_flash_uas_debugaccess),       //                                .debugaccess
		.onchip_memory_s1_address              (mm_interconnect_0_onchip_memory_s1_address),        //                onchip_memory_s1.address
		.onchip_memory_s1_write                (mm_interconnect_0_onchip_memory_s1_write),          //                                .write
		.onchip_memory_s1_readdata             (mm_interconnect_0_onchip_memory_s1_readdata),       //                                .readdata
		.onchip_memory_s1_writedata            (mm_interconnect_0_onchip_memory_s1_writedata),      //                                .writedata
		.onchip_memory_s1_byteenable           (mm_interconnect_0_onchip_memory_s1_byteenable),     //                                .byteenable
		.onchip_memory_s1_chipselect           (mm_interconnect_0_onchip_memory_s1_chipselect),     //                                .chipselect
		.onchip_memory_s1_clken                (mm_interconnect_0_onchip_memory_s1_clken),          //                                .clken
		.pb_cpu_to_io_s0_address               (mm_interconnect_0_pb_cpu_to_io_s0_address),         //                 pb_cpu_to_io_s0.address
		.pb_cpu_to_io_s0_write                 (mm_interconnect_0_pb_cpu_to_io_s0_write),           //                                .write
		.pb_cpu_to_io_s0_read                  (mm_interconnect_0_pb_cpu_to_io_s0_read),            //                                .read
		.pb_cpu_to_io_s0_readdata              (mm_interconnect_0_pb_cpu_to_io_s0_readdata),        //                                .readdata
		.pb_cpu_to_io_s0_writedata             (mm_interconnect_0_pb_cpu_to_io_s0_writedata),       //                                .writedata
		.pb_cpu_to_io_s0_burstcount            (mm_interconnect_0_pb_cpu_to_io_s0_burstcount),      //                                .burstcount
		.pb_cpu_to_io_s0_byteenable            (mm_interconnect_0_pb_cpu_to_io_s0_byteenable),      //                                .byteenable
		.pb_cpu_to_io_s0_readdatavalid         (mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid),   //                                .readdatavalid
		.pb_cpu_to_io_s0_waitrequest           (mm_interconnect_0_pb_cpu_to_io_s0_waitrequest),     //                                .waitrequest
		.pb_cpu_to_io_s0_debugaccess           (mm_interconnect_0_pb_cpu_to_io_s0_debugaccess)      //                                .debugaccess
	);

	S5_PFL_mm_interconnect_1 mm_interconnect_1 (
		.sys_clk_clk_clk                                (sys_clk_clk),                                               //                              sys_clk_clk.clk
		.pb_cpu_to_io_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // pb_cpu_to_io_reset_reset_bridge_in_reset.reset
		.temp_sda_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                        //     temp_sda_reset_reset_bridge_in_reset.reset
		.pb_cpu_to_io_m0_address                        (pb_cpu_to_io_m0_address),                                   //                          pb_cpu_to_io_m0.address
		.pb_cpu_to_io_m0_waitrequest                    (pb_cpu_to_io_m0_waitrequest),                               //                                         .waitrequest
		.pb_cpu_to_io_m0_burstcount                     (pb_cpu_to_io_m0_burstcount),                                //                                         .burstcount
		.pb_cpu_to_io_m0_byteenable                     (pb_cpu_to_io_m0_byteenable),                                //                                         .byteenable
		.pb_cpu_to_io_m0_read                           (pb_cpu_to_io_m0_read),                                      //                                         .read
		.pb_cpu_to_io_m0_readdata                       (pb_cpu_to_io_m0_readdata),                                  //                                         .readdata
		.pb_cpu_to_io_m0_readdatavalid                  (pb_cpu_to_io_m0_readdatavalid),                             //                                         .readdatavalid
		.pb_cpu_to_io_m0_write                          (pb_cpu_to_io_m0_write),                                     //                                         .write
		.pb_cpu_to_io_m0_writedata                      (pb_cpu_to_io_m0_writedata),                                 //                                         .writedata
		.pb_cpu_to_io_m0_debugaccess                    (pb_cpu_to_io_m0_debugaccess),                               //                                         .debugaccess
		.button_s1_address                              (mm_interconnect_1_button_s1_address),                       //                                button_s1.address
		.button_s1_readdata                             (mm_interconnect_1_button_s1_readdata),                      //                                         .readdata
		.hex0_s1_address                                (mm_interconnect_1_hex0_s1_address),                         //                                  hex0_s1.address
		.hex0_s1_write                                  (mm_interconnect_1_hex0_s1_write),                           //                                         .write
		.hex0_s1_readdata                               (mm_interconnect_1_hex0_s1_readdata),                        //                                         .readdata
		.hex0_s1_writedata                              (mm_interconnect_1_hex0_s1_writedata),                       //                                         .writedata
		.hex0_s1_chipselect                             (mm_interconnect_1_hex0_s1_chipselect),                      //                                         .chipselect
		.hex1_s1_address                                (mm_interconnect_1_hex1_s1_address),                         //                                  hex1_s1.address
		.hex1_s1_write                                  (mm_interconnect_1_hex1_s1_write),                           //                                         .write
		.hex1_s1_readdata                               (mm_interconnect_1_hex1_s1_readdata),                        //                                         .readdata
		.hex1_s1_writedata                              (mm_interconnect_1_hex1_s1_writedata),                       //                                         .writedata
		.hex1_s1_chipselect                             (mm_interconnect_1_hex1_s1_chipselect),                      //                                         .chipselect
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.led_s1_address                                 (mm_interconnect_1_led_s1_address),                          //                                   led_s1.address
		.led_s1_write                                   (mm_interconnect_1_led_s1_write),                            //                                         .write
		.led_s1_readdata                                (mm_interconnect_1_led_s1_readdata),                         //                                         .readdata
		.led_s1_writedata                               (mm_interconnect_1_led_s1_writedata),                        //                                         .writedata
		.led_s1_chipselect                              (mm_interconnect_1_led_s1_chipselect),                       //                                         .chipselect
		.led_bracket_s1_address                         (mm_interconnect_1_led_bracket_s1_address),                  //                           led_bracket_s1.address
		.led_bracket_s1_write                           (mm_interconnect_1_led_bracket_s1_write),                    //                                         .write
		.led_bracket_s1_readdata                        (mm_interconnect_1_led_bracket_s1_readdata),                 //                                         .readdata
		.led_bracket_s1_writedata                       (mm_interconnect_1_led_bracket_s1_writedata),                //                                         .writedata
		.led_bracket_s1_chipselect                      (mm_interconnect_1_led_bracket_s1_chipselect),               //                                         .chipselect
		.led_rj45_s1_address                            (mm_interconnect_1_led_rj45_s1_address),                     //                              led_rj45_s1.address
		.led_rj45_s1_write                              (mm_interconnect_1_led_rj45_s1_write),                       //                                         .write
		.led_rj45_s1_readdata                           (mm_interconnect_1_led_rj45_s1_readdata),                    //                                         .readdata
		.led_rj45_s1_writedata                          (mm_interconnect_1_led_rj45_s1_writedata),                   //                                         .writedata
		.led_rj45_s1_chipselect                         (mm_interconnect_1_led_rj45_s1_chipselect),                  //                                         .chipselect
		.sysid_control_slave_address                    (mm_interconnect_1_sysid_control_slave_address),             //                      sysid_control_slave.address
		.sysid_control_slave_readdata                   (mm_interconnect_1_sysid_control_slave_readdata),            //                                         .readdata
		.temp_scl_s1_address                            (mm_interconnect_1_temp_scl_s1_address),                     //                              temp_scl_s1.address
		.temp_scl_s1_write                              (mm_interconnect_1_temp_scl_s1_write),                       //                                         .write
		.temp_scl_s1_readdata                           (mm_interconnect_1_temp_scl_s1_readdata),                    //                                         .readdata
		.temp_scl_s1_writedata                          (mm_interconnect_1_temp_scl_s1_writedata),                   //                                         .writedata
		.temp_scl_s1_chipselect                         (mm_interconnect_1_temp_scl_s1_chipselect),                  //                                         .chipselect
		.temp_sda_s1_address                            (mm_interconnect_1_temp_sda_s1_address),                     //                              temp_sda_s1.address
		.temp_sda_s1_write                              (mm_interconnect_1_temp_sda_s1_write),                       //                                         .write
		.temp_sda_s1_readdata                           (mm_interconnect_1_temp_sda_s1_readdata),                    //                                         .readdata
		.temp_sda_s1_writedata                          (mm_interconnect_1_temp_sda_s1_writedata),                   //                                         .writedata
		.temp_sda_s1_chipselect                         (mm_interconnect_1_temp_sda_s1_chipselect),                  //                                         .chipselect
		.timer_s1_address                               (mm_interconnect_1_timer_s1_address),                        //                                 timer_s1.address
		.timer_s1_write                                 (mm_interconnect_1_timer_s1_write),                          //                                         .write
		.timer_s1_readdata                              (mm_interconnect_1_timer_s1_readdata),                       //                                         .readdata
		.timer_s1_writedata                             (mm_interconnect_1_timer_s1_writedata),                      //                                         .writedata
		.timer_s1_chipselect                            (mm_interconnect_1_timer_s1_chipselect)                      //                                         .chipselect
	);

	S5_PFL_irq_mapper irq_mapper (
		.clk           (sys_clk_clk),                    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (rst_controller_002_reset_out_reset), // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.reset_in2      (~merged_resets_in_reset_reset_n),    // reset_in2.reset
		.clk            (sys_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (rst_controller_002_reset_out_reset), // reset_in0.reset
		.clk            (sys_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (~merged_resets_in_reset_reset_n),    // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
