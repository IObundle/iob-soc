// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Io8EQ01zGC2ZEfKLkPllmuihSRIx18cXoIHmPHOtseHXdovI16MTHwCmEbcQnyUn
TZXUmsY6qrvuYzf3gUXDTHzVPolH2St7wVZb/7OFpRTxffpu+vTeU27JtesqVb1h
H5QWbR+sdnjSLNtA+xGZ0MGP0H4z6jxqvK0kDd9KncU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31456)
M9PW+fFQi4eZGUM/s8BmjttKw+wu8G0MJNLz9UE5E1XCclgh6Cpxnp3vzpKOy1zK
z8iMbsVoSypg2tDKtA4coFbfjEVYn7MTEiULLB7G3gxnnZfN/uDjI6blsaq8w5GJ
6NwCYN3So0sLj74zWmMFE+xq3HkPxMD5Ci7wgQiUd5FwwfGQoKfUDUE637DrxN3F
ya0fidcT7RDwaEgzChMdvmLs4X5TtHL79Q9iWLf+D8XU7rldmJnGq3IiyK+eFzTa
PlT5nMS4sakMCOkWajYATMDPstYjhGW8nMvPY2l0Wf917LwrAfZ7XUbHfJlCvkOJ
Nts/kLca4sGFYXsfiu8vNHgYbiPOsU/dBYhMv0FNX76+8puqruBIyJEslGG2ycqp
IF0ZC5fQdqRHoETA1lJiJ+jwRMZ/nzvUNmKwBsaVSzDUKVnCF0bswGFIpT/fdUtm
sZTSR9iWOillgxa5rf/u9lXiKgmonnRXPjpL9ktmtOvp9XRRTGDk1ntmcqjMj4CJ
Ofkh1L0GBJIVy1q9ms28pKtRpe00Gq59+skXdzf2xpJeZDil7rSsKWGq1SZgSpdJ
p8mYv3m1NVz1k8xsyuB+p1HqF7LSsY6R5kPCCA5ArETZ6K3PbQCniX+2IsFOMQD1
uWNFC3vIjaz6nQGkLfgbMXibsYGB+azmZ6ImAaqPtPGxnCQMsTBuSn9sMoX0mXLc
DgRV8D4VjDpmvyFUvGzQRGG7TJG/8Z7NXnwa+IPPyHPhaOBj6suxSOC7wLralVKN
iB4wkfW/LSJWbGPvrO6RIIWbtW+DzQA8ZK8YmOEASgTP8DtQR1u8FunCvr53WhKE
2/x338hXYQ+/2q4quxTVUz4Wpd3IkL2rfxvfFxr5UaUh15m472bFOeJxfjEZQh3S
hTn1fKhN3UfFPt2d+gTCn/4aXx8ootu99qikMw40F+4Ahj+Q2jiZaC9WxznGb5ZR
BY1Yv3R+UbVB+cNSnn8qGcnGs8SrzavYuySV4tALIRj0OVmYWWBw6KfxITpC1weT
jxgzZB9ejVbb5+fCymjsAr1MqMbIXOnbC7xQe7HM2+fOWZN4TsBZ2kUfR3sAWSeb
FDwR3rEevShDL2pR+CirNBfXtruKJkYssPlscm315iM6FGTaEKsVwdOa7K7WKgRo
EoVpfRbpgHCtqMev3F8EUk92s/Jfzdk7vVA9YBF9kSgSO+BQbwI14iyDkJXUq8hw
vFypkP9clAR7NAawZBipSiiuMP2CWfygt4BEjFBUz6JTmVjFv6uLVgwXS3nS3UfQ
gqNErvMZcXeUyQuj4CFJfXmJU1igVkL5lMTBipFT9RRGnwXaO70aySSlr2OItbVU
ffBEhAKhh6ovjZD4KQNIAYyOV48MLEkr/drSAyi3TS8/SmlIDyRX/P3j1rKHfhk0
hluQsou4ts1RWPhZjHb1YVqVSqLHPfRxFDmjSNMMwLDbTEDIMpdu4A27sRHU5fqv
QqNYrxCAqCHg8hsmw3fqtPW29MlBNv7+IOL1EShRTYGXVBKA/8dZxFWs62vS1Z8O
s3tEPob8GIWjCjfHji4TVjBHs1nbFhR8NqJsHM/fJl2lYz3SpdenZHPEw+BIXJmK
ppydCcQyao28ljR3PUUlQfhNS7kLiPtoaFWM6yXunFxXoGDnXXFD5GXMUqecF9jH
SqQLrHEp7b74QzcfHo8XsEWY2clPc8+J/53dJLmHZsNQQ11way61x85jNjO8IvXf
Np6EAST+/VJh7vzRcSRyE9CLfytPnz9oyv57mBKQUs1yiHqM/+TN2ADIQEQsmbJd
N5oNyjS6XZZVd+X8p4OU0u/aj2WAj6Cp1/LlFXpegmEljiaprzr1t5WLqYzhVa8q
CtUOcSMyQj94SKmt3gdsdn86R7ojNGdZovL9AwmLPzPj81SVoo4m2xgSzqAcfTiX
EBbwh64XOlQ1YbXykB9Ki9v5ddMoGbr5XAbLq5xfibYMjCS8efy8TkYHmlmeeMcZ
OT4vuqLcJ8iU79eqccsoFqOnAyBwCL/P39DIz3h8YATsre8ALI49blHLOv5wBrKi
k0nsPxDF//bWnqw/JeEIQtldqgVemuSxp/tjA9NIIuXRjtUV4oRAYBWUrMno+e/C
70fkfXPNLI3CO5r7B9CeInWsPOfUjK5+6HiQX/lBRnV03TCTy9TJZr1jvwFlXhy+
M4D/dYqU90qVY5VcvjtGsI1T+cOk2Chz9j2emNrJlBhw6ZQP/lVciFrj8Jk2ZN8/
11WYvs1VZm6t4jSkcqYVYd00IKXwj31eTRUXfAxfWcMy+pN/e6vhf2gZGDQeE95e
Xm+U6CBQX7m9sjUJzWAIJr8+2EZvvK8gXoJDgNmImgqyA/c4AFQVuta3/Ipf8FlJ
BYFSSrhS5PYVRZKNG+0laBqdOGefzhsmyPF6DxCOemxxqicCXhQcPGMqaaYFRm6/
J5pUHOWM7EfRdyYpO9ZP2aHkVO5KYsg0BYfynMJds7IVIOE1/1B/dSO2sHH+zNjt
oOyafmkOAkbZf09ffv1hy1JL+j7PaIkV9NSNduDvsTtQo+UnW53qspTD9wrWpePF
GW8P9RbaD3d2A4dreHYxoERUsZ2GyJzz8YJEIjpXjtaSgRC2bnKVnQl9kSiIVch9
v9Q/vcMprjc/He6RU/nO4mpRuJf/0A8swy+PUIeiSqme5M1yPv+b1R4M8qmKvm9T
rvE/fYzg0u5wfFvkyTk5okkZK+5OseG0M4uT8NhQHlBr4Ot2x5pxI5YHguBpOKwv
Wi56rCvTcaN6LgvZbithsT7OC5jOdRFyUPnbnz/j9czrN+VMs9omAyY9W88gpPTK
uUyEWHssmogIw0G3j3guD2oE65Y0S3LL1mEPvfzxHDLfjr4PbRB0t1q7CQgiwgLt
t5h1U9BpmcjFn4GkS25TBZyFIxS7evPvgI9TNilBjqNuYZui4UCsDrUI2hHj5Ow0
NGc0gTIxGtKU5TSwAfFyp7Tb6lMOKTYxG6kCK5eddaJYYaqwT/SVbzIs1yhvNNEk
4e5oLBGlyRhCavOZ+MONUbg/Ih5Debrdb6cOZmhTPRrFxkqTLMqFfLV9q4/huAJK
kAx+KBvBPwsogQ7vF7btnNfLBsu1Rx1ffPcOhLsDObN/jDaULR9tqs4/46Mp1BVi
A7xt2Q5JVTOanfbLO0RFnLKomXDGGDNPfPo5jckgG60NsPkBiGq0Ia9Rk6/QOuqU
9AXlEdVe5TfXtvMH/yqxARX3TVdg/k9cgibbLasq9RLYxifgIruW5WC1CwNgqyxh
GNjbHa/N15H/j8lDPHGr38XpHTRagjRTgnNsPmuBAKPNWoULdhpXf15WYTonLSfA
yI5uQPJTrRzosf0+fVrhL7/gYzTt1o7HVPI4BWSothhv3YdCdh/0YmZAjDlcFeYO
a90tZNkt/A70VX5+QVtS1I05CrpPr/+GsTU6p+g76RJwNJ09cfN1f2meGcIvKf+a
k6OzUmeV1p3BMQbqRQdkAHGNokkTuyvpBU/9WPZFeqjgz7LoO0yVJ0yiegqHDF3+
VBbZYPJjkR0SiVrpehH7wiowq5J/EDRD7l9MoETW30TtvF5paleAJIkMQmztoYHu
WfUldVVeYc7b829Hugzgw+I0R5nlMyOkk/SOqqM2d40vlCl8bfoAmfUi3QQ8ivqO
si1pORFGRwLCr53fBsyygmd2h5NfLKFjIZXKUbBa+FnkxqZ0hMNQ2PTWVZV0+3te
vupSu6QZ8kLEWYcUo79paBuGteOVy/KEDZOYW88DAP8D2hWW5zE719iVfLCvz9nj
uBQcwYgPC/4KMv5OWOvSv8lsDACY/8nXuMx+XFWBenio9dyZ2TBQNf1G86SOnqAb
YnUai25uDdX48EoEHy+VzPJey2BoKE1NZ+gS0C7XLT6UN90MoCDd+4Zp0Z/29LUu
BDJtyJ/8MKzSZCw70fF2zDfusA0fO588vyhpc1DOdAQajGiIfGmnz/hJTEghw8dL
L5Le0aOvqYdNfxtgxUuiF+xpmn20e1eGn6RheHUBO2STwAOAD6JoMFH8WS/IazqQ
seVNNBtPHpvi7VS3MLjV/WT4PVjJXWjxt1VNHtDXKB07mjPUyltLj+DdsU6/Ww2k
qk8mzaW7wQaGiG34/nPFue10YsTinL6GLUR1ZfeCrrqKSCeUJC1W3xmwbIy4VpRB
ys7+eNTaIDsJDiQ45lqQ0SOftJ+k0ce0JOSfn57cNDlgjuyUs+hSAaYFGbcjyprj
Ft4NVu+stGwnzOTWt8mNVwcP9N/d3FlRjL6L5DMxyr8VetWgTwy7PlQlV8hquxZJ
fXlt306pGmV64mWWu7pHEF1dzaWcHeu0tyB6v9EzfcHELuwlm/8ofotoTRb2tcLt
QNKvw4b4yVPrB3Ql5rge8wR8KLwrml+G/PtpJjpmdR0w2C11Wo8/5cg4cLRgCwho
9HZKiKHpPXxLYatu6pDStmKW5Mc+vVTYwV6lAEb55nxO1JIkIV4fG/Tv425tozgO
8QDZGA+K7vS21I9cMVoODfIus5G4k+SJ7Ztneq66L+dTPl5CAVPewyFql0YReIvv
NeIBuWsqvX88ANT3jCx3W7lLqGPivdht8N/ABJ7pBInt+oT1rtXZC81bPw6Djg10
FHkFXJfBNoRPSwjDnGcOQxomrOjHxsFBsSA4NqcIlIgMoGRKtJscbUMoDwqH5AKQ
lotlsdE/opndZAjWAoQINU53oFWshFlimIIG36VdDiIeYdBNSnObVzJNi8zOWsbB
TasFwITEl8MZC8x0Ij4bmuFdAm//A30fL2g7TBtg98lleYng8SXj4mNPcz+5Pddc
uE3v+HsvQX2faa2RWkm0kq+c22slOkLK9H3wjEcdFw4yQI81Ao5/uB9WYplMzhE/
QxZttHj11OlKZFtHBtEMBjSM88B35zEQnXkha9ljP3RgAdVXiZQDvJvEIVuRIb50
ZCWRpvAZnJxYTD++XsxHkUtGFCHkK1qBTPh6GY/4xR2wyNGR91IvOk8vlBAvkWQn
A0gakMlpp9OGIKMSLqNHldtn+cLIbu+TGfcQFof1jamVviV5J9m4fukAxe4U+fxM
AwP8Pkw5cklMowlMKih8nIwsM9HsuVnfuqEXf8mB9mB8U3QBEayUwYMXrKyody8M
Y2BI1Z9b56NMb7I1VwXSBOU0FagRXQu5+N42OCyPYW2EW+4bY9o7fiDWsHvOuf7D
4qg/HV6VlEOLxBSnRDKIDgXwsEKOocdlehlBjLZ6NULF/WMhEhSrThWhvgpigXcI
9FwZu/kQ9UqAxSD7TRa2sPFKLpSxGsLwGfm3e+MYkTHxeeeEjGCcUNR1nwiiJlqc
oFoIAeGCmWTsbD9LC0d3hlfgNucyCDyzblv2zGR/ICPACJKH1FPyW8+sLhPyZIMt
DcqqtefuZ2c8ZjEx9e7q1C32YgaGBU/Aye12XN1HoWcPdO8qmK1PD+0psh7WnfGF
ovR+BZRujtjbuU4YV6aQsyPLtO4it4PY3ARazxGMOOXinbfZ0qVM96KIcW2naZuh
FWREDvQmxlMH5Z6eZLeiLH00xr6oOdyzzgwyU4ODar2FRlWnMl7gpPimz+9pFxLQ
IbQJ7n6qcgs9rCKkEQ9DcdLUtnPkMSQI45kDAIUx8tk4WTM30rprxe6oDrqqxkGA
AJ4OsBwAjtCoeIPZJN/XpIarmJJ2YP8EasZLipfbS8/hdM5m6nTuVlCv8rJglf6y
r3RtlmaNidvMI4vZ5E+J1WP51NJJUJ2VLsbExFcIBDmOt0khtAabv/zccRhjWo8p
bThJYr46yHH7c1cHY6TiiyIxGN99liZDnzJOuPm5PGi43hH/RMEJF4NzPU4wyRQb
+tlWBpX05k03EEhBN9urCxRozh7JfuXb3URS/apMmsnMe3v++UOn5gTUVWWZ+vrj
4hJH57Kma7b9GV92Nob9XxX8Y9/y/AAglNZ2URHl//+EMqQi5RefdWZQ1UYR+3Cq
jGiHRaoYHaDvDlOETOj1DVwVhbKZqT5195U+17LqzezAhMwWcUmpQ6FxIhnqZbTF
YnZ8IWZP/fDhMe3wDTDZ6sEsnctON7/Kw+yhPpoKCYwrClfc8KsHeLgl1JlOJPky
B3uSy0EICyItoSGw65uxmaRX7yQ6+4muz1qOrF7DqmCSPRju69Y/R/9Gmh2aQ0j/
T0JDA5n6I7TwOrhav/3A1oTkrmAaMaObLmD8r8wvGze6gMFNYx3LnLzczTzkV2Hc
sh/GiIEJnNLB7DdNQVjcllh/98qpW3XexZB6916Xi8RyINSJJ5b7uwBkh4vSRhZK
frpuj8vxBpf4Nz9hB/vM6E472+c0QyEXkm93dm9WEJwtSzWnFJh3uU73xUVa7JMD
DI3EUxztGyUR+gsGyaxXFIN7dWm709xDws8FqoVgnQT1kyURRJyxEGH+3454CkAQ
/z6XHCXoJkY1xnbvpwLZXAGS3nUR6LI8URFOl45KJaWtjHc0Tsm/USdFUpn0FeIb
SjIAh6b5b5H6byqVCTQqdrVk9Povv+va6zJJG7f+EUhJ+kP6eV8YnQPr1hiNV18C
I5UyoL/PjCtq79ieNuatTFrZNVlHmhOJOxdzy0wQ7DjQlYe5GaIzVQ0YxHwU2vaB
FIiZXsbi6qlo2hMOkM65P5V74u35E2fSoeTKBMUgIDzW6VGAFjozg4kJ9Qd2SYih
Nrj1lbrJO1Mm79LLFNMOjrXnO4sBmwk65YXOv7BmI4tTlfh6VzEPuqCu0HDzR21b
hj6dLqHSnP9UcgdIHhL4UG/Yl47ZbGsrTGWmqiMZOtbPrz3VEXyNreWnvYINjnW/
FepWMg18pko+ddto+uL1AtEEAj/5iyWERqT7DII5zPPJdx9J/qHTitHxnElNcSsY
qyZPw//kNGW14xfjMZnZaMJ2csjBHaZJ17zc+K3JsA6zv+axJEmz0tjpbsRTKYNR
iv0OQWOzAqR4xjiq2zyfGgAzJofl/bh9atu2vPh3O8WoDKI4Z6bhZWdLu2ApVf4F
dazFbRxdsi7OkLqQ00iWHPSIrZXswF6VhgZcj51cRLvSF725yhjdSmZqxY3rlWBM
fVqwYe029mhptgdMTaHgpIjXd+6T5BJTeEvWocQpXL73WYhr+OnBup7gl0SqLPHn
pqxpy+/oM8JODCYEF7sDgwtJHHbI5kS/YL/E/utJnZGKA92WaIq8fA2zkMbTVLPj
JF1jka+rF9i+eH60fp7ecmpgnAk6ZgvKnitpCqotbomnjqEU6uYUtgLeELj2vDYv
0tqsKSrmxOAOcKtezZF0Ih5KxGjn+XIs2bAzI5onvhC5qXcTLCs3aZD189oss6dX
szvuPIXG/vESTw2TePiOwUZ81nHaOuXm8fMsw26gkuDWyJMYnjioy7GI6HSIRPHq
NGelLOvOKOQndZJ9wEq/nlJ3R+Rc64nq7I2rddFCBbaj2E/iZfYgeBcWijfSpVe7
a9atS9QoQzolVVt6NMQ4gdE5zPlqNoGdNHERYypecLiLjquhuNupw9o21+EIjIc1
X6DnwDpgtts6cogr9Telq96/kK879tBFq9BMpHZ+B/s+vzeARRThkG/dOfVKN7Rm
5Izt/DFyXin9L85g15SEgiZAvJfUUlK8F6s2mxQ79QVm5dlYycps9AacbhyQTB1y
REF0uA5+fgRzUX149XBc9HAGy5SLkoBlpMASrP0yUxeBrbOzzeuMTFAWFplMsA5V
TwfJYDmSxTXEBQY704+hfM1nLftja+924sR9QYtqQtrcLx3Tx9xmB9p0tU9MPQWc
QKioDwXszeXDB26zVkqpgKyEPv6LZNbyJFgadraWjsAiPcc/AC9V2KbJdmmgz6S3
dkGB/CEWvrEbpTje27WV7KkhAb1Rda9uta8nomUJBD4fbOsBy+MHxiI/F5C8LOFy
fl95FhkkfRdJvg4Ec4+K3L7zhvrdBcKX1AB/ix1BsIjD09BZffbjoJb3kHjf6dgy
F4mfHU2b+L5LLbtO3mW7xB+fgTv3Wm6aPldPSuLritr/VJQP+OaDDYcfmnSVz3fq
ZWhyRx87Wv/Q+AKzFj4+wEKSDKa8lAqRMHwvfuwLHtWWEcaI+nEG3BloEJDvJaEf
t12DI0HoZR7AUV51T/ExLFFleaverqjJvhIRmxpBJAmVQ3G263WsA87MI7w9s1YW
Bf6hn1QuB6CcXzHwyOVLaQxkrPT7rmVBfQyDK0pB8Thshmsr2z+B66ozI5sH1BEX
UU+0DYI1zdSmfz4xkTTXRWgS2gBiTZn2dUxFTGIGdx6CahDiAKdzZF97MjX8D7q7
aACC3IpEP2Zfrg2NFeA9nL8dgsWZWgkT/8FlVtNNHn3BJI7N/aonqMG1ajD3elUr
DOAiBJwYr2rvHTo00/vVtMa7HsVD1eQOxnpl13qFHF3Hw2aOHtkjiub1UZ52brlv
ygYszWOt/78wVzXAkO9DAQq0wRkIPIrhUX9zCRc+TWDCy/ohdhsV7lIxYcyagb8K
ARjOWSCogK5kLDH6VI2YWg3+XqGAaNNcT5yN4vIQLofo8GVAp36Wk06JA+q/jNQC
0Y4qiDsoT6ZHRVaaco7uGhQqA1y3TS6HXntWHZ1lYawaFnm6VlGmE5xt9Ka9qioI
hvJ1kvjItn/uRmFkgw519b+SDPGK3DwxFag6L9IwG/HWIuLZQyXRxiYGrRmQCtTO
z19qiugUb2kyf67N1m470EQGRjIfpZCI+lwjC8dPRwq70UgXhL/qZVNY0rgZYcWk
CjRoN8Jfc2wbMQVQOwxlLe0orfwxB5g6qF7b18sH28SwevNOc5vnAznyChsEwtrB
+OSGG+7v7xUA/0X25lxXF0HkMw5ie0TG33jzZ0JMCpNP79U3DSs6iJBXIouSE1lA
T3CHTx2wxQgGYftJ5S0yn7FWt2IDPL2jhe9YhN7btNva2OnPQoqZEF0V3dn7Mag2
QINlkMkPLaHdvQdMJ0nK53B1bfPVixPNEtWuTjavtb89PO/U7nPmxIpZ7L9vZ69F
cPRsCw9GFuXgBz68KX90pVELeDqpa+jD143AXc14QwzmMKG7NX58/9Ykqi3mrFLt
7qWRX6oz9gL+gU8XaQ38Am5sVF6ENATmSZrbSw9dg8caWzEa6XqWpv0pnjW74ttF
tHmnZWeqBpz6Vy7dEtICH16AZaS2oNlLiS0mMWFcoVbIrzO2uLGG9CQgk0kM0uZY
/zXJ7OM/cvzLkZr/nBM4uwOlHkgzGstBz20L4aMb0cVvRvAr93BIvi3bq6jryZ34
RPPo0mD8w581sgPqPVmuDQIE4pmaHH97FdMMUGOr9B+ANh6IrW4kPv7sv2zWBfHC
i/x7e4uokzLyh8XOyANQLMHcQnNuyfpbWJ0aeqJTjgQTMEbnVRBabHPHoGQd8glt
En4M/jiwaOwam0ONOhRAw4ekuRe1bjO9P0KOxWHF9VWyEZB8ecpkOIM0vw4MTyAn
JrX2N/+5Ih8zeT1bMStj5WJtrDIqAGxrJLv7HWjmaJwLBvxsXQaJ7PTkXAOjM7QN
D9gIpO961lH0EYsngE1jWEBDtVtItvm5dckeyjCuumfxGXmFkPB7ZSrgaHL/V6x1
iOaVLwkKtY8NyErIBhR6i/2vgrnmeYl1f5NOzAZklkyTSb1fOVTjEFnw0mCU9fXO
+rDF+aBacgVffholEU6j/2Yd4az74wwnzXAMTiscGjR66xfWGdSpefzuuzSmzpxP
KCku2JKql9zUxN2HJdak+Z541ETxJrz8O7gmgoqzeq5h5Ioq46I3tnV9VESm9Egl
0MD6iQ+v6tmP+6vHuB+VOVEFdnX2JcKci/AZgLheAl679m70k47Jn7uoKjaBmV8j
iYQ8GYwbXmLmdu6tifQkAV02cIcGwpmk4mHjO7u48UHZgiTBsCQJm1K640OY+gJy
g9WDjEe2Ux2X3wPXAhGvnzS/9FFoo/hBQHcDtec/7hlAgpZQkmzVXsiX74CY8/t3
j2QD53G3fUBxnT1Zis1XORw8LKXshNJWODFaGKubDUI+bDclSRASExAXsjCE32Tq
D1Vo4PEMrSnZt6l8j7jzGb3Ur6nUjyzrx7T9u7yKj+nekFljAmQ47xXZlKlIqaug
wPrDxypEcaliGdBEbrxGzoCMnOS8wiMmvuqfmOCM0VXe5ziGQsz74Tlvd1Fmgblz
E8/BOZMNVVD2z8S5mQFQs8Kzi/Vmq86edJ+mGv2CkChIoli6Vsdw+nI5iuzKONh5
XHs2Na5y7BbN5rQZMc7ba+2i8gVFc1s034A4ozC5FOWywDakG6g7DSzSBsHl/eNO
m9cK9XxgFN7WQGYZ9mxpMoFIKwDB7hu9wOMDVpi3jY/a9X/yzr5IuYv6NgvTl+9v
qIgDzgsbUj3F/3UpiMOjKEmWaUHBjnkSPM0U6NF8r5hAX0QR8fEZQxtdwUsaec0o
T+FU8T+555W8eO2iWo/R89urZk+mkH+LvBAbYc/xRiz7B9CuCNzFxPOW6k+qhUK2
eQGBg067WQdFzdP+FLRYkGbhIEaduBteuSr+KcxgTHBCwbA69k7r36s7CB448fxv
aFKXRFg3OSVgSsCITKgZkaZQ36E2yC+RPsBoX/YmGleYtUqzhU9S+SOVh6OiHjEe
arpqb1UC/oxwGBudnF7auq9YZI0XWPA7P+EmYcSEwy62oOEzO3i42XbpapFfZ+Ks
EcY7aeBHiS2us8u3dYRKmwbpF9mH/DoRxX2rfqKjTw88PbM23BynHf7hp75KSHnl
BJsS55cI48isJ4WWcTT/NjeokFRfXw/jfBFiNvmWlaWoXndx3FqOHPKP/VPntlBC
bfyMpxQUkMZlWZ9zNFDDxpLVprcL7RhsjdfsR11SBb5CNy70PfHtEj9SJ1aq2mrP
HlM2LwB52+MHM4poL4VH+AVk5D7kfT0IGxuNtkp30snLsvGHlENx2M4kIgmY4nYq
ZZ8f8DS8OxXBOHV7POwDci9BPp4GAFUOgHQCZHAsxYO+cItKW/iUD2ol/d7B0JOo
2yvgVgpRHrT5ByKtQz0wwEJGRo0FOZyWMjNZyVYluW7CeBJTT3fSN2Epam0Qg0pi
lWCN4VWN9vCl0ZZU76NCsRu68JengGhalcTnFkTVw653TI5hnkIKwj4w5kEq4ES4
vvAuo8dbDXVHwkMJSXAxog75hAlPwVTwFgBm7p4FOMDgUfZdKcXUVMkNbsYT+ug5
thDK8IzYt+CDjvxsiYhVsW62y1BUURTq9TEc8Vn1Rfj2k1e1op1S6GQq/7idq/qe
2Gnm40td4WtmVd6X3t5jM6bogwl+9zgQkwA4f1yjoeTs3+TQD/sV9TY4Rsg2uElR
irHesknZOq0HOxxYe+VfoAMGMpvbobN4deGkNSI8EbkKER9U6EkVCIpY5XVRXd9o
EXA5uys1WouYPg1ZAKAIPCSCYtdVhFBticGjP5K7MmB755A9EwZMGf6CHRiug+IE
z6LDdf1XTYiomr0Tdw3+vXMs8TbhOMubHrulxTMVuOwW2Do05uL9/ZB7D/ylQlJg
iZEFmUDTmUsWMBMMoyC19c7ixieITmU/qbMVrNgvIDdAu6gkjB9DaVodTB/ffLMo
Xx+8nuz+OnIHO6GpvYclxH3RyCYWN8D09QCv7SBoSJBh2gBDOfMzhmRao2Zo4d/X
KiqERX46x/H0s4o+/6nz4ipCd5nobwKCmw+b7+w38O9X+zepE6AhzBPgIG3bNmfB
Euk6BMiWkf4y8qMt7w/+gRmgRBgnlhwQZTIoA71ey1Nns/z3BuEQTQX2zBrhBFcW
ydNjfLgMkKT+UdCp78YFptuqnLaPzj/6w89c1WTlWDiqON22GM776nNw32fAar6X
E7UOVuP8op3GG5NfnbQgMqWdsjvbS7HIFrK4urbWHFV+hpr4bEtV+UkiHuJSpOLd
5SNDDiBKqF+xgjkyaMbp5e63NiMaUOxkmcLpaQpsqAgiBFR7nvtwSHfl33krovni
tL/raJr8GZq0Wrg0tokMsrk3j//kvEfl2VHNN9TkhWNhWWXiBKIJu5FVmzL9Qrp2
9NoM59pOBn8oFLLHfgK3WqRPmlmXBq1HzN/wqPjTFbgzpj+HIrooCtlh4nX5d5OB
lao8tDHiA/kA4cCOAAm8wfbMAmVOYX0dTM9roeUnyl73hf/khsk22TeD5oT/+cb2
T4MR4u/3d999WI4JrthSs4nC/83tgmtEbo1edANcXotlsx81FWPcyxVPbBalpQir
fdpnCfOv/i5fJjk/3uagHYEL/ybPEuYymqW0x5719bQ+nA62mbQNHnmcAnMgY47X
ClIH2lEV1GKyXYRb/ll7aNpuhGAPawc+jLlDe2CLzzuGaP+jwvuwulYfc092LWUT
JEcMJNs5YEngg8W+d/Bjb1wsK0YKlEo2GL3+tK8qSq03fVk++JDYHxODbg7nJk2e
8/uxljLB1ICAaXlrImxEkCkLeLetlrKUO07q38U4c6IOty3/Tp9PaQr0qeZgiZ94
7ofE/7eYgpRiTzWbBqbN5cVciyOH9wATzykuiRwXB/LJsxcGMkpl53GWAVGyoWca
KP5e4HRCRsyAlo+/10x98xxJ+HwprPz830N87rsB964Ht2SL/1X0Bm7IJnrGo323
EACIZtLnlfPeU8Vkry+1PzzX9DuFPHqdAGrrHy9v6+SJoNElV2MtZOpSE5pQYW5+
uwICT7Uig933DMVv6ZCncctBtUH5C2KusTyV7mEEQ6w8bLOuiHGi66fMDNWpb/qW
/VeIpQkoLFNsnKoVfCzVFiFPIwQhWEfy01K35IxGCWtcLO1MBGvYCOoyMox91aKb
m4pwx83TwGqGqufZ1C03rRZViw4DIWOo6Lz9Y9pOkVSa4cdmE23o1OcSamZQ0hJJ
If07m7iwnPOHAyoIhmD6d8swpu3FLCt4TXxeSxsowPxzuehYc+NNwxO5HiBc1oW8
9VEEQvI9/3rWxGn9pzSw8jI1k0No4DWEV0fVly1BznknU6MY7llYvtkLnzJE8wTa
3dS96ODxnFVduklZrjd+aoY8tdxZPagNeSXWhcG9JhOKDzp3wNn03dn3pXQZNV3z
uYCltoyy6t0n4foTEPpH/CGDqyRtH97YQc2ZH0P43ZiCE/KjkVVmWbHguQgk8Dd9
kADPIkuKijyrrKuAX+G3juuP+5MqB9xsUMXr470NdQAsjqcQs1YGGxcuGX+JNF10
h3YIQ/5Yz0A7e75Tsx6m95lK5SWxlbeot24frlMyW4UZ01FYBoeRLTWraMwhyy9H
1jnxlyj3KrtT9FNfpdUyFvIJQ4puS0Rv7pJaCVDgUIU+W9WG+JLwPu0fku09FUjY
qj0Ozs8kj6L6Rtd8CRsyOAEkctLJxbz/dfA2VFJ5ZHbJA7TaE1nv1VjHRxuxNq4e
d8ZbBZBrBTftezp+FabROAkrJ03lllMAXxBileTnZ16Zj7Z4NlgG8X4U6AO+3gqO
1jr9nYf3fIDupvPEjZRQSiRn+0+POdj2Sv1b7SLdZHmaUmJTx/chOEbcu2AznBwv
gK7YOh0AytF+QhJmLS6Ei7Wr2f8znZKwtcyktpfULJM89NjilELDmZJOxf/ThAEW
JQ0cj6QWAntNTyPCKGHD+evxMq2uFM9PrRW+htvqVdrMDxVSHJfDRIrGLk1rZ3qF
vEOfRLtyzi2LpTs6wpP7RYrmaXmU10sfKjodxRV1JlDBdzsxj4e/a0Z4QIuwkTdg
YWV2agX9Mjk+snoW3y+dbVHLH4RXvJ/X20wOpqSECO0wDEoSkXBmKMAfFXuf9Kzq
TizNVLizCLM1xVU5i/lXX/kgMpFWyazCX+61c0ymwO5Zo5FQrCC1ISMCYC87UoLx
NhNCWbJG/zT/sAfxVkZ9SKuz6rl6yuv2IUICk6BYlmD2o7xi8HUfHAwyEpVQLcAe
JaRnuWkaWxNxgE0YnYK9f2w0PZzE9HxS7mO/E6Vn43Rz/DM9xsDn5auURUNZy2yl
RdwtVPM+iSIlRlAN8ig+3/ZJVlSgqh/Gm34fsd4B6/i8p6fJN5JeuN1Bj3XxIits
2XT7FUWq1y+GH/qj0RyxLs2jvIe0lDLvjHbZa8/22H+srciqqzK4OVT9xcaWfe5w
gFuB13wyYNLBjt2CLSvSyglFbDJk91VgdLIZqjrMXOXkUbO0CmeEMUlPbhf1HSpH
UjbNJtweLtcIIfNFP0g35ex3LDEyhtw29clxKVbAeOf31k8PHEPR/ErprR/oUZtU
mz9vEBcO/HLm/xgUiU1l9GX00cClHe0XAvH3e0OfoRXIFNVSNs7EoXZby09vux5Y
Ly4aT6a8DDFmywVctnqzyLISKe7H9A2g7cRiX1niAdUtk8JzOKD+DbxQwEvoSHxK
0GYhi1YO2DERmfH1DufHa9lQP9IyBy29u0H1qCE5uapdkYjjWcnJZcfHVPeUal58
2e/ngLFqKGxh+NK1qoIk0FsKj58mpqN0o917jxR5Vbhl+j1lypLXqxK9WLryjH+E
a/PI5xaGXXDZtSTmDRJkDUCXD3e41H9yF8vRYD7YKpGmJH73sfU8s15Z9JzXXDMo
33N8quMb/MmduiSgDrrC9jc1MsQxSSE61eQPcz9ANjxY2g2bQlEtDcDpClfh7ATQ
KxfmiOWHaUSETlsjsiEx9Mi9N8azoZwr++HJ8RssPKbz9CXnXw7ZorfXL+rT+DKM
hF0RSE2GfsAajWYDwixB/uiwhrGafhClopiRjBLlEY+Mg5QSJaXWq0aWJxxYtn9c
13E8yMRfh4SyNdmgkgscAH+wbg8XrJcuH7R9lDdOovIwwDKq8vyqwdW3SBwjn/ap
ey68ivHEUvtdZ0aq3CbaRYnY5S5yXnFuzQZtPhPtSFmfV5co2bR6OV3GPRy5h2WC
q3qfknVPJbkEAYR9nMurFYWr2eytHhs9+7aIRx6OkHTvTJ394vmSCiresAk+ZoV3
2Vx91gA/olCC7qTWlNbXK0/VxXNt4VvatbzNpgcDikNWZgF5gO02TXAoq1nN7NbX
nFrcakeEaZv9v+Q0R2vSxYXJyxwhsWLv5w9LlmVxiqNo7t2s0ZjsiZxBN/hJJBsk
ZsdnDQIcEs7SFq4t8r9LigBRyOG3wfsOoesJo4xRmzvhK5uOu6DKvplnoZlwAlcU
55uAq0p5hjcDGi+b8GjDwNhYo8+sMrQhff8WGmlqK410zIkto2oLRDJVoawYoatB
6u9yhY6PbHW9PtohvvqwJCm2T4fB9sSJYDohFABgEPlJdJzrgmzb2ims5dDe9qr7
J1/urSH2trnS4RY92VWcE6/IaJlPgdWzuq+5JE3w12gn82/qzLAKG2PbMTlhV/sM
Dnz1QCavLubPpa/QOWwY/E/zu7o21rCYDNBYIUUmuVPW1RrEYQ8LonWIA6tzjr5n
Uiuqne3ckQtOo6RZNyFuIctmAr26PWyK3LchFEaR9chGW335Sb0Zk04Xt00nxEdH
T0qAS1HSFUBph3iAnWDK4sBS0jEcIQrmSL9MLZpOu2VAFw0UNMbO1PWzJ8Ccy04h
eYFYCw4vYMGxLStRrDLDQQHMeWdLBoefUci/CWIaVoZiZToxhUY7is1WvJ4bSert
4vfxPIAnxi00e5KwgVTZ0pAPKySuC6nZbM5Cq9vjNYlc/P02PXeiyG/9NrefrT2K
OFneSxoveDUgtlVppsfKkzDxwaCBQqUSc1neveENtQC8/0lmq5ZIOJ2iWbbCue6A
jYrFE14H0rlVZ94adkYuNhEs9/7KtydcktoDN2MZeAMfQjeZGZqPMGWSWsYfUNUJ
CVxByCLIvxKB2Ep7EHBbF+/nFXwEVBmUNa9LNPFgxDVxVW8D1JMTVaG7cn1nfGEx
kpumdZ+luVwOlGnrmkZAM3mVuwirmofMOyjyXbMqJNZ2za4metkHE0YS+HW2R608
0KnhpgZlLf88osQlADOsMcVAJiIwBIAb0S14XhbKj3d4RYVA6vrTA+pe/dk66abD
Vj0GA5YFzfwfVxuly7ckH2o2/5Tisy9iiSQPMax9mzKNiDwnKLks3iK05TJyVtxO
LjXg8Kx3MoHdmetfTMsx41LbVFx4La4ITxYsdQJvU0TcbUWqamSEZ340OY5QPRpI
yfS3a+AXzCX33r+2eAv4UjhIB91Eg0A6dx0zsGw3ruZvqDvX6mXRqkjqx+Kt8o8h
4JzxorhllugwkrPjWXZhb295E3WSBxVNTp2yvd2FI0FS30v/67EHfkXa1DL/Y9gG
HCSLImSFaK3zeYnQsLlYYqlxtjbske0qX8ZJaJM0HaOXm2TnJo+Xv3pIbJ+82lUn
O3qc8VSj3hXC89vmYToJgbczmEHYpWTti8FTmsk46WgYPZMxNDwVo5tsGBRHgEKC
Y2vXXdVIU6gvS3A0IZfb6mNgTtcAWs6+J9Q9Sv3TIcNY4wJD8Q7rpLM5oW8Hnfnn
koL+nV+ZauACa3Q4DKRN/DgqPWOy9qdKHyJ/oSCUZt67vfhhmjGbJHLHlc3H+3Hs
K1eT3EIQNnBv+KyhICmynlrC6ryHIqS2vds3Lv1kd5yfMl9Baqjfm2jHhmmzW6aF
e75ZT8039s9KJ6TVE4HOtKEC4A7vRavITYHKzLbZ3j1hgP/ONwJDlKiNWw/7dE39
4+sekygACGp1Py8r9ytjyXRunK/vWokzpAOjrxMMtUy2rwio6ubBdbf3vYtsZ1nB
rWBZftC1S2IdBMSqUI2wB1ZPqwZckffj+L/NC1mVSCg4HJ+YZTCmT5G15tpaBAE7
IVjSZfqLXH+4al7vda0L/uD6OzTtFlxVaXlmb7jrK3u2UaGx3G6bsgahEagIGI2O
a0dLkKQeR9W7GaKAA4VavjKwPnEofUng5h7WyLdUxf3Bmp4k3PIFgaZzliUFMgoZ
KTVWdN5qXeCwZ9Sm0Rf3UtXCfu1y5Kd/PErzR+THHMCf6Vhu7btbPtVL7dlkCyqZ
6u7vC/OAEk3kIMcQCV0O8IxVxsZlfjM5c0JsJXQf7H4xWleT5lNc+c3zYsr3MExI
o6q5RJ08JlUipeV1YD2VPpv/SlGIVrbVrLqqwM/7qbUr8kUzp5xXUCyXADL98u8e
+WdmTkue+Zho+kiT0KaTdBYLeQZQN0XF4pKi1S7siOpRd/k6o+aZ0ML+wu8DVM+d
GEQOxyitsirUf2HL2pohDPNbTUkRVm2jlhj9OIVz3W7Qk1GISETZC6XhN1yuH+fm
6P5F+YknQ259qYWqeZB3FxxhIr2ztWIw1ablyLH44ohY7uNfJYsXmxq3OUFdvWjo
E+yvOxWnByOTOZrmXb00HKS5VlsRxTQhOucLUqJ5IZq8Kra86gslAByp1j/LllXi
2Esh2ICOfmZr7ZDxfx+7iDPFEqClLZRHPgehZgrgsrWapqJej9OQhdbh82R5M4Zl
RomjvIVRVci8rZ30vOkllGq/mTk6xyee3fzqcIV6+R6gHGpq3bGwPdL5TBIjQ45W
7RXY63v0DYhiSX5q1PphehQ6hwhRxNWUk+bTQjove04ZJ2mVzb2daBLl3ih4ddvZ
ebhvHLrde8oR6gWTJL/00jkCaQAg1Lt/v7Rkq/RdEVN0+EPFvWsJhHICOA6romCc
T2gK2jbC/NVv499zo4IVZOeQF8rZk1yUfW+ZcMfpEOoaQSFtmkE2PcSpL7n8uFTG
eTdA/o9D/swDt6nSqJrbSWgGpA2IzFp6WoswICs8zOGKu47C0pFJycwYtyE5bOil
jZEQHBVb0/jcVbhjcgmdjRnU3h6AZXDfjr54JxFDt0iuXZwhPWdHgezuhCU21IA/
f18N9Ib1ev4Lu41G2e7lZU3zFQmqONTXZ8deDMkNgobo2TBs8xPQjZRkoot4SXc6
sZ6DqGc+IYPHicqTVqINJPVqyy7y4eGXHjQiud9F43Ici02ergZYomC3qNt/xM92
2ztDqGTEqCWqiGAcNbDdcRabRduV3u34fji8P0gAjxGhk2MrhnPwwaNk9ZaBm0ln
I2GvNBerKbTG+BjkV3nV3i4EXemM670v4QMNGkZLxCb3AhQaRUOfWR+mbwej/qG1
/RCAdKW9obnD1GyE66jDsXaAEfn3MTBWpDLtB7I259dz1FaqisDDD+SXD2mKMPoL
82zKAMtvq8wy8H+V7eo7y40LuXBJ1fEj2crEfEKbuO3NAE9exDTfkvfrUA+fwly4
5ip7jf68pJyRq935I19u1niaTfTJgSgJmZkQtUODTAHqsOaiXrcZFMQCKTgvbdMp
L793UWOf+ITtiNSoI1PKIc6FAnqeM6Vq4HuP7OQ36d0FheRJf11xKpFW+nG2PIZG
9gBebmeDz4C/zA5hbjLQAZCEHRg4FMhpFlxsHxwdeRtNTKcv0O4M5STG8/N0fwLL
N1+p/sKA1TJQOnN5VlgzmfwuZA+ItvRbWZwgMv/ZB4AadYkcXnlwhaHMg9r95CI+
QevkfBEBuQqq7KmIB/f8t5Yzc7syamcQ/1Ws4ENYGajt35zoaAipmUFjzJicvYKY
rmiOkY5Gagr5NzHE5eJJhsKYYgUgXnjASVN7LcZ2c5bY9FhZmyRk7yVYm/uufhx5
YJYFOQQ+IoKDH+vvneoWTXqpSI4WzFaPp5QcH9K4+P/nD2FUAiL50CHLJoDa9IvA
fDqNdsqcGRYjJnGNPQEuiLWQq9up/xpvcIECuH40GKApsh6IiTJtTe3p4hpAQ3Jj
7l2Vcgzm+5aDanOncJSUeKNwd4edR5KBILSK7HjaTxqY5m1lNsOjejTogYf4ZU1m
UM39+6oZoUTiQnvQyjsEJIlx/7bO5NmBZdccGiH0/twrw3DHTO4i8cFOvGuphISQ
Qvp9m0ruPl9MVsxgOlLeCRmPt/xlYtHZNBB0+JY5Pjw7CSlnqUbMN23hl9L4rXSg
W874GX6VAc55nj+2JlnGPXY7tO+oJJZpEolokL6qklVOHzVQJUvfO3z1PppKqcOh
1hXHijn8ZQMMEH6pmmTxYHrVFv80PqOxgnFR/a/2avF79ktSOAN+Bc8uclzp2Lo8
aURIRdOSIMwZoyrdBWvX7s3RTk8/yGuOOTKUuydSV1QoeO1TdDX9bCpysNiam7wB
DkzLXHqU31IMHnVVhRt0gJUtPGR/OyUH5xf/EBVJRw0p1mFSYczUpvWWmERAt8B0
KgUXu5Nh7dexI6A53qVGTJVW/DEkAfdBpazSKWp1QDKOjbChLOM6ZE7iovoOjyVh
l4aoBy6dXoaz/gVPzZjLmI7JkM93RDaCtzzjpm7Jkq0BfQhRD7e5mINtpgn6qiWf
IEbQvpPSE3pxZBq2qrUEAs3o/fIkpuTDJBNCA/Izu4S+4VxQiANPk5gwz2WuR7NN
zpXmLFSAUoe/JNqsKuODchXolip9h0az3GSVQLKIxh6JtLvYA1Tz+8pRfSLD+g9e
u5X11T7W2ogS2vkOhtLz2N+Y6Efly0T3YGh1MdHeuvo5qSpb9UCnSbhnC+kKur8C
c0dbkkj5QYLIT5RpyDN1NPFtIMb4j7fZvgCCVIhNK2GzEo6tX2rO5XAV+HB4l9x1
0x/cUnAEet0Qqfsz2LxA6kpOAE3pxwsaBkTkfibRHPqXNN8tIULHY/yH3UNvmS3F
JuvkXZJGU5wmDON32/ju1IK5cAcbBDBT1g9OXH/MmslUZfm/7Qqc0JQcyKaxtQ32
WC42u5RbnCi5gsausuOLy5GfiPNR3nt/awGDUmK53s1x1Uwx2XlPf08K0LulOQ2U
ku4wG7HtziERd7hX08ILgV2HBnnrn8gGtV8DqdpZIxR8ma0a1OO01+GOUa4KbnRX
SJ0sMN2oqitrTYpeYgE6/LTGSAgdny/Aw+gb5GOKQwDnbE4CCR+eotSJBaotu4Zz
BLvY9CZopesW2mcwD1i4RduqYI0qoC1G2s4o7YiufRZNk15jmaU6yVDoVNKDLLLN
G6qo0LJl5PBn+KRAzWZqw29ArVdb8qzUne8UrK2kvCG9Q27WkqbNnxMp2Kie0szy
aY/YCpxiEcz5N8XUV7V/4UNVFs8E8aygt9+yz+FNOEmYgBePR44dyXrcHYYMUQnh
yfUAHcbpqFxlczZBLWeJ7EfP/IbOypMXkD08l7Ocs9fcJ9DzB6jG1iudtpe+10xN
6zt1tpSDw/siSz/6Opi97xQlDBbBC83wttU/YWkNH8+RnYJBGiH4WO8/N05ZiIZZ
4L67pHF9hxSC4yeBnIlIrAgeX3Hv5Juei0+eY1jLItTYsfYH0pmumiOaHfkE14ho
AioCyW8sn8kWzCfD6ojkhecmJmeHdOeGqdUdi+d8xV3vD9GzJqAXUJIT75UyukdP
/c7/uxba2FKd8PUF/+SXYqIUwWIvimF425Zwp8+ByMuiE1hCxqgitbf39gf9D9i1
YoFUQH2RYoQwDZAFlKqXBUmjJXikb2mpKUu7nIBMe8OSv8E8O6AcoXkf0DzMoKxY
zVqt34oG+GW2eWJv9DiTMNP1eciXq4TJjZi9WpxLhSBbyYbFLB0kjw8EtUKv1/3K
xoEyIObumByNR/CZ6fvS1P3mvWaOVOMpCIEkOfWtL3PDUT6wmV92DOInz0NBxVNM
F/gVwsd0biufpWOugtOctSAon2WgTtHskzWfsyveDIUEM9aeI8/XPidy6zBU3UT0
mmOQRMVrTuMwH66d/Ry5c2F0Ut1gdjhvDn0tI+hvnIdTIikEisooG1524dOY+f0G
KvCBmK96qGUj51dv5zE6RUMdAJ5+4g8QF8QV3TQKnUU4pOslS3f1mDu7ra5fGaxz
KH5JN3pH+B5bAFImNUv95QbiyVsTkvtZwqDDhZgLdI7YQYY2vR3nuWiAsbbIQSb+
CU8nQqEM8pVGD2iHpOOndQCDevhN6x0J5fgo0p+WYPkW9oRbA7AjZXNGupmZY+rZ
5u+WsqLJnGV5cv7DBN/hYgRZGkAPWZxw1jMMG0JSVNIkjn9hE/gkfToxvXih7/UF
cAb8S8xpN2oDIdBmr8uLE2+LNHniR8JRpc820itj0W5vg0X8O6eubWKvXg4L4eSj
ZYalJekUsMagtPpmK3sGu6hXHUQTXcWS7JoZ2eJnckGTQu4mDmQrm/Q0mkXfxL3M
JpobIn4Wn9HiC58gzeBIt/gY3K9BA4IBu4ypiNw2mMZgI9Z3pt45z2QdRTwnWY96
0f12LW1VfnXrGacah2YAeenwr+vDP5oZm69hdqzAK7+RER1UKyXQ0dkVNT9lZ8TQ
yGrCRp44EvN26yOWKq1Tve0+7OzmZhoag3vSOj2QSlRJ+Lvz6q/ZPIsIY27VDk8q
5Q/JuiaR9mZGp8PImABGD3PR3k82jAcBX9CVadRJlt5uZ6rr7W1qlCUoBnLq5ml7
EDyXvyLzGRhRSwsJ4bJf0QSBLP7O4VanLGsYX68A2GZDLO8teIaIeCgsfYlARWZL
O9db+p8Dy3df9WLb+Um6KpSx1t0kwyFjyxDvG4gFVYJzsZl9ZOXg/2vIoHTtxYuE
PBD+yIbF1nx2RJ270/Cm/RiJV3c2jWRKIfurvXgdk497RLZ2V+DcrBP1yQIZUJkZ
SiC6ujcp4wb+Ga24ceo11Rz0ER6nzo0iPZ+1jcvHYIjOBIDHjRdc35g1Ky/g6FYn
HdLvMyaGtCBoPn4P+DiQ5iCd+mLygxUZjwTGNi/mAd9r0gSUjnSQ9SeB/SLH1l8g
SW6/iQ/0adGRyVgmFFugWYr6UgEGizE0HPTTtsZTrWGrrFkxVFlgwtI8PbcO2obx
TjL4f+yufeQEVQobh9AlwsdIpdm5LGYIIUqxEKKsrNq+/Cpwhr95Zzpk4r1I9giP
jnw3eX8pLJ+yTgmeRyFCCFE4YSFpcFNrZIJtnbfEQcs11KNts7aRF6LDQvS+sye4
dRNXC/BeCBP9+RJ9qmSOQi681A6Fam6AkvoKLYvGuxIPqXA5zGeR/AFKUlqHjsrS
igQZ9Csianbx94zksocp00Gt2NTg/UP+C3YLeRXHZIFslIhfMpfcpy4XItEoELVj
7eBN8yxiliOj4Rb6FnLXgCvbbUpMgdeKWZ7T4XrtA/+54N/GfUpVLRAmtsu2tbBU
2MFw45hU36fh/3Vxy4cLatSVBtAhysTc25WcsPp0+TB8uTRu7t+QjUR+Jz6xe6OW
pg51y6ILJiWRiDpk8PCrJRvffAA5rZt9wheiqg4x7k9yGGCpHzHiMcu3Y2BM1uLO
HIbeQthyoeKV31KU0R98O1cg+befxqhqBffesV7Sgg+xGlxQylwtEUp/BhF70ojm
dJ5jbnvGr2e1MtMMHaxuK24yUUAviQU5YcNcGdxjYe0gwLJm8Mm6jy+Bxu0YnJPV
WtXtwY/VhudtkvESdukxIEmeGg2Hu8o6nqfjs9Jou1W4PVf/r4rJUPdRpfSOaji0
wQoLYqbK/gd734Bs/PkZgmE7u6WeT2DkyeyK+dPgTYUe9dNbAZNqaK8j2lj9o0Cx
voKldySssFACJ9cR0J6JJbpyZIJnd4Nb1HSP+yFOUZOzr6HSmSZwllOrg/zbfI5X
NyCE9AjP0CFJUY/DS7TIDXu7WWrcRxXpI2m7UzovY8QZ5+zIyWu0KvJzXy0LcmpA
uPlsKf90j399+PFw7aRIKAJCnZwSsU1YUSjOT0P71lChq583aS9D6sVFjaU2F0Vy
A1TYsGD1P/zqN9+cXMW8V/oS6Wn1JJde9qeXzJUrYvkvk4GASxOnLTVGDEvMeh6Z
BIS+kluzsjU21jMDF3TJWTfTjv/g3ufcTZB5tMMSvapyU37I+YBs7Z5UkQSp8axk
nvXN7SgVkm1yAQ/x+hMn3R/gGIETUmvRsLpml6GWW41paLcJQtyIqAnk90zj7xlW
Hb0rnZ6wn9qcvZkLxs0drHFOusFgKG31l5jOEqNPe0+Ct+FmYx1ixTdFPhhKB7gt
Iew9OjguT31bQeKtjlzrI5SCEaqqQrltBoyoaBbBeYNlWKJMLfjp79PNMFE1nsIH
tdjznYw1Wap08ba89zyaMANboIzZdlJCTNaTgIa2XIEfVQzrVpZdxLp2Rz7TnGrj
laOiP8IcZqgJj841NEzZJ3RdQHLDpYitjim2n/XGrD+JnnxdtaR1CXl3ajKyZUgT
/rMe8PIvm9Tf8z6GAIwB6ZPUjwlgQUBQUgTE6xXTfNfgzBkY5IRZOWRXiOYmZZpM
JrvwauYhZGCL088EHOcz/EJrtSQoeF/rx3WOs5ik2wZqceNuhbOKFDcQrtod6Dwf
/xxB32bHIO2gYv3BXUsQMQ1okFnKQsanwkdT7vYaVwWfV6TfsOXKIEJhYOTBjZ3n
0+y5/+FsdyCqLQyvGjKBw48uuM9CyLRs4E3miJIHJGfxMmr2vw3n8+lWCwmxI4NT
rYLs2Pmq6PL8X4/zcKI8SlWNMLIa8aKfdYyilozPH/127xoXw11PO88LUUW7M9+F
qYNHc0SG4uBZ9WfInPJPt6fOx2htYLftXLCnI+mX1pSy9O9DoUZyWuWJE1Q/qF3J
ZFZgdeZzjajcaUQjtDaTY1H51mLiB6fX4L284gFZYvW511UgxIWbQrvqdkUsgETx
W23Ann5tQlYU0LaBF6mEC47+MdfGJDTbEa5XzYJSg+wcUoKGComwdUDsLg/ebOac
M4fBhbY59HnByAAASfEGJE1fy5ubVVyK3R0UAIR+zWdR1PMsFUEDFP+UmU6AomG9
7S17NFo3yFDoovJRpmgPzJ8asuqqnQo6qTtlHnDpRZSkQQZJFpcrLUjq00YuyFPi
JhraOL/NqfKEDgaUyYrpQVeUXbufu5/yTIiVlyZqVD4ZeD7DXyvhiYY+yIouBN5r
YN07XD/TOwWo2ID2Ou6twrxx3WHKaNrKaVQkg2K58eI6J9uKIPyV0W9KVpvvjs0A
ei4NxdaNZtdAZg1lZK6t+OAL5LHhx5YVSO6CxS7RqXJl65J4XbPnkeDrV3oiZgcE
Jcl3PavENqCkfGIiLe3NHn1QQP4KkWeEMfC+eAZbHDeg4uUTbogkTyL6C5UImQiS
2njJGWu8sgPVzhnSLXbQefUnOqxWttyOkrghz7SKmPCfEuc1Pi3fVI1Nl69jA3co
L6L9E4ZUQ4Jk44YKzEAxjdlVS0QWT6ke0uwAFP4RwDw/GeArGBPtZqbqzFeuChoY
aKzCWChGDhDbUxm3oqbX4ZGbzjrBo8ResNTKd3GNWzfQhHXJpzrBtz6qO4awczAw
ENVXpYIJGO6fQpXxqXOYKctq/drP/P4cu2xDNE9a9UZh4hjPRCr2bSs8aTUmih2l
5YUWChOzpDVvXed99UvHwax91xHkRvcGHGLogyE3U3jYfBAef1L5G3Nu/WEDdftj
eexvlk+gKa6fcZDTEKqZzwTmfMPnCyvy3ChHvstrmv8TvgK7dlOfqt8a3QBjbdgF
lPZXxQVeEk0OtAezwU6muhjBz8ot4lUERJkPIpyh31M770N6cjkcjSs+iaoEiBbe
WFcZkLOsGBlUcw8zNzyJv0EU43HzGghqgx+T7ifakaH91fQQIWp+8EDchoo8Kdr0
HKw/pBOzTjEprTFdNiIWlbFqjNTXeFQ6h8PgN6l0Ag+JHcz/suzxHUDE8a+rxh+S
+lu2Q5ESG9IStjQmDu9qkxwi0fDWKx7gDWm0G1CPZVoSXzQsDr2u2h6bQ2osHjWc
R46a5p30RN0/QjS6sMNrKwPnj9ulm/ehYDDG8ixZ6YALkXRXafv++vOv3Bt9nGyV
XbplxXW8X1k5XY6uq4s3/tTQOEuOc0oMAFSiwrJLFEPwcRfdHYjNIL3cCL6uaLlh
l3VLT+vX+QQZXWNhp2j3HrdO3k52RfuB9mg1dSc+vphFaFFVZDtaq41H6jWozeoW
n2cKIv5gBE20VUvlcBEdQqE8uC0rTGeTaRbpzn/LOBCG+xd/zyDgIfKS+hkZj6Rr
hB9iBQtOEbKfbqJadwlvKUgAI5GyX7Df85jzwtPM238CJticKUixquX7xpKl9/Qf
lKQCuyNbhoZgXij09tO+bvtQj02ZRV3uhfsNWCxa+8UP+qYsskB2lERm74IOjasE
EKaguuOb6uDUuUTAS+HaC1cG/w323RegC8aDmU0H/qQ8cQxb8sUaMSAocJ52oa3R
U0w4KPRl1yM4vH1zqIGF+Hf5AB33oxdFIPeJFCNfLIdYT8nA1WuzCdFFavw9f7+g
ZjfkxICgSLSwonGV5XPEk/1hl7WQ0emvxkgsrrJYwG+VIEoR72Kle/OJe2gSnfoY
mNtfAf1Z6EJOAseEYgjp3sml6EYbxkqnEBqBU3vVnbuLrpq5WEvTbTXcgZpf7Y7r
zPpYJ2iWYcy9GL/+JXrtoKefCu44GQpqD4q5xis9eTB74Yv99o9RDWo6p16yS75d
K9mvdftvJz8X2PVFhAAbTEOMznBgYjvJ1dm1mcB5h5mvQj4cuqSM8wQfWm6W2kVg
nsWnJBF5ECBOI0Ta+uPc6SYXvZh6owyqEvdA0rie3rdUZtkPzOxdlYpD2SB6A9BM
+8L8VqEL3Cc9JjPkIUtPVZSh/pmG+gz6F/NO4gvjzMlua9LcHG+wbeABzH2g7Qvm
OO1SfGTuD2HDLvz0dBJeYOrEOWmndB11illiNsvWvD3onBFxWe71hP4ytjhOxzuH
+sLI7GcKPgstqSmMemuC8aWhe0RAun4F+dHNcIciA79FIq3nP/eb7NyrXxUDLLyw
S3Do6J6VOI6y8RgZKhX2wkNtDWTlpTi0yxCTzWESuOMd+klUj981B4JXYoBbFmwR
wD+vBk/37r3NX+nA+9YweP07aduL1zu2PQFnSu3q8YLoZvZRjgT3k0DFHWhEc1TZ
e9JixQ1rMFvcDthFBcNHHhcroftwCFd/FjgQGJWZEdA99LaqBICJPGS41Zh6+Oy2
L9aXmLR0n0LRu4vh+SOlKug2XNe5n9cwM4HWpzvZ2DG6d+ey1PfU3i5y7NoLi073
flUabJbpVOpnQpgthOZtPvOld3L8LIFTJwwYx8zBVIfEqqt/MViycgh4JNOAcXtR
DbP6CQ+SvQqfcGP5cbaTFg7f0Ch7OfYUygmhCzpWNToZMoP0TCEgKqy6XksnYiN7
9jedNlJ2T+/XqvUfhVvVteQ+PzyWx/Wwpl9qa1qPczaQxxbcBkICXNaFOx0LjHqJ
I4FjG3KEC4p4IZ3VLkcv9PKHYvreDeBWVaiedwzhFrs9675ZKdzFwo1i/eWQYLcd
QV2EJIjdbSu+w0raWm5Pw4ZsmlcsaT/IXup2UTFQiuMg4MyelKWKZ+qTdG3IZk0z
WYOIfOPxVltO73jC44rq7ZmcCzknFOEeS+3AensAO/ba6C2zI23IpmB3Ci+FmX9N
V5qj51LwruPXdNy4/Uagfrrdu0uW6lQI93ViPzeEEslS7v+4/ziGmvmscnhOXhSn
fPQUvl9dNJxDlYRTmRA5MPX6DeFEYvFE4ciBXoMyrd9Bl/guGBCdO/v8gb8d3a8t
kdyLCNFte+O9pf0JXFNZgix/b8w2Xm/rc9O6Q2v83z3qV/OyHr4/HUvP0QDJemqa
aWdtnomz0RnaIbFr8PP5EHFBPXpEZBavVBmarznVNB08SiwFvWDddAlXf9/4tu8X
SMhtkbygl9dso26Vr8yn3wSD+pm8gTltaOjzYBUh3NLoNf+/7zs1UoApExvHHMjy
e5ZZvAgPxhbkJXYQdFZoeoWJGBNkILZNyVfjzkiEVg7QYEBOYSbTZ2u2umfoR7em
1juMUKlCboZyhiFZXA5hhzikMzRd6m/WZb9hecZJDHqrO1XK0nr3BhPAeczS53QV
kCD90NYctA09aNYKlVjJ5eW404/r3IXHTUPZdaVDQvocxeS0/KHoCOdYQdLFCeGC
hojenTCQ/X1C2o1a/00InuO7MO3biBbX9VsxUz8Tl70zLiTx+z9eVUbC72Tzqb/p
X44f/DTWK87oraA2bIMYLUbRBym8CX9nYzEnOb2dEIWq/lSQoEWrreoo4UOSk2Ss
if2NZoeCdlj8SfddG00lmnkJmXuCp6dLX3AhmX3AsdvL4tcKPb7ECM0eApmjZZ1f
LVxqY4kFTZ/nZjYph5qmY30CwrNDlKThxhJMqBvKd5C45fjNySNsQmnbbdth/cOw
/2v4fjEWy1mXX1s06+/2+KKFka4IV+9QDGWWTzJoJk4KmRPEuqUu1FwFVXGy+BT4
ublzKq9dlwKIVcj1DZ7CQSQ64AInv0WlhTy4d4h/VpXFGS4+9fkqWZ4aM/RTyLVM
pitV5fYqNYZ4lnsnUceNLlu93mSVYVJ2fuOBjinG/KxEwJnLjCyG5tNEAJfUykqi
zjckpJVm8R/gRHoU04igBns8WGqA4EmNANDEj9ukw5UIeeU1+qrd0AVGFWJHoOqX
DaOsD4L8+ifLW+jUHmapAloE3P4QJzLTmJ5I+NDoN2ncQzMyvmbBj9J6EIyNqXKk
uY6iqpIFXVdPAzFDxIt275O6g1pwQ9vVuTBrLBfVq9A12YWfRyvPL+xLtgVU1v07
axzQ9T0y4KslpEueezKAzt+C4koTQ8cikn12ochhR3VLu3Qn+FocwBVngxE0gl/v
SP+t3KSScKD6/8WXIwAsjv/mcHUyGiz+f4NqjSdwloxYr+WrVfH8SOYfOQ6ZD7lB
BH0gYfs49iWNrF4+vIEy0UmoLD1D+F8HwW2PnyNoOAXANUP48Mw9oUjUEcJQ8afA
w5C/hDgklEH2xLKCFlFwf8+nlqcHJUyclCkNfbAvisV1RdLy+DBzqWmUHn7Ir6rT
uyYEQE11ASfG4ZdJxrLByFSMjv7Py4YWVkcHfarwxyt32x238peS0fejNfRo8Qwx
vUWN/w/vHXZyVc8VEjef4tUD3YllIbQPaf0VXzDC7VsOp4Jl+CVE/bH54WzxetNw
IMpCci3y0J+vvAKF3ubLRr8B9Z5zh3alWmnVni5hRX92JeVEAVf1uk9FEdAhEYNw
jOs8b9JP+78CULupuEbzx9uNtdiH/J9MTl72wdyhz8EHqCQjndofdPBLlqhZ9ygC
hBJ3VwbQcpokQLViEG1Cz2wmmk6vk/GIvAzt66YlNJVHXZf2AhCTS/tC1jLhrMma
Go/NseDvs/Iu7LG84uqdbBGIxcD1NLXRpY/iUHoU4ukROoVfCtOQ2wfaATZN9f6m
AYErn9cNJvS/kHHkNv1z2jQs9/WG24pv7APS5sA762ZXe41eigE/+kVLDUCbvTxH
AfHke56RJiunxSZO+6EQfrWnBnAuMIWX9pgyxRJyLmepN2J2VsSQGOY9e/QuMo7v
Qg/ifQQjW71m5ihfXprvnpXleojhZXFU+Rqs/RFuOGkzsPxVp2jNn35dC4aafk47
xGeGVx3kc1d6iiCVPgoFONwhdkJY5I+WONwfOOv0ZKJLkr2qMAgTCSbfpatnWTfw
9N3za4a1356fOiT+ObkKFnMbYl9yNnvJT48XjvMaxTeu+FMLGi2ffk5gPqmcLPJG
74t2qWiYUewvcjgh8Sfd4LCnI0a/bdY73YF+rHeev5Lef0hLZO+P/JvDd+M8t2+k
TaydzMUDIP62NNu9cGzNY03lTHAk+5WSPCapkWdVlehKM6ZzRWKzemAdfh0Rja+L
CxeWyAZIVwV7SPP+eFyUq0cKIONzAyE8+EUjM0zUAUKTpvC7kWR9T6w/BoyiDsb7
bGR4gHP7QPO4Nxix3M8Nf465epWzYHqsdOABeN43oIaVuowzZfv41hr2jwNITbz3
ndXd3KSSRzSoJk5rteOsQl+83Mff4FUo7AotXG1j2arEfC6MWjya8hsS5CrfxOUG
/8U8OaOJxyRJGDc0Wsz88Fr8yQKR4qjILeb4BBom9rXLH0d9l4+kdU12xuihSZmZ
3UCXsWImEXowFEDRMoBNiM0HWyzjZi82f2u99M47mftkGishEtJOVDvk5k724MZ3
Z740DqdvbKA64keJQXEbjpT5Ims82KEGT59Vo7gdUs1Twsmm1PyMMONxOKjCD7Fk
RI+3TS0Qgv9/m+nmxO1SI6xuax9MA55xB5i8jZMhJly7e7QeVJGCryrRZM6bEHtd
d0kJXZ4jkygOOs8ibn4ssgPXwUrbf5mnxGLIMvFvFGPwqWtRPmnoFePmdsHBLMag
QBp4vnW6V6pvtIAcQiS/GbijZPiMZ102bGY3A2xlfTvWF4NAJ3m24f8uIBXmjOr5
ED7RDoNwat7zRinUJgdq85WIMJ9eabuWGoctwo4R7/mSMiVRWpaD1U3G1y3z3M2R
NN+kqoJh6AKok8TSwxFbE0yZE9K8aEQeT9C3slIKjqqQ6i7bOzFsvFB5elzgGkz9
ELFUAOENCZEx3Ezgw8+SyZrEqQCxAWc2gilvREOPst4t28JFRaCzS4EDSzJ79Z/u
SaVieV1uWbhyCOtIkzK83m7GnShflUmqWVPh9ZqytCiYCEEymbe4fSE6ku46BN6w
2Tj2BEh8XXFtF2wHbXWDVYUXEgcpknuPyCuT3+1wsI33ito1Ylw2RA+i+1ZGlCfE
0g84hlwiSGiaBHvjnDneBqq8IOuYw0b+SouivrW8oTGUN1se86G1vuOojq3O55NX
riDAcb4T/IjnDsCGbecvB/Qg7IgfZ8b9J1Foxynvdsr30s1uNHWjwVfgkyZB1r+O
uJQydM3HuxSaKmKag2eNB/iv+wtOyKf8Ln8s/NoaWzligSwDAhyY6bnyr2Rx51I0
QWxW+oUswQksErgNL9Ondxq8OkPgXW01pFkx512XUukO4gddJAojgLvB0ioq2ZVP
nwQWBUafFxZFmyJAOiMUfgyQZcf1RrpSdmzF4z5Be54s3g3BrydtN8Vs6vEdAJOP
5Auu8iubt1qxtyz9kJNIfJENaX4/QQbAx0ZSpjudFB6m779oCU4yjcC7zr9gZier
PvdNDmCwcCOFHOuSJ3LEuzdVVbYHIRTpXW3ZpzF1SDKHXfOUMy6Lk1gJRjytjVzG
bw1Svt8mh8txgPB/PTCNE5LCg6BqSRNzUXdeuUgsTTSbwkElh9WZdMThkuKo4SPm
RZlBqOF4Wf14Rd8448Zjsze5KfPHQKQVkhXXwUbTmgEo7C7W5gD2JSZzEtZz/iRd
V4rOA7KSdTxlqZIJ0NfbqSCVM2Aew9jqzEnIfPLuGM6nwooHT4il94aZ3z2EFaxt
NBDXWVANCB/zDJ5pbj+Zh+/+8sh0LgLBNeZAWYYUQ+zGY0kA7E3Eua578I6RmY4o
PwQvyZg/HKv2iFS751W9MrFv/JaqiwBBB44vKpq0WfmEN+qltkzWSNwbR0Bd+UBA
1kT126pE459XkI+UxV9wSs+z6ydrHt8rMFkYioG2L1JgDT5DCEU+rJiYU0BZPRek
tGqNiILOAlxAhcUGZRSDqEFiN7vbpKfxyxIf6wfs4pgY+ZFL+9G7kEn14Un8liJx
6nwM0HOteiEQbtgdqlfbpPqQ2Db5fGgpenNmSTF4fESll9VgyMppM7mieMXMqS2W
DgA4MWz9LReNNoPdFwNJ7ok6Z4d6ct6W/B2LPTxOZ8sQHlkJHuXZxDCb5qe2n3xO
m8N0W1nFHN4SB6ZUN95JblN0spkc9Rt0sF5TCAip26BhgBMTh+RyMBOio150bT/m
mSeKAXoGx2Yupyc6FjIv+iWTopn1plzJeYZYBls0VorD6H0Hb+YfyxeI5e1RPbSB
qsU4baNEn8hcL076Tp0JOGDZNl38kFznTHkh1uWdozFiYJOZm/uDuQvSPuys7W2u
gI1jxdiPOzbK1ckbkOEkMRoSFA3qTycxAjyI+8jLrveAfXl2ZpZUy2gO+8MEVFUT
emjlUkpfXxdTorISNfy5TAnHzI7p/Kf+ZBjjHkwaVd21BxMfHbZz/epRMMFjOLNI
NEkOT7XEclrXwuiMLXekGO4SXzZX2EqrpI/6/QexxKcF6bSCT+BY41ZNAE7EsVMB
94/DjuPFKW9ECw5TLE1Hi952jc+DmjeeQrm/ZZld5fLp4R6GB2gg39uWiEsWYX1m
ThKncbWrA02OTSSLYJmURMuwrlvPG+U4LOH0OgdSNgsSCliS984APlUYJZa+C3bZ
qcrzg5tTif1cp3qelyj1+uCdf/Gx67GRd/Exk9KZuh8NV5tUPt3lcao9vRH9r/6F
IuQ/sQbge0QzQ96Sk3oRzlFU66oQg6FNaP0mLvh+PHYEOLsBjqLTgg0lqcG7otSE
/uKx4wxGMnG7SzJQ3eGYtFvHDygfwLrdcotei0X2PNBcnIrGdyistzmzRZTnwbeC
loQYvcswjk5KsVfjNMGZz1X7Xiq6nFAxlRT6jTXzNCaQ7jECijD2kGm/NA1eTsTf
e3n72wgK+YsjMxAILfFxWCDhhJxmJS3R0boU5HblHeqnnMX5HkmOrrOeE5oaNmuF
dFhIuBbSaKXbT+nsGQb4Ox9qLsNhz6hxWbTBI+CAZ46YQuc6KZPFfnbG6quelbdU
VaWHH2+h1uYiIRCs4hXR6NN70rIcBQkKRvnRguhS7RHJC6/S8Ulk7O27Khdi7oU0
IGz+65sv8ewkmqmvr80Go0/Km8BfYh6PeryJEhqCwdMvhwvS/30cnbdH1HJN32t+
J8XHW6myOc552zVOFPC0MyZ24QNS7k0NfupxF/1bciQu86TfvL4HY78z0itd1ki5
N5MXURNGr6OgQojsq3nT1XetdwOXpV6AU1DeVmuLr7jMPhS/M4mxK0+d6FZNQJDa
1W5jNiLNXEp0FYwTPT4lsGxsXc5lXVdmN5+m1K/QCkOLtWfxL+fYRO4Lz6h+SsB3
iu0GFfipUw4A2G/W5FNpUTk4zSdh2wN6nIb8NuVvz9KLuHCu6vYnTsDejO0I1a5j
juXFx8mZiZFGU52JaLn5TlLB3YUgYX6RM9ES0ZcCHXHl2d4u+SOXIuQgI94c/wbR
iFKI0oJXQSLYpkW6COBPy7NcaLCrE1dawyrnapFjJZeWc5/7pIblnp6zbInea9nd
xe1IjF1Orek8Sb9C5GqLLSKDFZOgZNN6RG8Bff00bl3JuZnJISdVhNB7NEhyyFvf
01Gk0T12NK9lcEridbnEXsVwiLCuLaZidxoxOIkhMx+Ng7ON0Zj+ppslO3GqMvFc
d26MV/doqSrilziep/APM7iGLQnUujjzt+JAXWkiUCPeCj5kqdeAqOzRKyfWX2rS
btnIGIKngTE/BkuGmipP/jM2dOmeKBoryFOBblBqoJ4qQsK3qkEsHOrFDeBjqbkz
y2agPLtXTMIYZhlxtWOM6ZB8xP2lK3xn6deEjTZcs8HofXDBuV7z2hcpc9CgeWc3
XLxOM/8DFlVs6ShFT7935FqUQFZAge3lPskTRyTiz85lLOOVNpPoCn5AvqLUHxO7
cVFGlli/t7NMT0/GnWljSIsuSoyvhkX1Jot75jFGZDKrlZ1W5XEPFTZ6mjTDX55L
m6Ac6RmqqSZEuaZ/I+WiTpLIhPnY7MlOqb4mcZF6UrzcezL4RN1y3PR5M2H0aYfP
2j+gkQVlU+SLTnXc+iYO07wCYESZaTe/kyihBGe4G0PNceekmJIp1a81M1M4SSzb
ApDMyMXBMNo3IuTItp0wSwJo1CiBRw1Ynl9Bh0qfnHDekPfPZwVs9lTqNEPJ/cig
8bArzM5O3jOqupqliu8dfdxxGcmztxb/zAKF5SZzPR3LLKIdvv5OwpdqDRqUOpWz
McMn/nUJVTPGx2l2VTZU7pa8qaOgL2eced2UEBt55Gu72MRteajx7vXV0oHQzxTl
MMicuP3zutWEd7gnqpDZ0hWGEw7LtTcrK0/EDFMpUceg1J61VQntYENvluUGDLL8
QzVVGjhHmaU5rZz2mE+/P44lbDbcy6jQN07Ro0M3GaaqoENIeM2tFFPi8kkE4Q/s
DjHqK+5zAhfPhGJMhc9JEMMRJxiUOMqbuD2o+9XxQnaxOVqgUQoTQbXygUvVSgzV
maE0TSQHeYHzs7JhdLOMDS+g7kuc6fBc0q8oNrmqALOCi3etR9Nfljd/ChP4L8cu
59hKlScBErLdmIhjtqwE4ycofIMr0p0SvioLKyAhzRUaffu7PAjTDf/lzTmu1Qtx
BsF/7JYbTesZSQouXEkQECv5aALmG9lZ71I1IxiBIpbHGyeBk0FGYvSBTXBg9kLd
IFnZviF/J7JmKYxDcWt1lF1xbQ4pchdYwMPO/IyDbTotcUSwabyepcvfAc81lAkX
IOk1w9r8FTkxTOCOIftovO8FnUeqJQMYekM+1yy1nFMGmDn5+uLfppwMKrJEKHMt
V5AD8aWmUxOzDVGiT1D8vncVIus3bZ2FJhv/nhwBFFz12aTzlT6TjpGr+em/sDiJ
Bd1PKoKlseDGhjhLu6863gLAHCTBlMz0HEn70zBmrRCMMRGwFrTKn6j8bXSA8/Kl
O+zFcGKtvQJT9vWgG9iQW1GuGE39gOWX3iTVsaNbB5+1YlSVqx+xKF/Jf14bHhD4
PtH/PFtQWZk13+0vQHq2fSrG17zVa+j66VVHjZ4AUWR5wk54qjx1y54hAXgS6QBj
J9Ve75ztmZSxfJ5gwBERDW4/dSC/xbntm+a9UgPTnZT/igk+jNUy5+5BkpO/lHRV
u08btL5DAP9EHXy9djlduYtMzvY0ieSq9YaG4qbP+PYYuFZ3wgHkmxwU25K54XDv
iS0pzRcIpAkkLyDHuYSNKptdLa+CdUSWt6+GLVaAuOdWlpV7ZU97RpshknF3d0bd
WsNLhvrFD1QLi5PmM2q8uNnoR9zgVKT7CzqO7CDE0++jwN7qFEpDVUzWGAYn5aq/
i3f2QciKkc8IPXdBfK6hLPUE++WNdQo6JW3PpnB7DbbFTDyEvDAMkABQL51Dbg/B
1h6hNIpNEVBSiowsZ5/v/l7lLCaumssGLU4sonXjfszy2NWgkAeL1PC+rff0oe/7
pbLDcNT+t+S2VnJBpbWGgrKnpyIoqAGTOvUsZpBOCMvCAIAAX3h6AmQo7Z1l0ag7
QBWeqJhDudTOlZlZ2o/CZwIZe791iW/cxXx0MkdNlWq6zdfdeeLK2vfuIyv67m8J
MlAvjuNbYIqImTOZgEc9BLvFNVlt35etyUyRIdV3t1/HUw2y9eMBJnE7jHQG6R0E
QEzFV+pUMusZ76tSQAsnp2VEam0/fZYxSbpXgAYLgDeBl5+c1pEko7fiZfMZwMpq
hlVh9MkHpCScn2wmOOsIhbfwZhitb7mLkzOt0HrTJpNJDNtG3QjdVhBAvc/EB3lq
uhAvqZTQhmGyAYqGndWz3rMF4bwrs+YKQq4w+DmXUX64isZXmGl/BjyuOzld0wqW
04NriIdojEreSz9IFYFOGytV+ZqVycckg4SUMAUI2B2oI3/OugV0Tx23Irf+A+wM
MWqKibHjjNmhstPQQve1RJlck0z3mgtaSOMgZ7svNCh0SujJdXvMf89aeLmqz+EX
gVP0rTj41rqqVltw1/MoD+JYHBv9MC57J9fnlVVL/ycCsepIlB0Vujuj4CoN3zT+
gE9i7BDmAuKVDs/9N6hO9+trhKUfhem1MGfuApeDwgJHaWrrUldhRElZBQI1wNeI
9jiitlIB4BnF1Dc/HbxscRa7SSWr6ArShs2lSxRnymWMr3+W7xZ8REWZ0ZRradu3
odcW3McOuw62GjwtRy/XJLgmcfz3L9fm6ZVZ+Foek+Wdp4MfqlfzTkTho+rJaSHW
6tnnyJeI2Ag7EeByjTVCUJkWQ1sER6kkSxMRLrKXljkYP0HW/rXE94HLmjSmXbT+
otUQTu5HNqB8iJ/N2/lA9w3yeP4afjghIngvjL8HpOoLhFvL3aaa6K4KsUnZpIJ6
EeoeHkuZSb0hwVarUcnY7/vr+h2VWly7vhljWFNJmxUZYHpv1gV/fjbxi4CIRpz6
evvzArduwVWTY5XnwLCR+A+vTjs1JDV/EPomtv0EulO6LiUaY2d4SKqMBb5uNDE4
uVgnEXa1HKwJip7g0RXVWfJzYRLfNf6iLxBBOr2rEGbzwDWTKlhXy1dN0ae/eXq2
zapxTnB6derZjwA45YRc3W91AUSEfSVkOYikaQJkDUMDC3+9itZXBDWaukbHbVgj
j3N/v+XXlxHbRJG1g1cUFmZxCn/y4sxPElsxbSS85lQ14z3ZsqeHj+Skp5XKCHpU
9O8jp6H51E+XFUknagQPaBzF4ASKL+mMPnJ83MOOagsK/10bKe6feQiuhvGAUzYY
hpXild65B80Wfi6cjtnYyArs/zx/Vsc7fVzxUx/zE5WWSHM4tmHufNlEqucUus5K
Zz16c+lNm6hly1/xLsUIYnrw9bJHkoaxplazxlNl/nEfc4iObO0gU+wYDojFQUif
JpBEy3r/1qeRzBM9mDLYF46fwVfH5dO1Ze9Ry6LTWQ/mz6R/psC+AUslbEK9OYKx
4tsavyVh+6hAmI3De3mbyhHKrLaLqxvXChW3s8ZS7hGQE2VcKog7UEFMdmtrgTmz
qZhDOfCMw6ckfzZAa/SAiPhDi7eC8Ht6XsH9HekfbknVoSX9Osk/6sO0pdiUhzSo
8Le8niCvmKr6G/x6BKTjsObF1dkspDgA1Lpbc/a9UEwAHpBmqVXpXAGPpVM04f8p
xYyYZnkHx8EyKqPLrfI770v3+6D3Z/n9jYQTCy/ymGkZ/4assnI5XehTit9kDt0z
JTkQX+2lXitQmnpLPEl73ltyHzWOltLbC3PkRoEZHGFdIl16vcj4rUUI5PCOHCgI
0f46AtFY/7Y3qXBCxs+1ombGF7pv3gXGW0toH55dpVqPB/GUwA3/BYzlpHoMiUYT
xa5yQql19Cq6mtWY4XWwlzJCB0/YbyXr7dlzV7xh/f4+r+DmB2YLuS3r1iiecGVj
bqL/C0ATtl8L7hPjXRgNBxEIDGL1+cIdlrzJVEOdHNxhEzXih8Dyj6TkOBWHlCC1
8CpkDItRXyTK4Ug4az069WjRCoHziyWtgwZ33+PLwkeUaJ9RmCiCZKPwMKqJGO0R
YomtKqD2cOO+mTdw/L7XWlouRMOhNAocCT5nrRb/D+uTyYQ9kCvSvghNLcoYGroI
Hh96uIXO2Yg2mgN0DA92BaDuHtGV2XF/Re2NlAuJIqGioI/nptM9DviFkoAjUMrP
4+LATIZXetdBZpOjlTtslPqOwldaFceWpw4HLfwS9fHwLjV6UEpNXDlnTHqorYRr
4IVVKzCs8bz3QK2y/EW9zsclOb9kxcxkLvY7avBAKKFzyDZUTtEmo5GM43jBiAFH
BrfI4q7xN79nCaNC6nmowVjqksi49WMllClFY+Az3/oXRKdyaJE9AcnjtKPWvZcA
5Y87Dlg9mz9lQ8oMJAB7rOHDj5TSxCoqXTgJtIP6v+e+Pdq59FRMwYWkAmbVxRQC
X3GjEopBEUlXl36d4PSxOY7/1qXlszMATDJERXyvVUDLhdb/IwnucG79pvZhZEZc
QDgZT63BDYsTcVPgca2fluLWv+Lhitj9Bp/fMiWoNRahj1CN0727HjUs3uwT7YfA
jbctluAfpwmiVu5H6yKk9WduWg7xNmGrkh3UgV4q8GuzDVz4Lr0WNiVKYBSMqbmX
Hst3HoqqMqDeMba2s2cSATbRrNQ+525pF7N4jue4bVgvohjywGtJC8tREGM/NT1H
8SJgnK4/p1A8NQYu/Cq3K2pUzDM0HLqIAbA4qSJ/f1PoB7Jv42VAmY5VFdQtDE1y
+yY7eV8P+YOjKVBEyJqiwC1qIFkj2wn1gF4fqlUNbGm2B+qFCCuTgoQzC37SXCWS
jwEY6DVAVacGDLzJQEcUqr2ce13vfB8DDTAjmzrv3Od1b9X5/S98BfXaO3i/fOyI
RVKbt/yg58DpXAj/KOzUUyDviLkz8Ksc6eMR48T4AWW+fOJJqJGNM2UVSNG+fZQu
U8kNogWwO4zXZqoATwR451jK8X71/pdfh3+3WH44s1CrWAtVddb8uIYfxitx2IAp
xOPMRuAlr9EvG8do4Q8YjrOxsIkIRj35k1qD/5vqgeLXazzKiLWUhiCG6djuU0ge
baANxt8UTf/x8d8EeYKATaZKRUMonb/yuff+jcb44uTmDCL9srw2xMV2jpCD/wg6
Z3aFPzXFADXQxTztiLoeIxWHACe4DAQtWUc7SdShaZ6lOHBZwn338vbsr3iw+FHK
Spoyq1O6fUFeljUbQYmIg9hmVg7A6J4VJ81o6ECo+JaadXxJ/KSgOmlDxZawUT6c
wqVrO3JLFBJD8b2a9zC7TPgDPkaN9IFui+BOsJMErlN4D00qWztttZAmvvCD/pwH
jsU14kXMRl66rqC4BW3S3caASFA3m+2wI6QreMxZkRDoQe0S0281JG/MVmQsKByl
Dmqq+Yi9FElML8xhtXkYR3FkBm8SbMmtiFGsvvQZo5s2ZmDwfkIr+gB5En7N7kMg
glcL5eUkjH2d9nEmWGh7+4CYN9eo+uQ+tbj2O2zRvuxFkBlfdaG3AyVWKjDRUs+c
0DUuMYvGgxSlsQwK/W7VAqBxm36RS9uRZ7Z4S4xK2bvxMEYAk1bJV4P4c08Wv5X+
hEY09dZsINNU7eFOFyq1QeNs5pGKn+FU59NkYVfQOXhclmDC+FRkxdj7eE96PVqq
uIpVqMfX1Avs3/eKeFz0L5g/Wp6YcfcxkX4ldNthnPA1MyLZPfj5HRcd2+lMyBd2
+aXVXCgU8XWPmlbwbQbfds47Npf/nR9F+DFa36651Xb3PNwc6tdnIK5/MR2Tr9YE
0Wmxh6X8h4KuGYCGZ9g88qayDqr+NOG5NDFuMr43qYzbEIKICHn/OshwZSeOw0Re
+xfgUlpbWxzOoDuv7rrXyHuFRndqLD8mn59lB1m+J2cjcHo4hMYUEa2r7Rbsmdg7
nft1Sin/RhwXlfVUYJWk5gaHTC55Zss+TG4XTIAMoFCRLbuAUOg0z69pq9tN0wJb
I3DZJ7KCAxahdsjyEI6wFv6uNzBKD4vVMkQVzQdn1UaUBL0TXDUtgTFFIN6S1rdl
ZT75AfRm6rVWxgq7WN+tvUq55Dj+jDpaWDNW4UA/hDvhMWsVLsyEqH3U5jS35ROg
x9WGf3RwG3c3T1mugq3ZL6r6vvImDTtZB/Y4BUrYK0tsKMrh7N3HN4M7hl17ha0r
Kk7xR4AlWgNiH6y7dPbhuHvuEhYtWrLBG4dw3oj5oVMGubqYyIwyPTUva6xHZfYb
/8xKZ7Ap3yomn/1bscPG631v4KlqOlH1Uh+h59OC2yo1MVp+txx7pGj99Q8wbYfA
BQIMy8qAIqBU3XIIH9TnB9DLqBn6X8GDhawVhgqkasNo2eILSZEJfYUmWTVkFeSw
dTzX7DRPL6AW8xYlfjq9ude7Q6cqXvKupCY21AD05zuyVFjM9r12xPY29Icn7Rt2
fveQ7jVhlkqciOB3ZLpTfNHVjFGJpTi6lgdae5A1JQL75DJsK/zpNKZNWrztX/3J
Ce1ZJB0/sILlwjVa5R8E2aq9/oXpTMWvvFE1swywD1b5V2jtVwteGwx7NTzhxgI1
cSAuPMcU2fZ1Ku+6O894BV98XaKRa21DM/V2YONedBM3Jk3sBs5u1jj3nIo4hM5+
Sd0kgmMPH6vZh021xRDLewcxM0nAQSA93+BDAkR7CF/n/QXlnQL5RJFBEiCbo8Ew
l7wdL5h7h7QVwaWm1DydWnd70uejQx5wRolrofEgkmMSOw1N2LFXdPFv2SVyhOmr
pj5yaiNs5HBNtW1XiEH06BX9qnp8YqiGSlvmIxd6SsPj0f6eGVty3fDFC5oErGgG
xvMiEMr9cGstsLoSCcgK9xeC+0cx0cEt7JvdSwJmXN05SRmBrie3eJC294V+dIw7
zctbE3jx9wj3db8+YDa5aW8MqpvrjNVELPCOdE+JZIZND8D2W7L7ojAvfXUvck5M
cSZBJKUk1R6ygK/Z4qWlkaoY/LATuVotxuA5uradRgjvQ0XyqXgZhMbFV/dwuuri
LL5kf7/IRCknVOWNLryC7xs+p3GegQKtnjQDBpZ8gyaR5t1KEPERDUQyj8WqHS7R
HkNlOulAqCvO0u+9WzjocKlA6dacUvC2mRwowdmoEV9V/Z9SiB2xsDRUYC/QiNFR
+8cS7bHs6z/FZyVeoxL6Hk/MLWUhceLuEavpkXNWLzGnEuKKuEb1MpuZzBgODisH
ytJJoRRgab4uj/yUNR9Fzr58nPgKRHyVOyzEGDrpvoxFgzOvudu1phgzTpkfddqa
Dp58Vrj1Flqhg5vwBc6GxpnWv8OcanbpeT5vfNSnhl2Qg4xZuCUaGtRxVuHdvLpQ
hjfB49tkBRiJLkzk9xOzASdBhpxM+OrTT+rwD8MmXYrG1wql5X6v393oUB1gbAQb
IFCAhvkf+hFl6E6BRiTn9fGUnzkHfiicY5nk7110b+zaa7M6qDDMYW7QYT9m4vsp
naayRJy8/hfPnsuQmzjUjX6+8pPBXcJ68VaIUWngAU4Cwje78JnSBzFa70/MFDTU
ctjMV6DSa/vusH2wxrjQzpiXVt2ftuvGONEGOAz88PtEhCmn/Wa/mE1baWQJqjXI
iR/C1M+U34oy1muk/EsUNZOOD/pH0D6+T8rWM61txRMi2aRaZjRHAD9M0oIN7GaK
neDMO4+GRZIdD1ELSorxQ0MyBJWOxWjOwAEFBzKFPeVCcZDmENAMpRSnJ21aoq8n
UJQ4mdUa2t/690BCTPDw1m+8VLArv0LL3gv2qIedo776IdxON7ey37Ai/uq6Pg+S
/NwY25ihx5/VifNz1oQeAtmjDZ2l6e4+krVQ8fBYC7R/lCSA9Edt4Y18N4LEd+0A
QmVznCdetFsIMX/tBe+e93m7OggC3KHpDbK3/HQSh58I1xwUQW+xRyMGAnbW6wVT
+6i6H2i6i0XtI/+i9VuIKFRMqF/kMM1MbE6kr9TnsyPQWNelzIRuiGJPLo269nLn
vTUku47Pub+U5hP5KQq9OMcdMXK0GUxXtgdlsVOzjySVl1KaEoX0rKhhF7M3dvTg
4FgyDTwylCYyd0tz2cGwuZ5JiSkY4asz88w8gVh+iz7zmeZ17a7fmZxJcjsJwsRn
6jEf8J5pDcxeR4yaoAvgTcWEDgSrypDAT3Z/gPqB64XRXMrnXrf2IRIbHF+cKuqy
T017TiXJwavboILgVitDQQ4nTwc4HC1wpDpUppliCTFeer+NHmd4zza0Tm4xaZWg
dbda5KWMjUJjzM+IR90E3EEJnM0RsGUrs9QBmv8J13uD6wJvR5c6K2wpa+HmaY8O
/1c2ZAWrIhTvvxKcOvT4017t4ImTQbKq6mcb9gPIHqHnbVI57b6JUE9b6CM/1QBs
3ueb+Q2zmAM6AE6Io+PKCl0+k/04Sk9FJ3SZ2MS1XYwsRT98nVVFMTRxeN6KWNGu
LA73gWQoyfXFuj+XAH78d8lnj3SL5LH2qdomhJdZmSrwIe6s/zC0M8H2HRpP3CNn
RUFTZoQPLRnmS4LrHMiyAVxjepzODf7TUbp3PwE5+GxAh+sR1RP+0x6lZs8AvqQt
N2dEbaRKtErdixN0Cfw/Q1hyDNkRAMev9jfraq8/Blpf78+I3JQlgjQTUBsentsD
ZKk4GohIP8TyXIB59yaCbhA3yWRuOOIXC67rO8MHP++IZIv07r28m0R5H98b2BSd
NZ6q6/tuVatpm3KlYZRewLQ4TVOne5fU/JwDdECgLT+l4NW1Kg0KeAxBW2Xh9sUg
7G1D2IGw01SwvdK8niTIMAxEJe16spPOJVuLDMyYr3u8DBTGGP/+uocb8ck8XxZI
XZrrkiY3qMJsgm3dzNgA/+3s+ZPoLnhVSiOb9OVJejFvyjpLGuXpry3amlMNX20H
Oo7CggA5OwdwLZRPyGKeFkvS9aaP5gv7aMtV+8UiwB7PIkOkBGy8QtYrv1Hikyi7
gSF/OMLrWIF8im04t2hKyeRk7bEPdbZki1686Kt0NDveNVXPIIrEpLvf5dC/fNTK
h7cs1ReECEXiQCoJkO9YIwD7u3ME8Dulvl3tYMk+uhkU0FOQvzoPWEMq/ldvCKjQ
aTaDWCeHEcj0Z5nIyQgb7oHvfRmmboHJsx21JojFacrqpbdVdQPdag2iBZHl8Ytr
fXAdZEUdwCUVczf6ea5lQEnl+hCV2dJS+b/lbYzTScDSj0xo2LwSYDw6SfItnfBb
t4FJiTPjoxzEy9blaFusmCDS7DtAQ/goZcoHkDmlLvuX8w8kLGxrkFFF8H9PFDi1
/CPmL9OirmH6XWx4FokahGOjTbXcoaQXqHklwDcV4Y/OZbC/m6m45ynMmy7OoaEO
xPCGtsrKzDba/mI97o+yY8uRtX5YTDRmVp7O6+Zs2jRExWO+6IS3MAlVa68dw/MU
za9O1sUCgyZiePECqwdPhTjCfWlLR9Z2/CEUxikT4ecNQqjP/hJHloiEw332L9La
dwyD0Un6JcHDsFiGiytfSQvvXvB+eDmjDKxN/OGVbxl65epn2fLHvbug4MGaNLCX
FB8c2zhFj8C2Bq7XC7uo80wVwChBaxuYi2fNFxkp1QeqJ6h7v+UyLmk3P0SwOknD
hVV46W05qkFqvjNNC7jihTiEihth+fYTbot0zBiHFB3p2WNTbKZv0JqcwxgkgKCc
2Ty9C5OTYX5c8+j5is98pfBh9xg7vPKVYJTsdXJR8DSxwbxxMRDFXasBXtVi79fI
OFca9QhSF97MCZWgYbWnhWKOShHZSieNcHyudmn+AZ036c8VeCHaozINXY+cQBj3
naWhxijLJ4tdHfKZbVQwY3fAJ4YtokNv3+xIPtlvmnY4xXTPdcTi2CAeGuaFn1Ss
pB8RvId0zXMr7QQSJkt7jYYf4hANo6cKNX+yZtw9zArpNbD34eF7v+84eOzr2m/H
ZekXDliHYU+nLPmh8fW6rIaEjrxqNn6N8K7Kyc+6V8OsASDOR2Ae3AunD3+kVNsd
ffRWIRrB8Y0/Gcp///mtcuUeCaeqxkTWvjwiCbdxJfNwRDS7a4JxbwmxGS/OhTJO
t3rNrdFTZudxiK40CK1B67kmKboiCl59xEbx7CXGLVdE2DQdKcDsPJO/sZhfu4Iz
RcP0yLYxFAhOAZh2fGA+nvv2YuhjwNMddx/05Dbza+cLQI9d8AQHdrriaunSXA0R
MlYJ0VPvkPZTmdRJt0rTVji3/htg5CLVEgAxXJFQDCQhtpd8rwn5zOeX+408GH6C
nV7Dq15BEevLnYGcaJDe6/MD5d4yRDmdviB8dgDhz+l/TU0D3TfL1QZVszDoLlcv
QF5dyuCdJov0EmXreDgbRYCG5fWlcRg1Xpb8SX6TvsbzT83JaQu2zBAVQDH2J+1l
zIy7z1/inWpJ4vIZbyw8WA==
`pragma protect end_protected
