// Copyright (C) Altera Corporation. All rights reserved. 
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 12.0 windows32 Build 178 06/01/2012
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6c"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c/GFpcPHTT/OFm/cSFsDmqXro2f5xHiIqsF4UKYzKc6/kN8m6qQy5Tcc33tl0/+a
QvbhE4LgU9GAc0Y2dNgrpSihTXUD172i19pxQuzQXU4R4CSTCIu61ozEH/OlsuZX
L6dga1J5PYjEry3HxvmVkZ1S/oz/Se8DXGU6giny/6g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 128528)
Vzw3txZYXroSfhfNym2hVB/y+rQO2o3IJ2bP9AWQEfbR7RgWhrKMFmKLfo6OJm1c
aNTiz5Huq+1Gfx1xIsc7CuoZICUJf/9SifMVYhf7p5WopwN7XOF/tdxyHCJsbPik
wGy5FlijZ5kTKQphZ42rZvSTmiTrU/H6rWwdiaOjyatriyBdpJznr639rWB6FvSH
bGhDU0mpa35CW0v/WaSVUT89WMfAQ1g37/DD4sj9OrCIm6+39Jr/0wmBOBTDltuc
Y1kgUoY9SyETjJ4pRPKStQxQc7hl+cTo/ubVrfxURdQr75Ro6S7+iPmUzC4s6rYK
JIjkIwYZ9DP8rlY/FOT05o98q38YMCaMasL2qMmhN8kGPtEaWrm23FuHd9c5JuhB
VtwE/kfD2+Csa7eodfgzChqN8z+n2mFF0SUKcS/f6ezTjBzq3HScfrJWyCxIUr8r
p9BvZNHdgETEqHZh6XMNgAd4dYTNW2gWpP2AkH5yi2OGCye2eeik4xYn3AWVc0ad
ubKQKCbWz9jG+J5THCYfYLXOqX01+LpGnm3q0JlZ0iYZwIVqH+1ThLo2LBEJkICw
6djlZBbcyR1RKKL5zUc9pjT1WbVtGhDSa51ZWt02qouxyNEbzsUiNIfb6bU3PHOP
+zC6QeunnlLQkjUp1JAS29wVmha2Xbhx5IuXP2/xeyHlVXJfhgO+i1EeX4pK/Gyr
7un+V98LLze4HlrIDdm6TeIJfD65zHmmf62/ZVsjdwcVSWSm6i010mE55VIfBUk2
QIyW3eYD58Qbtld2GGohorDoawb/pdwax5xNG1YkCy/FAHG5lqnPH7DsfffoZOXB
omt4PQhfNsXHgAbKrSwZ7BN8rAMi1DllPsRpRIUmN4cm6lq6B9vyv/IFoYVTjuCB
Ib6g6H0MX8ZIjt3IJNF9YZrv0prAKzkc2OC1tlLdoRC4lFUVxQ+GtT17W/Mqb6oR
25W7ibG40GM1AsAe18BKYc38uSpsilDLkmqx4xigu0IJWiAnWYpGpEeXhyAvGwoA
qDDUpZPI4LSeUTPLa8Oj3cdqYPxxkjcKM/l8PBicU7WOO1F5YtIeRrO4ANsx9GcA
io6ggfREegP/bx/HWdsZXH17eprmclCU4xv9zxdZ+qIuXyijmzNlMFlJFzNZXD4g
2CBH1Z2kmpG3ikIgfOxkSUVksKNtKsxjuR1YA4Hg+0JTipyS2xnhHlOe7KzkJ71N
yiP43TdDSC6QDKAt4jO6cPWXRG4c7ppLpmoAZ4bQl0uyT+bvCmk1mGRCcPlX+ReV
fMTuR7jJDiEP5jBj+kE/7ICcJAqJHhiRtK1QWvJaVvfNJzLGFglX5pCFsSdkJeSq
QgspGI+WXJ7kpC1L/Bso8H0GOWy+dZwk9gM1ykUgFr92u6AxgLa1LQcpkqYdzuSq
Ee/RWFq3JYw+0dPU2JcB4oxMLOF1Lr2qbtU9fa+ORaDkMcuXjAsYTyRUt0FSeBj7
V/ZzdakDX/zfP24EFs2jDQ3kZJWYChT9tbDp1zERn0qE+ySUuLpaYsisg4thcXaR
NBkqqfHgCkNUyUGYIatnjekvF2z4MRo0jhcFVXoFwGuDy0laIUzV0IG80Hbfrx0w
JmSumdXxZ2zJqoRRAK7xLexl78e6geIIpGbbwVs+Ymlw3D0rmFOO+zFStHTAWY+I
hvig2rm2e25g3NFMThnwHMGXllwQtd2IpOF7Y/IUENQPsbdyDFicmErGfe1eQ0bY
zijOG97SQxA3VDzOP2iDelYwU1j5a3XhvnLjbcbOP9isByiFw7K2plSjx0mM058+
4n12L2bUyWSibu9noouNZMRPBO6tnEu+O7w6C0k2xx7CM2oFilqEOflw7yUnbXFs
ffacgBMUapKg0tJGJLeQbmH+gO5Rsok5QIC4BY83Rj9WyHx1xF2nyVaK+0QCNJbv
0Dwl/LKB2JXiXhuY6I54gX4VliRjd5SF5Tp0ur542whT4aI69MdNM5kJnhmPHCZQ
iZXaG9dmRaIKZLmKwZgftPwz757eo5VpJ09i/8iS8tR6K57UOJhdNTz2ReECJ+CJ
6ZF8eolZ6xcvXEJOIxTOisA6yTEGqmMbb6HZ4IG0AuUYy5eMP9NcUu09TSPSThio
9q9wgDISNuSyQRPhf3OxKPOEfc5/s2oTlE4U4YD+hDLsqW8UOvcj9BlFwfXkj4jw
uRWShseaQg/Xu0GHAOAKpx/svWGJax859AgcxCgJiUfSyMjAn+yVxqagValPgl1E
lKzZnhB1s6hjTAzOxdDjILilxp2MO2Xy218QR0MUMnN++arwjGpN7scLsl/149GO
+QgwKYGZuk9V1CXiciy97tl27ah3hMo+guOs9WGzItAmr2wP+ipQz5+Ekx/a6QDq
HNohur+qIzVlzRMx3m9H7dWu1Xj5izCpfG5P4CtkVl1s+G7959wJmLwVL6r4aOya
v4sE8iLfXFFDv7EPaNfmNKT57ga62REQlw6aV4me+XR8x5FxZZ1d9XsxPgspHYk5
hChotkudZDWdA4qn1MelTWAqUaoxzcOgF2mdrIno5Bzb7qRI2hNMMwwgmqgiktIX
Ue0k6uPcGanHu7gLY7OpZ5w6Xg4Uy6cXI0s/DSBzEGUQIBcIQ0MdSQ2jwS68RIhZ
w41A/grYnjfY17ESsHC6q5s2QTxUNOzNjpiqjVWsmGcoG780UiBoufndOzLno7hV
/bPzFiBAQASjJW5w5dXLG7Ko7qJc1w96Cm6igTjKKjUKVAWHJcsoBNwXt0E33ovp
zXlAPXjKNTnipRPVNPzXEQVRxxY4WBgVKXSZWZmXw2CNFpowBybvrrLpFYqKQ0fB
+vQjdw0pEls8X2dPswZR25lUxiv8qAKmRLH+RK7/oRfZfq03Pk39z+eO1CXWsnEt
aOmq4ZZcp8cd8qM+BBdq9H2WQqKFxbiIMp+qgi76FNFFcVQ6UXbckZ0m6Z9XKgeT
lFPcrRnobGxaxk5o6RhELgc2C+cHZusC5r5Pq2o+BH0dkSMwby/PuMrZcYJ63GB2
8xZFbrIeuTYpvEhL8nXNL+oh/fOIbLeaYcXbIyfhPK7ha7z2xPqoM3sVhrwCiuzj
jv8GTTXAfGmHnJLohvD/SFWd8P1mbj0+RKp9a2JPCy/mdYuyeahVjhQewKB3xJZ7
LVGZvkGFYYPESfqr9TS8y1m38jQ0GJDQ9uOkVdbp0fjepZ3VnyuuznxUkq7F2tGL
0AvI3JIAb1QAmYf+B7fP3JOKTJhLf2lZipfBVowMNv9ql/sfsCxVa5MrAdt+fgq6
DysPUoHQR2R5u1VhF3+ZLXbS4rCrZ1wcgC/DzeZDwXWmmo+hhzPmOWjFzwSwrOB9
oQOIdJAMuHlQwgbcms6gMk//64X2Xac/nGaWqumoOHEe6UVMKtnKR5MahnHbjUZT
8AJdr+Wx4HnqW4wkoAAHlkXZ70xy52d3PTtrZ+E0SOJzuY/pK9HG/BvcwszhAfPr
Vk9XpCKAKeSlQc4g76Q6rDHC8EYMUbtQTqzIXprGSruXZcRgOZCvS99lqKO0D4dm
zpypvB8YvUil+QRbZVqTLtaBIlo6hC3lr08KlZNO9CyjNpKRaJx+x/CH8LrMyb+Q
bk4ueH4b7OmSkLh6K9o9tUpRNtzkLSERiqz3esTVqhhI2Ha3sJSkk1EjE+l9FKuU
a96OfWyJ4qdWVL0S2Onm/sCRcs23BIdtlgcu525nJwL0PE1X1LWeqm5PmPHzoAGR
aSTW2eA3Il56qecLGRIHKz51Fi3unSDJqifL4l7awmyNBaOU1JdCO6KwKyMmBq+H
44HK2BMpq54fbvfEuvthXCBTgerwIbbYbYHpFf+CUuoma9tpimvvLfvLxlaynlzf
1C+cAC/igJAbjo+YufZmLGIi2jpT8NJ6dFf5Qyw91Rf2tHAnk0QgHbd4F5kZnr+3
5fH4XaC+G/nh8MCgj8pJX2qM2W1zSQgfEBIWngDSrSsC2Gfqo39l5OM1xOTxCkXp
H45PKwWOBDH/4m73ZujyRs+o5NlyGajleNwXQD9ubg2WQ+5tv3deqv9u7PF9rB8t
Kd1zhtrKfjJwQiZFqWRSdP9UvJsk6TFxKfVkyH+cqwPdm12tWrJ7StUNsmO6keGR
0d+B3Nr27ODUVtkU0cYZOwYK+evTJy0lzPHoAbfiBn1EQnEHmKixzHyTl6e63q0B
tmlCTKwhxUL1pd55mHj3zAZ2X6/DtrrzO6ybjZLrXd9uG5oVMAEPleE4w0hgg2MJ
kjox7m0h/KUp3WhSIh6ivUBi1zBOh6+D1EBBaumz+WA9HOY3aqvOFVkzFK/V7HTU
iXxfiUaMZP3QGYuxhHMTRk/33Xb+HJUhJ8FZjadhKQAXzf+KOuF2QynxOVzTOcn8
lbaDLdXUj5KKdvhDjb+O9Aydtql5eR9egZ/tywo5zw+Ssfjebz6RXkgusjUTH75D
6tn4kxpOCgVLBAtsQg+gjOmduADH/JYNdZjzRUjJtO/16ceOrw/tPLJhmT8x6GHR
NN/T2uDmKYeBgUne/14NEb5qutD/P8xD3ILtOXaLEPmCTF7YS8bNzxpE+NYmynCP
8plGKZAvg8qe5hvpoH3cpYs8ndIzcTifSNLNyQCUDEKB1V2mx/wtNIFYkiYI6ULX
yYX2zHYqvEfYmPOLhit8KR6i6rAg4gweYwmyMfO5bLnw+gR9QNS9F8mAb0H0ltrY
eXUsAU5fXZA1ZrqmcuRQEv1RFDGPRvxQH8RGVVkG44V1vcpYEhgwr4Qp4W0JvRjW
cL1ooKssyk2G3IwovudAQinW0AV88YTcMR9sj3JeHcVcVOhOVDXg3N+XL0AfU1WF
ClJHQqOXBcsfW8sUC4p3iANWpbDMWQe9W/ClH7XFUtprNrvD1qNavW+u5mnr0Cm2
NnZ9Gl/CjO7beLgUnxag+OuW3jcaJbBHzKFxdQiToFfdWoBjs/Y+Tp9YfeSQ0xUx
igeAx0WBv8220LJrKl0DjEc2JHXfBFHSwedQ0XLnG85yNmSvoHbUryuwuNrh5yRC
WyzeBRDZwjrNgJ0pT20gwk8ec3wWmNSSl59SEOG3aapJj5NjV23pIQx6pnuBaQhg
6W0htMjkVtfrt+XF29LD8SY7GivzNwUhmBH6K70MpdVoTpEanfRWu3ht4piT0/xS
QOPstwXgkN4yrHwcKlrk0U/aUXpHDOqq69Af5o1s64+G6nFBt+EmnYwMQ63HXJ7q
PViZwX+Da2JLYqdXjroCGPwxqlvdaUJae5u5XLkyyuP/axwq6lQC8OSiccDNVMST
RrOH3X6PEvAoWilWVbJExufPf/0SNsA30JY5r10p4wdTKwo0hAOI8BjhbQrodaAm
pRbK942DO70U899J2/d0DbVxOzX8eL+/lSYiqO2awtxTOM8rPUb9xxwHlzoVpaSU
A4EFonAMF/wojhFU0uLwbuDSpdl7ukz85yt/GQ/ETZFn3Tf8HJBd3gAx7v+BEYVe
jgn6Hy3UtTKPp8NBViW6dmnY1cW/ENMdT7ahZIkHwIoCOJ5Ax4mIErx3CZcdcw3S
eMllBMHB2mlZXzaZ9nuTHocwtu9i/XYRrB830X1MAr0FB0DO8Pwg9iIQ6g/Rtbg0
bznV83u/b/EhYRlQUgFaHJI6+Gz9whilHOCretCHASP7KEeia6C2bXsU2qKjqA+g
4tlXQtbbNrDTzjZtYK3aqY9jtEAbpAzN9aj46uJ3/W969suWHs1rAgKEIMJaAuCl
b0sBEwxAVzgUctPW0MnQDbq9T9khSr5EvZL70JqGnpscGCyEtdytOL8ksdDW6i0V
6+dW2wNQtJuzipNZm4J1zMyopO5DYEhF5bvkNuoapJuSNLb+2xXNmMEBNMsv3EHH
LAU4kY78yyV7Qv6YroJc77LyxS8Zg8qZ+nHfZ2hvBkXjkvEIvSDLPieSDIqNHjg1
fd5SR1zBrWmcdIWjppiu2cKz+vUk0hMk563wZxdFgyYykousVfLlWSonALi28NzW
4Og6ve8hKR3NixgwzF0pfUN1mKpwXInZ3RRDHeXA9H/+IvQx+LRNv+JF/uPuEV3O
2ox1Ppnxo0yznY8RYzboxAUcmYtWdKZT577q86ChwPdnDmAmq8n2WGUuiH/v4JHN
YbphGcATU1W95dNXQ0Qn9Wk4jyD+XYmMfSuTAEOkiXf4UaSoIef549By01Liyzcx
6Rbltiq7NMEHfk2deZtGILtvzrVjepq6V5oyEzB+Rn1ZXghdP7gRxYt+mEmJOZht
mWdpsPZ2VHLPEf7D0PqgVCLCRQ40nc/moFjwOvBI10HUJWFeRwsgJFUMZVThbPts
jz3SG+A5Q12KniXIydCCB1lx8nFn5eyiFlNtOCI+ecUMGtxMKGUhfH6thoZqAJaW
EPASFpteOrtVTn9CXZUjZerpprau2tittIFada+E53TL8g3Q29EjPECO6HraCXX0
zSzmTlElgekfVs6L92O7Pe6og1FnbxYPW524ok4io/h+WMAMcoC1V0mfW9JCWJZF
TIEAwTechUjA/ZT8E8xG89FC36zbuyB3GsAm7oymlwQP+1d9yrcjNb5OFtb7mpP2
tvtQYh+bN4hvvt8aec6So0qnov+hESBd68pTS8gVYZc7hxWqWeRHxS6T8IS790l0
CxFRksoUw8ds7uTlCVeKYlfG+iM57JSKbkXc09OqLPD3/sXbhyVqduvl2Q9BfZ64
+meKWzzdzYi4BU+EUUD8cU1VSVIJ1ydhZmgwpBRi3AGv3AoKxFBQCCmVyHbomvlq
1EueIpqZGZ4tlkN7PLNs+d97cinpFxZ3gL+bFajm4OOF7/eY5wrh4520m76DiVoC
cmlNI5jC6urIw3KgxurMC3rA2gsnQHOkAOm0IsxL0ctp0pKCERFn0ke58wdxb1pJ
5SmZ+UD1+9/8HhlrrE2N9OHN2zaRbnl5u9NgJPdde0PyJ8FwdqXmvh0HAWV6vKmR
YYV35bLy5TEmTawVwfgoa/htBUNN0t0Jo4Xepay4L9IkhPTCy3XyWZUId386+NLF
3D4L+EOX7QjONq0S0VPdDjj+SMZ7Hg4nm5EC7kyAym6u9Ot/aMwLIE/8c1bJ7tMV
WYGEQU1qSDQwpzK4eQ/usgF7/yHa8Y3ZsY7F35CRiBemvJH2181lw5Lgrf29+lEA
zmlilqU1vVO1o/xLVB266z64X5th9bxAsjj81rd+zAuV6K+lYrmt+qRq1C/DIf2v
1KbfEu5SI3ALRq+0UcjQKfDc+RszYaVQy++xzuL9BArlZgCLh+cuQr04nT5oB5Mq
tk4cpMcueTPCFXPBdkhsMKsIDDihowJoTxbVk3x7oEP8zVnc0ThKM+1npom3ac9F
h3tELRkGgqL/rMOl6gjHDulJISFyb27F8OmLNsbpyQsglmqJbvjKt4AjkDt9dZRU
haQ4BjRYTW0JyMDXN809cWqsKjOPDsy6cCbiWdMPvVauo66ZRXLovfBGl+bm7Syi
aZkQaqP2/hGp4rqMXhbSbyOeeV+X7CfM15rQbQQbg8szY0mcvsM4mqr7jOH7V9BR
wHe4q5W38jnmBbAiSuZD/qfIsevcICEOTCcYq4CPan2Lrq2frVKDaNZdJn90sk26
kDVK8c7kJ07Oy5tRNQeUdu/0mt0I5fspWEXPfHHWxI8oWcgDYECxR1GcD3moWhpT
pmnipY7ZzatJJhi7faquq8mwIwTc+dhUWMDVoQjDqWGzAA60lYffElMFsWDrDryx
7GRMdTTDSCl/c6u21eA8LOqilHfNinBrdMuuXuDj/FLg7HFGwUpjWKbhqq0TCunM
JLAGRpPi6cFSm8wugZ7OfN9v60n3HGJy51NchN+VHLEjwvKbe/hxXbxMT/Js/Blp
r3endAgzd0DPM4IwzunI/0qvcfCoWZwwtD4+7eUuqU+JMFZtGGmi4UsGHKnsa/zI
OB6JwDYaSpcg8QsH0GJhzk0Yu245atvc5k+V8m5ggWhC0julMSvDYeJP/In6QC9w
RFvKyEGcaggyqx16rtVQCs3NFSncKihACmfcUEHJsqHPy4vGGM10t/Wli8176Y1b
qjae3E6DBLyEeyJ8+21aYb47Xr7kYGVOP1NNQ9xcqLr6EZFikz41GfvwDr00iJIc
ZmUAoVsgAxniEAK8plx4XLAnL15YMTMW4QJimcGH7vG3HTjvperrSMt8gdc6usCs
Xz9RnCAWx+WP9L4Ck9RHL6u9hdxLPcEX/5eXL9FttnHHbH64cm+TP84qKaEa1aMj
jdeGqNF9oGz2uQuR6kXVqbp7LPfHnp5YPIjZde9iHHlnj7fltxl5Dv5IMCjl9+ix
illzFG+ut/2RdgamWtdax37bVfsmf4x7sD2AMGg4xkyBSyej2Tr1YUh2e3LmWRr/
milcibA1ds4lMxV8nVVhGECAEbeAPA1PDuVhTzup4RCsOGgmnc43G5ej2Q5JCLjy
s57ZSjeXsfx418QiRbplxw+qFnliCtrLUDk1vEYQc/9uzYpkL8uU+5dnVHGtgZWw
kSJMeQjGQ8f/J5q5F8sbjWq8mYJO2ljhBKYClYAyIlHYil9gC9W91vcfU2kuMDbs
8QwI+9rpn46zdaqVVBhbxijq8NnTPovAtHnXX/mWHXz1pfrvu7QqUMB4/xyLcz/i
M7zEBMSsW1n0TFxa1yTXZ/KjLIGfBk3WB67fpb1R3KXecFUFh4pxxerGgslxzaG8
3iVABrrXECtwJN4LQ+QZD0t5evGv52nNu7V0nx0gV+3aNchSBT5zDUJB4biPQjrD
u0W3jN/+R3VrE6/+bqe4bWIU8VP9PPT+FtP4kO57HRhrUlpWpmBg0q0dlBC44CYk
72VU+OcM5Gz+TSewnhyqKHY76iCt9D2anAh7MHHfhwOYKmkt3G58W562n9lb/n4H
zUC5bJErVfHDBNy0Ha7nKU3IqSNo4SKca/jfCJRO5XlXlQRmNPMNlL5XjH4+U3ur
jdfhjhUFk/3Eo2g58y+Y/FD5X8GIR1fPEofgTMrUamukU3FeD2/7Pd9ItytvR22a
DT9gq3wGVy1H5WiLHpy4wRHM1E0597tnyIuNOuWBu+73N2CkYKSUAW+1+2MBwRZ5
HTK02oHhe5zjF6lSE/7YMToWgHb3TSWrRnbJ8vSDC4bkRmCmDqIJoqjuG9GutRPp
wqylTVwDhvBpbMC3z9iywQD88wUUUCpwGRxGkm6+DMRwS/bnhayts//f3Sk2xa6A
n9GmK1rKSI1BPQMV500w/bILhb4NH1N7gkr/hZfSikrCDIEmry0OFySv1b+YUopA
v7yqyRaX711BnBi2aFXzlApI6LQ0y3WvginPQrwKjSsR4VfppnNdV2kyBX6fovb6
ffKwGToK4hmbQfvGFYgwX39VGm/e7QNewuTBJBR4YdAVB1M/c/cd8ZtkVARFB3vt
xNomujHo2SwRk7aPePscEAVF4P9XcRTlJEnZAxuIvNj88/zq28M1YiDoPKTFBdix
H6wHJR9DgfKM5kVSMALmTAohc2T01wF6lT0VYTUWOlipDQFjyxIxrL31eAlq3ZXc
A403sGHkn4wtFXhGW2vCifmS8T3sCvR3RuUyW2+GnyM3ifT2GbqBmiPbzcgoVgr8
mtbbXudImpB0VDkAkCQYY7eHSXlLgppTUa8BbqE5xbRCc11HqQTqCesxichNBlQA
n+0HY/YLVA1L8aqFaCtdeMbnq6ibI+cFCtGT41o3hKAdzAOVoLlOMg/nPaaOKG0i
A2DtjqBW3TT7jl7PUFsxuPjRsciK7lRs3ZY3bS6fw9qKfuCrqeqFgtmQJaSkpfFg
2Ao4lltAaKIxKV3dEgKcH0xfAduMIk5vkzG7d4d1oKL+gQVhq2DX5J6HeHBdCZi3
nvnZAl/7TrWTVhm0YBVERgTc9cBkDsSByu9BkyVlH7yeuUEXT6Ir1P6s+2ylMr1n
82T+BJy+vrIgHU5PJHaE6DG1YUvTe22NdvybkM9z16q/YhvBm2qdE+VVv6BbQxSd
wnGBoTFNcs+HAz/medihKEkZWtUYKjcQAI7pqJUlHxO6Fz3qgCkgZqJB8bd6F2v6
dDc9xxHwpDd4to0cVIAao9JXyV19oQQLaGkV2Y2S0WXRp097YZcGSziYAPLUENjz
PjbSzIgjuxjf7VqbeZTRkicogiKxcuOeCHSXJ4Ey4gyNd7A5AJhVEpLeCE/yCCMW
Bh8J9RMwQOh2JZD4Xfe7Eq3yTDsiNJJTpaDaUq2NTG0sqmAZu67O+Gkaw4Y1dnC3
i/0sqI3+6whA4f2KcAKBW/xBKFgIaksZfpLZP5IHq5Eqr0CW4OxGRa6+81xxIDQm
crrCzo2ILrH4YIcyh6EESCvsyVFH9A0BzjgI+oMIQaGVz2rhWjGVlYU2wRICTdw2
i0ErlQQtrhmIz8P4E/ndAH1xJrohk0DZu1BeqsAqJvRqVNwghovR/CZoRIH9lFw1
jiCuP7Fnk+JR6TYUYInUsOPmvbvA/jjo4/6GSRRkJ+FCzmaW2uQ+xDbfVdceyltY
Q+E+i7D+gM9LX9ii4M6ANPS9hDSWzzklPyJG1UB3WvPhVOLwQd6/clkIb1m4+XpA
7oGqt/FHvgQWvj/EV+xy3LUtnuHcUlCPgBEya+Is71VBHdJqV2lcgSjlXZYA0E5p
Gu9gjpAKucJDVOsMHZ3wG8p8YQzywoBijROEy416ZdmOg8JCiCGTIaUO1TsNLDPP
bc3fXo3iSfLzOzkA+mIPuA1EK07W0pOFQtgP5kdK37fmIkSZ+ew7OmCvqie557HD
CLYHfAlMeWFxKye2qhpv9H+8s0zN2vBy7qVf3PaUec469KRmJaSdcoKZO39mgD3/
uqMR634X2buedJ4xfpag1NJIa7XWX99w92nR3VSh4J+SwmjMpDn8m0JfcNnq8Qhy
2Ir/FA+kBrWu5mxdFsOvi+G75FX6Hgd0iCQLCC2yQWIg4yWmELrbAF6GJ/c3as9h
SiId7LAIj5x5tc4IXh66Y8dWVjWoOvf+bD6Abp7qG4MgLQfRwUW4uK7/R3AxhG4J
1cV0AC3vdH7uDR6yNUDXt+3r+V1nNpKdpnT+lZhRCczGnDacFPE2m7yRF+wntNDO
axiILURHDWOpCV5M+SbounsqrPfpGmGVyhEHirX5V++0XDytFsB8ngf/HlWW1Tc8
I6fmwNr7UfvE/S0lipndLBNC75vq7OX49ByH4UQa2AheD67EQ9V7SgXi4z4qCvcC
iM042HACUjV6IYfrXK10cLzotIeiqAPfm0BTZ6KfiTKdhBRfnLvM9WxmroFT/Elx
BdO/d8MwlRzCkU6cJbUwB7AbrQxNVjLI7iMHxxiyZd3Wb1ivwBlzfpmXtCQKrzeb
yO5FpN4tlanOmxEqHFeaxlL8WlykB1WfyI7ppISty4vIrJLN1ABamTYhJS7RTKRw
VZeWNS1kbUK6xzPac3ij+7eVaP9n13rf2rXizT6FzvpG3/9g0HwAFbiCt175+1ec
LLDy0xpmVRA568L4qAehhNY7Kl8YuQfMZLL1J+q2Z3lV7mLZoQpmr4CAuXeDHbag
NbdrzvUnFxA/FITUePJwRwnVva2DNQRXr1RRyp0Mb1dD6qAOla+qujOAv0Jr5tLg
zfc9ELfGJVG+58Eeib+3fWYPaKZa12ZUmzQ4mvWX0rMcJr2GkyBf3D7r16eTHIH2
pxWnAND1WJYIyGxuT8jMXj+sSgsEFcpyb8LBXKPn31F0CvLsJE9VuFk8Xwj7f6I6
b9US1jD+z0rY88bp12teRXWdm+uuWZOFsVRo7tsg6doQch0L93ADuN0tew8+kjTa
ZAmPbCxqWogBDwcHFx3FLvPq8I/CnfsyYT5EEkAmE/a5YY/H4Zw6rDXkMGnq4s2C
T4KZz7/LVanpoqylU+a61Kx085HUE3oqL6QBU64/cxGaTL3yaz7n7XYnUs9IXGxZ
i2kI8CFPBb9mCFhPVnz46CKnUUpZNC5RxgZENDuuSZ98flhU9B0PcQRTVSJZRXAx
S8UUXI9e7z+rztAeC40mHr9WxhQXId2ic2BGMzNM9PL2JznihhpOv4Y3mKENYCyg
bLkK65foiV+PZZEL8EJn5WNi9E6cg6Adf64PYiQKPmSekoG4eF9NMu5Zk0GxdnES
jMkyGp9XSEBrZCYVshG0UBXj3HHXA5MwF57/s/3qBE7oXVUJe7emXvZGbh+NCY4F
i5KVDR84OPti5Bm0d/jeo+iop1ONaAK0nzJBpHh0xKWCnBkXh+Xxr/8YB8PRJUia
vDYv+FguWx2rpxirw/Jl/SqZeahhny6V0Eiajj8/VsUp3GsMIS1KCgZsQn533Y+3
5BT3LaI0ckWWed7X7n8iGwvU4qTvK/uySSkW4n6srJ++XIbEWr3llP9Arq0fRd4/
yo14WAT0lo+fpcCUeGqHHjl/s1lKgaHb5jucpS6cQvG1LCep0wen297m/TqrZCA8
YcLZuPOAdTAXZ8W1hpX67fCin8+3dlkRUhvBl6r8sqSwroueqOoVBkmyr0Dg794B
bNaEU8IJL1DuIwVYbgeUaCUU1KSVeL4FL27QkLkKSYIcVpIZI0FpZ9opUAtrNfJX
T/2tNByQZNrvSIwnjwIEcfRvsvS1E8NfkcRC0A/JkD8CY5HttAT7C1duYunbo6bS
oiZrcWXrjqNWHv0IX1zY6NVHvpgPi2p4c0TpPsZZcQ73OuySGh7cm5K+A7gJzKLp
UW7vbv72wNwPiJjwfjCykVhU7kTp3W1EqXQY5uIdl2pFKjUuQ37LuJ2Sx/AIUYUC
B0998GPF0JUufpTAxkdMpv+LgTVS4gee+IkJXWvskoUzsRRlQAQ+QXsGbmy/no79
g/J0YF5F0VK7AaNeMimmi7H7rGeZY28YBmGFj8X5jjNU8hkVTeff97D3QUVhO1p8
aTPfTqkob9+f0Z7Ow2+mILdSRUCc5J2QIS7vSBLF4WhthgRK8sgkAnZFLWcPGiCJ
2SsYT38go0tbClFGh54U5UYX25Jnltjli46K2IEBMm0KqBxn5oDoGG5VzN656LhD
jHH4rGy11A1eDnbHuIpAcc4miHuZ+9vifA37luzaD1gDO+Mc4nWFsBcKH+5P1435
1eI1ZjECZtPae710TEb4qVqvnMJTZCMuPI7kKeg2c0KxRxLzbWjcfzSLksnflPCE
lW959r5kB9V4bx82i42SeYchT7kDexm+SjG1n1AYo5WVCGowbZbk+pSVgLmqN1Bf
KyjH9nQG31vtMKMlvkq+n/gk0Puvdnxn7i7l0ZwdeZCUOhbp8XgtP20xw5Q2yQl2
9pSUl09wxw8szFXBNrbxkt5a03Wo1wtLjyXLo9ghggx82eLRvzreBa/9MlSLj2VR
IZyoxK+jF05cthDUSVoGtXWJfBLI7fPWT/KhWy6/Mv/2UhTpJnH1YUL+XQGQqJUi
F4k63FFpKLvxoVpcOdvkfiNKCyGGHiYI7J4rc0eg48k/KsDqY0KdHZ5GeiL7dpIy
YAYCfmsK93eMbpCWkMSNvpQ7uAZ/Q28JHewiuJ1uAXcq2o+wosZB00qJOkpe6xxv
eLhDwqDEwodZbZeFf2QBWcY5pW9LRdAPAvXMftWadl6zaiAtAlFFweOvNd2iFWk3
vOx2HXyPiq5GfsKs058Z4cb+fVJtDMBtH6KtfB4T4fChHJMPPhV+QpFnQfV8s2LZ
r2v/yqCuFFouAQyA+E4HO1UIGtyhCqnM+3k4b5ghF3mgQoYUM+OXFstQzY0NyVQZ
eCOH2VAczp7pZcoybEzjtq/6Cah1upue4b7Lk6sqIBqPnlPHZlKJK1az96AAVc6h
2XDzKjbfSVLKeBniUJGO0QMGqtBsaj/3S0ckHfAeoksfyZYukQIE3cVjCFInTYGI
RpIhXljFz8G/NvUvFk/SH6463klbO7lmSXWlQK6hhd+XheRfxrbqBiGOzOihYo0k
/BLcoHE9NenSTUkvH3hCCEWBvj2fczopuq3T9U0ZZ5MkDsCAdFh57/X1o6uKcxWf
BeyFtBLF2cI1CAyWIHO8uha0XJq/s31EXs6hycIpX6D7UhYoppGpKsgCWis8TzWj
5A7jl7VR5uNWFJf9Ttq5o34hNGwewCOO/N8DH2sPXVcO3b7aPgQixXwocMimKPXe
4cwg/PB8NwkrfDsLUGvOOtp85SiAgoeWkWrSCKlUEgXM/6qq2Se0aY86FDGFrJEF
fjHBd7IOk/vwbn/0XDjhvxSKNL+gO7NaN7ocIHZIvcp9jn0+NQ+T5SuhHzruuJlb
G8DaK3uXz5Tz0EjwxpTztEviJzrxLhGhP9HhrHB+FDGEnOro1ty+ozWjazGVVndm
r+ycUpbvde4nMlKtYDrT71eUNb7J0+Ph9v+pjkH3dmbqBLgmQ+aDvEOsDJFeZUct
AQBovDd24SksrrkfgTRUA7IeJLpxo7ek4JPXNUVH00XkilQXhkSNOPekLTANTAEN
XXYEGd5RiEH6mk5iKD2CwyScPAAHEENbffeDbnSCo2fS8beYz/myl1fxLB0z6WGc
XFmd4iM8RTUMokpl1AxY1wNFTQyDwQWKvUCa7S5HJWTNx24JiEbfu+1Wj+rR3bu0
2zOSh3N0qM/uNywMXmAPge9ED8RRvdRjc0oL29jpZOGdMKv1JFtSPi1LHV4oMjrq
IaDEwaM4kgUeG3Qd7sm4nwnK2zUm4j7j7HF+brw2Pbm9jFRepaLWbJJYdsc6wIAw
HNz5a73rg4M4LoyXF5jl4RjCJ1FjdqoYJTk44VlzSqnkredTgHVlbItX3Qv/SK27
RvJjPawhoAVrEyIXlDS2Fdi+hlAnCQlIf/NSJqzqS1LuKxrTEBG25vRDRRSUPkFP
Dyf/yrNOvdsRa4K6sCWmHyH2Qw333zabNReAMdetAui9JtxIWD2yy8lTdWOk1UBk
saa4g5niCJoSgyWHl8Y1ygS9o6musQItGOUtM9TAsQu6tuuBKaNcxMwvAeufGJRI
Djj5Flo9zPtow21YD3+Vrdc8denDpcPqLaEmXU+udEFakMMY47qqJU74nlCbjizN
6So/UJRvAYJAlZYmJUv+AZZqd4/d7YUoJZ83Wa+1QarrbI/17cuSJNe8wj1Ui12I
j5/qVgHlLu2Y+QwkOHzdCWYnQPqkhkHf9Z0t11LRKV2UxcwTiV14M2/n6sbAQbSx
pLEWEV9uZguarxiPMiHKxlcz5Ij5moZf6TYLtexo/P6tZjtu90T8n5U1tRA4mGUh
THurX1g+TXxfPnM3LMg6kIauYBuUWtVFbR5F4A4SgYKT5x8nFXL82nTz8/nVs39W
MhK6GG/GT79ExiwxEkbZiQGgsysD81wHykvfgvNyseeP9SG5EnD0QYue9ML1Nvyf
VG0+4DtvRfF4e70Wel5ZQ+ftUiDHk5m7k86EJj4wKXDGbtFKKXq9xDqrPOf0JAZK
f9gU+8ADIpTOZ3tM6AKwWqOsudlog3EPyM+gvujeMx1ofi5cXwqGNNGLhRNZwdR9
b8/kw/ONcCFUn+gBvP5qMLBTeVhaaoUh0e2KiKPyIgIf7oapQPa/RfRYvsh+UMRD
vR2jzElrG/eN0l8kRW+L/ud4OlLiAh/Odcxp18J0k3ZeJmY4OMB5HfLYhHWZeHUh
GT6joWtN/JobN/QY6vUUHlY9+SaETdzGbWl7231i8OzcdqQsb8q4abYP0HGSJJ9k
/xGG5Qx9JG6dI2ewjzTc+kNo7MPwpzJuMTOYbdJ/1By14tMSM9C3zqhKMZY+PvVa
rdAgO99wrvkTMWYCrvwtF9vioEpWyu/vhKWe9pZ2juSp8J1GhzkNcotJJ5dkAxaL
c1qMT2M9gx97Yno2854s2/5LfYDwPXkwQG/tNrGTN2O7ts1dc+v9Eyozb7heI4+X
aAUH/vSzEs0AjTsnVfN97KZhWxuUne5fRINgHqjTXVc7J1+lPiELyZNe1Mtr1p2p
C3Xd4nJMOC/RAJsM6qoyDW4r8w8RrF3F+vDqTI0Vu50p+QqbRXB5o8mwkcN+mf+k
RNMzpPHgHUOsdaOGqZ4lRX/OrzJAEVVqJBkwUYW1bXV5kRls8lJ5mfUbUyQ6ScdF
zgHb45TgUqjynLk0DfFHcFNlPV5ZcF9UgkCW241+1+WszIFrWkVW2qRegiynJHtL
/Tzwy8KhCH+vnVH9TJg2m+ffjL9JtyhMsttvAUw3B90QvSBl8wjfrc3qoSyfe6gq
E02o7BmwHSc1Aw0kVkIKUywZzEdeJdg8q3icwRDLhnH+mPTdaUxL61CP0zfsnnm2
4LHX88X9FOKelHw2pUPVIHEsakPZQADYXkKquE5Cy1XC9f1N2dHzZVBytH13aSw+
3VME59udzh81LjjZPV3uGwmC4gmEDODdyx89+l0lSbTe4QjqfxoPCqFrXAijOqeh
LV12V5kyVMtTC2HuI4oRadx7i4y04X11SkpGbpxW3WvVczB9kqhcWoceAefNyntF
JGiJGO3LlTXsuUw7gq80hKYN9BHy6rnx/4hY5L7NDGBT0nzBtq0LJwp5h/HKgNaY
/1I4COOccLx4vnXk33fu2awJZo87pFmKx5VlaJ5LT94H+T9J09Y/sdevWj5e8BZT
r08cDDI7yo5EjiQw4oY8oqF9HPkxd5lsuzS/bcveZSX03qq9jNMXF8ZeGlJKkA0L
rJxileyO/bj8ZOLV5wG4swf5LfzH/O2vUDDzxrAdWZMiFFGnJJME8KUCSa8LhqhX
9TaBnC5UyPNKjDqT4ceILzuI8Ql6GJ9wWC6MaYdtckqXC6PAkEssmpkjodQgmRDJ
A9BQhxxJypUOrRh52S7VuQzPQxLqSCtBDTJ4S77jyvyjerJQII8TNfHD0XiDH8C3
M1Q8RsxhI245uzIneIDekYfwDQHSYy7eVIp7dR4cCKP18h+S7tZrd30gsy7tmOYG
/pC3eHCizpx/aDvyglFbR850f45XNue376CYU9EnfF90A54JHGgFHZIzsi3fWEdd
4oG/Nvf8plfAsIu7lGBnFDwnRTIt/MDXzuiK0Py30ohNLGtLbVPW1p5uVziSA4Ef
F4Btq9f5pYw2vu/VJXhUdCv+dgStOUqg4j43Rbj31CrGJSWq0DCA6+Cu7YS+7sXw
7B2fxHUahep3/mG56kIOTH67SsejTxd8R/G1tJ9XAhJRcob3ulaFb0WC8G2cIVVz
BYie8Bnd8pI/20D9bhpm3Jzlm0k0nZOAbNTZcckDEu1LJDQl71wEkFzPONVbga4D
jLZPubCvx4XyaYNxBwZY15hQ/zG3zjp5N2gOpqxZNL/Xk5rqNnWJ+Vi1Ay8W75FV
GYXiU7Sv7wL4TLl3CIThu8aVv6yGHe+aHn0udgNYyUdUgjejMINYbahsKeV51+Dy
DO2Kw0sd11UsK5TRSsR4PYcMk/THDb3lJEwSy1XJbFzUlcDMxhWNi8Ax48+uPTGz
1lfPqq7ZvhENyFASFUc7fPNzTx+aZaMtwrq5ENoILjG4iWUx+DZo/HYhVfzRV4sy
oqRjQc9VwG8zCkDGAWEv/k1btzS/k6zxL+4uFxIlGFCuhgz8Y9X4RFP2rIiT4EGd
b9cBZJIJu9uiZsu7kG84SBQNvZD1TvOw6Zyqh49dV/EhJMyU37L+yiw5c2hrlHtl
ubaDXVtI9TUgtYyBgvl/lvifndnxC7SYzVbXNhWRZ8j6CskEfaEKFSA4LspAAM44
PxcARU2lt7h/jLanFXOh8lSp8II87qKrBk9o7yZ+I+PoI8nF7rZ/r/6JnR3tZBQJ
RtHt/pP8CUGCRt573K5yxBmlid3IKAY1X1FNJEcl2TEFXXb5KJR8lerOsm+rUF/t
mce815cxKDEO4F1+CLSttTbFXtfIHQhg8tlnG0ixJ+BpMxpeLaZ0Q1SicMrSwL6L
vwM7Ld7Rh8ndIHRFTHGerri5cHeNtq9MxvmMstVEX7zgaxnNh2sdpZTWhxlcYIe8
j3mJMPln49vPY6tC9fct6MFtIeFokH0aDuJ4rVitSc+758/6qFXt0ZYbmS01t5Y9
klXwJGF8jn5cnrW/uU3rnyq6j+2WGsvfZEWv728v/UeOsit8P5AjQXSDcL8ZdvI6
3wZwzRsGT0pMH4O8JrJg7FaO0OuvS+c4ZtDymPRWSobTZxju5W8uQWZyNruqsj30
AI9qO12FlD56Xn2QxrA58uxuGasnjoG/raE0qigVKI4hZqZoxwiKmSBE1rHPYeB0
7kTdpdJii7zheMimo0nl4OBEnaKVWl9JqtiNKhOSBPEPZXU7eSsB4i4C6QMEqxW1
pJTH7gRKw8KA+3zR9qlo9aTU3vJOkWX5/fWA+6VSU31ytIVzy6UX+2TTIQf+MVCp
vzvJdN/yUvD5OgfSdhNp8u5NTyC5VmWbx6u1UzXwWsH6gsPDeNokYZqgrIuYi25m
AGC1tUlrXfwj9fUdWc9LUYyODdrCdTzkpRze67PS4dwY2gL1j0EWXkaKN28VkKZj
+BybeNlAAgkC2JKHL9tT70yu3zs7WmfqIovxG7/SgDZKFwjqVVaqk2dJdJ90+2BT
7sAblVCS0rnl4k8/WAZF/wRoy/OPMFWQfOKVTz9wjx6bjfEpk807nFRaEg549gq+
sPpvOEJfFM+5l/cRBgoePqq9hM3e5aNFWLC6JWRT7sZ8aH/kZMEveuwtvfKAht6+
SE+5Krhg7r5NtJxOS5A4kazObjS5C+9b60zVthl13eDlk/PpyKu+ex0O+85Ekcq5
Hy9OSUBScBIAQhH8xBVkFre3qAlxryiORiZCBMXZ2rbvMAnGg61rMD7H8R62CI1f
tC1WIOy0JYOBYYC/ITe8sJK1wJxbUebiN25Evpqz30GJZtw+4cncO9cTZMSm+SM4
HsKyRCG5pL/U7Ts+Y5a4qnZFbXhnyakXIAc6RyJpVyeL/9RQihTwqPK718zAmhRE
inLNUgxWalf9Hs6XFZ/b8icJ3DGExphTYixR4cXhbxTVsTitaJlRDPIJlhOUoTe1
J8wC1az8VN9IAx/fzkMhIag18Na6qlTZ+c297Pn07GZelPy2kOUHFs/UHFNrirHE
X/w8gkIHWth78C802HM7wgId1f8Mgl7mIp/erfmmWFxgipBj6fpRpmysvq+DaIM3
nEobDcL8V/ZKbsUybe/DNb96q0S64NdmlIDBm4VNje/W88jK0fqgeVhombkty5pP
Oxq4DO6pLm6U0iIOX4lhrRevMbThsAxaE4lQBS5NRb2lBCoWmfkU/02qK43/JISx
jXhLBvaZp9R7gJeJz12UtK5Ym6fNdga/3wI17AaOtPBwzNQQ9ShmloIupjeQ84ys
bDN+IAFoocWfPQDCX8dWQEAljFW5OJYKOrRJWsm02fMJUheX6W25LkHcH00wagBP
0EN5eh1ishKbvKAkPDWQ6/bDF+MzRYXMtQQHv5/ZpPUCVHxhmE6KOR3EH6YfOLXd
j9so9fayTvr2ITn0Z6xyb+FkxXDZXugIREkbRNzl2dGjJlmBRTkJysTQ34DkKsjX
fNsamLTt7v/78KdclCmRE3juJZBv1eZOwvTF6jTxmlXLmsvCXpwlk1AGKjZLvU53
uSIpw92M1p1nFdm5hlegbDGQLC1dnUTsYcOa4Rkbp435r3S9QJRpdtQ5z94E1sWi
OGCi9tBzEkZKdcx28MFeJu5enH3OJH1XfROU8bvXYJgk1KelyvCT5KrDHlKEsiqt
dPXGD6+Qv2yftZXNet65PyOESsja6MQrwWX7CZsEBvhkb5viUP1yzmsNC7XFBSf9
LE/103t43QaSHGgxq2yyKIIFdnL8KwrkdIy63yzAOifuYS3lRM64+Ls1JiS4bWu1
W88S24mcsKxXZWHbFPIyRL/FO6txHubBT0ni11iiJLXIN1gEE6OFwgPodRM/x6x5
GbVb0zvgM3uTWbkM3CzhNmNYUFIQjj3MoD6ZNC3oCmhEWhM/JdCw8Q0622/x/DW9
6br0roTdIrp676UdHp7cKPs534ltlFNalgLGPwf8bWe83exBgja5K1ww1+SCUzfh
3hBQMJxv9o3dVCNmQnUKGTQPu8gggt8jmq8nsWNz9bHatRbkVIeD6uy5MlB6kizf
9lPJ3F5rJDGhrzmKNmS+xj3wQk3CWj91e48ayqQIoSd63X0Cdudu2SbGUT/7Eqk0
xOo1yrld8+RSh3uTyz/BQads1u9ZK6jw/rDiFGxIzDGVT9/wkLhW67zYdv3b7Niw
sMzqUftYN7DN1AtNCSk4iCvi2lxBpHhOxfvcwK/TdlhKPWwoTkqYxp8tLOMyJ9lO
V2ld+jRrm3m+x24ShmhYqYjFs+cqZB8VVFNYsuEtE60MDmF3bk17xFe50GBEjqOF
4RXaa2o2hmwx/kKWjH4L3wwK13yhw/t9CUsNLz3rTjJ8YNioH6MkqZT8XRaj8Tb5
QyfXH7SMqlVEt4lVnravlhDBnuLuvZOKgUdHE+vZoB8SZug5KI7/jiJ1wqzug6oT
npSJQR0MLuBKiNn+AvVGRHz8yX4o9ZW8NRNyAwb4faH0y7oYjEOalNEE57r+f9Nv
mGLS+kKs51Nl+FZPz0YGAgz4seZRmcj6WixktzGrLofgzSCX7z5oTip2IAS9Zppc
133HAVQ9F6NFubMGA2fWM/XP6QmOLbLChtDvV7Lq/IISVXi4olKpSnNb2FIG/+jL
U47TCcczzb5G+l9MYmqrNLm77pKUrkzQoHhRqF99xwkYVjwM+bk7qvr/BxlYw7f1
Db8BVBoz8H0eNpShmKA1d7A8hWKPp7YiKNTkcz1NxzDuEyMjvV0tKUtPNjoEilIH
F9vRIIrg2sEOKk497JC12M+QmIfaNjfeaZTMOnQNY695awvjqJTHFYlHEQTvhTy3
paM04jAnmJl3CVCT5z10sh2T9BSSFTCAJTWHdv9C+vTdfZbxwAII7OR8NutClC++
bjUOSKQJdagJudbzFaAP8Cp7XhsFPA7WkN1PxNX3VEBr+rDz26BnHtuk3Vvulz95
1KnuO9kUr3475BRmuhqiV82SIY3LYu3bnm1e7UvQEejx8Mbk1aAazeo+lTs3wgh3
oRuc3h4jJ8/8EWn8I1Om6d08950MICnyXQfhNGzrYM5hh+KkBRjLZx5jw4DtGobH
LMbiTkq9CD2vjHAjcw6C6HzX3LPVmsaxfmVlI4RQIjAdsFPp/mG+d8cq2pVKHDX0
4kGS5aWqHKqVrUcmNM3z6UZQGiwGz1/UDn6m5UvLHuD3x6BCUQfn1vP1YWeLUI7+
cTf2aSkhse7hs51TvOiu/ewpb5qs9kMDDXZEMgeIa2Hm9udYG2ahnpzuaMjsG6bL
YxV+rPUAT246yAlZhmxpO+ryBE6EW0ivm+YnBkdKhYNFa1T6BeYtU68AENeZFHiJ
K2f+zYGdUPA7FwxMrNQdN+280CCO9PzzccQs6HoIH3MoAyBF4bL0ztwqa3Bdpk7I
R+9hmRKmLVmFM2wKB+U30UlcTDDeDYnmDgSL7Fpox1dFYgc0DI2jiRLqCzcomMlK
gNvXKJLESnH18HD+5vLmW/xxrG9ka4fsn/XaKU8dwzWTxLvncpJWkooVTG3XJqp9
QgwFuaxWIXBNc6ZY/XlObSDtocAt9WWrl8O6LhS02Rbk6tqllpp1OvbsTjFho8Wo
BiiPlWj5NENNIha8+YN/+0JnneLTmCdoNb7R5hRLwdSCKGGqCukzvWXM2KVXzVdx
7CJXzEetw6cCpv0ivobGq1GyQD1Vid/4D7SnLw/NDWJ0P6gektoWbVXSvC4Vt9Jx
Y27E/+oaemuWTjcJgSQr4TDuZ2E8pfTKtHIdx8pWm+wgSmxeQIlX0Ia6INxscD0j
2sOBmIh0+WXLTkUX3OiQOJ7C5IAupYjpurTf/dN6hAy/D33PnYX/WaNvJqEx0ms+
+ovb7h32jYHV6ExH9s0zY1t2H0C5pdwX/iXl67e+5PAs6EK7UOn1HSiArMN91psZ
GGmFzc/2M73UtywY5IARZVIeiOs+ITERcrlRHj2qUu2jyZkSjMOchi+1JoRscpcb
D+Sdw1fJKSyWc6tohD3HK9LiwhGve6Otbn3lB4WJx922aG3beZpSRnk9zJA6aQ4Z
L9aWlqJz/vvhCekmBqoHaKGLyx1IyiUb1qgl1yLFF5/squIoP+DVWwR3pfVJW9+o
PO0MLFAHMTUHLnDiBolkVbZkogp24CIA1MqDaARJueNV2YTwlsLR8fmHqLIcnWf4
koRoB+eVTCClwOyg0H6Bw4Asp0ahjzbm1Y8cc6uhZh+nOHoKTixBA5phtZ1Zc/pJ
ar5jDpjZCMuhjlvGiUGxqBzwhYxgFSB9cvilH1q76JQnek+PeQ7ucCue5f4u9sJl
289wHRqgx9hqD7jtSvJjQW++TuuBi7kCAGs0PXT1wck4ExoSwweb5GZcRDD8qIB8
HRQTzxh//38enrZSRTMwhbjFh5qKBg00VWv123DM7Kd07EEXzf7aG+ONbYFKNgbS
SUW/bXAWmSbyDzc5TdqnWYFNxTR/yZg28kZRfJOPWlfDHSj12F24k2wqgBOiTh6b
Ue8S4jLjABubMw1Janpo/9rSzATN0goXsBSNSzP4mjEmrbYZqS9a49pQ8KQBoMxx
2N7BGi3Xmy9/AirKk/IRNYN5V4vlDNAJ+3MIIgEtnHKow83A7K742wiHskXMzlh0
znQ6h+CtU0CDxwnw/23GYHd+X4QgbAic9/rhjvrM5ZQzYiVD3Kj7UHWvMJK2/Gza
Acg2B6OtI/tqgZ8lPIJfAmZXdhC/x975qnCDzPY5lXeRAzFS1KfNEa1rX6yGudar
4oV725FD2NH7vL2rX0I+NPnf0SByYo00V0/1AJwcfEzB7OD71lGN+Q3iA1bs2xu3
07SCLj2V0Wn5DqpJVqKc7YV/dynmx1YatOqTOTgqcAp+zRIw3RAXEU0IYQbvG6al
6rDjFKrsaq0E2O3+m9usKBo4Y+m/EHhB2QPjRzMbtU/NBB+o/voKXfBT0zNNmmjD
bUMLsdzw4CdJNwPpFsNzCtPTmDucZskNw/LW7RrM7r2MxJ6VOerUkklVkv+RjJxz
nVdyiHImyATJ1t24vLWN8jQFRnf2EXA1XHLd+6msH1hVntX0A5+FE7ASQ7Blso83
uCTC5fNgIBTH+0kj2Hc8FupHgFDty+gBu0o2hBCnSkulvFEaTUCN24dtL4lz26rA
zqTLOudlSOgSzIvGU/OmcsYyvagTYzmR5XqGZMm45qDDEBCqJFiq9nJEw//yAiDC
6TvycIlr435M2QI3qIRf331YGy+4K6xCfY4jGfXCSPVh8rTTMJem0sicMAYrOLkp
naGHiT7JReAMZ3u5Js0N3P5HXg8DGGWAsAV8As14b82rtnQSFk5W2Ff9ujW8Fr7s
cAgiKo6RWvid60n6vCGc1wV3mJkevnLTT0td0/reIbXjv108jt0Zp/0Wj8H+a115
XLCWqU8NbBzYF5Dt811lFD3s+b04dLGJ3EPjev7PsGnIKVx+FPd1enTumtouHiPU
rw0qXlMtPkRD8w247yuWGDrqXfEZlJGn6KRdG2cqNrufno316uFB0Ii1R1nAXuPR
7fOs2PrkS44v9U/jTi5XzBiPhEKp7DoVDs1qWKQtP6PHKnuu857ZVKjm228OtyJC
QRAKlaC22kBOPZqJ+5OZMeom1gwZwsATe+hIRvflWBBmlIQGSNC1EaKmpGnIZ4xw
eL4tTBVYmyFh4OiETGSD1Xfmh/sIpE7u6D50IDif88I02uirQZuZuPL3nwLE2XbE
bzfE7joLajbgea2M+z+5w+skvNRXHCDeHS/hrxfN8XaWtEafmIWCfxdfmrGdHxe4
95usdToQqZrtz/m5xUMlbaAL0MTVpujMwAltbl+7SkCv6/HA+abxq0NzWTj9itk0
H4ZrQwyEOLt/ln58Tbv4VJDBNUMIyAfgQZG2wPGwN5Hnri7UeUJz96lCLpzPF40M
c/t3ZCm8coXneQuh/dHMPxS36BP9tt7uQ7vZmPB5zH24LlMiqF3yyi/bQ7Sd5oYh
H3KdBxS9Pt6mkTm3Jc8NkuIlDGx4hAZvqwl2UXmB1hcgdQQ8NRPh8IRhdusP2/cT
N43ognFwq8OHfCbZCewcPGCendzLyMCK50RaqbmbgAJmL9jA5tlrSy8GTTD0C55D
lZbORL5cLRu3tE8mEpA1h1IO6xTP0hxO0gBjBHuQfwRg1yCr5b4J6cOOc9Lf14np
NQJLU2YTPiNugQwKVkHstFnfu9gU2rMtIv4N+gZ45K70MXVYmSnhOW0Ads4Gaiy/
sLwL4cB/BxJCao7fkJg0sfpd/sB2pTl+qsduC+iZVZY48Tvh6yFf5FnpXKRcKlaQ
0HR41NOnYqMawG1a2vwuOS434EiQRMo2IUb5EN1AVSGlVzBWPCtMNNfPkSPSH5Xz
u0XtJmLcCwt34CiRAHXY3hPgCnFaFY9UoLEPHZn/cpjCJ/blZ5Cw+/hovHMBGbCN
IUR9rsCzC4Z/EvhjMYRDkr6q5AUYdfN92ySfyt5TFvm65cJ1c3GLpGFgwMEprc+U
XFDJLEfXT4mhjndQUeJGwORoHuq8JGd5OS9gXL4h1dQNQCOHoeCWObSh/lN/WeR3
3nb/TC48dYU0erAyaLeRRgQBWPQIiAUFph4j6JEOUWWiKg53fG52zjwzOni44CBt
xUqr6BZ1lqOdI2nFkuZ3Kn4bvP/GW2BdmtMWakctSLs6f20O2xkyzquxe1cAoNzc
e1hXx5bO6JIZ/0Le3Go+/724/k9sBtzeh0jQhgqG4nCuEbcp6TOf6PeHuQny/8Qj
EatqdjYYD8FGkNORzYf2scLkzvIYB3NEY/No53k3G81NjPs/RwmoiJ88qb8d/cp0
h8i2yJK4m5/DdH0fkGAkJ9eoqERl4oZERTLj9CgLYPeXK70IFfGqzqbzgWfx5YyR
vXTgFK0G5H5EFVbzSEcq822aNQvmBZsnHWbQ1chQ0kqF2+RfqHzuFm6n2Zx3quQo
IKinHdOEJ4wIgRY0QSaFDoZgAkOJTNEQ9wnVET+XnTzKy/pNVjqamgPjDqDEM7RE
xKytYAjYwmWgD32nLEV/Yn2Qm0j+Uzjc/Yb5ETUUJ02s7m2Jy6dRQwFf99dedEVc
EEtF6CtbY/7wq04/0+iwxu8HyaR/b2U/IdmWYAxSbMiLNiGE1NuyESYJVVliCpBe
Ixwi7y+IbMGpvoRRHRj14Ug3uQ+btkHRU/WGirLa3Y803jQ4ABIpPCCf0xsHlYnu
7jIF1u3kV8Diqs/vEtrukQzPnLqp71mVEfcf5wOlL+QTDLjWCD/l25sWKd/28hNJ
1GgBG+V/Hb0TAcbdP5FEXSIniYFKbSyAxJZOGvKL+QkEz4A2W46Y8/qD9O/xkvEP
FhDnh281gcpL3taCaAAeEJutYQhppWTxhfyvWPC0o2ryZ38JvqeauiwueGuhgk1l
OEVXpaBFoJVl2xj9hR8I0Vm15/SS6tIAQvkBTHwnE3YBcQvEVpjtptgoI8S/mIsl
KGuzUyPqoMwUpd5ciNVCL6+3kkPNL66cwwVpNVAZEZhQW+UsO5EUJ9EfdRgfG4RI
hn2dnpa4GCsQxmP5TRnGf36O8Cr4bHt7IkC0EOplSYSmKj24pQj7UNRTIa64tH+G
QZ0nxSgMlDtT818OtCCJgBa+VzVrvCcxbTaqX44BZGgKRUqTktprk+a2fkLVBxxF
qPl3KnP6hJLMh4Wcd6q5L0bxdcyEF4pzyGn67ZbTXaT6Z9Tzt9TVcaeLLNfQAD9+
ALs/yDozS5qTC3AEPJ61226Uhhu42nSno+hqVzQpgk/m9PCRbO3+Vb1taoSBJeyQ
A7xW4qW6s/yduAs7wgBdN6LqKwlW4fP5TysBzKV/6KncU56kwcRJqA5fFda20vTd
Y3AhfUP2G+AKdbwa8m8pY2E/v+UfKDMFHKUQYIDJzw1yg9Ikw6FAYyi7ga6usJqm
KmFgHQjBvMyh8tV/kmOIIr0S+ehpl8d57Q/U0j/sUkr2LbDL78xmsw9zoQg5ErN3
H+/z3SfBUOOXP4nqdc+wWmW4hsErtuSgebwSzmUP5N+liDKOSM5e+i5GGO5dqyNA
OYYXNetH7ZAeCJIspxHiRIvHGlLZW5/RJ2XBa12Scw+/w5mXcSEYqBPsl5JTEhQf
XBgtu70pn1U4XCB/ImURk8M5CU95XOkGLv8hmfn8JJojPwAVd3SbI0mioCvCFRm/
82BUgMwsznlSXvSYbWkwJ2ak4lY148ksIG+SNu0TOLggVyY9w/y5t6au/Ep4wels
rJiW0w+0p4MvfLRkrJrD28S6PQdum35Ka0RVJ9m6EhJjncD1Y1qW919LBinE8fIH
AedjNy64d0jpmskqfwJ2lBuQCohJ7GjuN+S+RTzKelZM4EVomdtnlS4UvppllAO6
+89LpLq4CjhfpUvYhTBIIWHDfpjS0ZzmbCG3ZSi/5Y66R3fkIydO2qfGFp3gMWGG
NA3vw7Phy3TzqJrCY3DbpWyrHpQ0ouNv25jEly0NPxlgTbg5mH2GxNuBUFoie4eD
hUyxfJTkzY8JXt8WOBpGOSyGQRuCoxhKJDHxkBafFY+2Nd/9hbKTCyX4w6w36GFU
99mx+SYB6ss0RskTCVUHJsxcEXy39AFs8FvKxF3OhfPF5JJMIbXMCBsruktjnhMr
rfjFZkz9YUoEIK0dB123lfcN/vS6vHKf9MkBw4FxAS1JycRMG0yy/QL8EQhVZ7nj
8QbRgEO3ev5euN3I2uPbN2w7TVvQN1+rZ4+CvK2zQJ7MWLA5+Uybjd4tHlLYBGyj
Zice85ZAwBZ7lqLPGHjckbyKEzKwJPlW8TUrwJHfqRDBLrWRjBwAzFK474BS/gUL
Mi0R2X5ife1TP+Ybg3c5kQnkmc0klEoj9re5/iNWIPoJCCroOCzgbZHE/Ki9nVta
G8J2TrzzFht1S+QlDhCIYbeBFXc5GUPG4vcQ73Se5AB+o03EZQLsAnBLabhTfl53
dCMFa/B/sTptQwTuaQiOWKkWfcg/b1dL+0NJ7pGUqgxDQNP09HQnhI9loYarWaN2
0rS90vfVdLMx4dUo8xVP9XC+hJ0Xh0gfHKe6ooMO7Oyfnhwr+M2SqhHgCpJArG4p
X2TZcGR9M0LKHEHZft3KQlRb9sB72wjxnHikzPm/LnPFaurdOk77Bu+XvtOjdKOj
ht0x2XSkNgRxNuFs5XMRHdbgznGVAxmQPcQwtCNetQ2oSu0xOT4Zg2lnGZ1bcsAg
gXDhPLjQq8TjGIdv/5BLhAy0yNaEZ6Ha267H0sEghLuGuZGmHf+2Elmg67g307dp
DuOKksn9hjQ/mTKUh6wPb2eU9J12QDRZdogvfVLG+K6PHZYU8Y/mB3nIi9ECFtho
ODJoFzGVed74mftTqOjGNtLbIXMDGL47z4dlUOFMHXa0mZS+uEm0JtUxEoocPWIm
XGdCWcyXz3Ieadg0ZE7OHxT/nuDuPuBT5AfC0inu+HyUWCs4IL+EwDyeEcuB9Tvk
cTFgG/BJNjf/92ylCj2hVlInvumLabPabfbTqGTE/6PupFAnQKrRTml5SFJX81y4
qqLC9NZmQvY6aptHPNevXlxBpdOVhMWU/TGSfsv8IPWl/8V0xgiOFDrprRBZ06OP
/MqxdDAI9MxDxI+ZaxUbi9Wq1vSW8Hx/sQTuRVRzRE5m6+3SlUi5VqZq3HaLk9CI
P2JlGEX4Qs0zRs7iSQd82dv8gdvl+eLXf1kgWLHxj6HuQ0AJSGE0o3Cxv1+SRypC
BpPoYVnXkdhBCEENWV7mdWoK4YQXWNy+NJuvSe/nJCJAfBR1JJvbBQGxKP4XwEt0
INau68k48XfK5tLXpCmQV500P8pdJvBfvDHckXdFfFBa1faJb5DC62Zos8sTpMM4
kn23KQ2NMlAt0WCB1Y52a+dwqNu/rvYMv7UuzmZvXn0aHkrN1NFKdpVHDj3FfZ8V
7gmA40caaQ8mjgA1dwlF+yEO6d46C/KT2vmaHK9CWrQ3cSPSLvX8DwIDBbwOhnJP
C25jgLojvXKgV0UZhxLqVII6taFZkzPaW6qwuCmki2aicZaCMsNb2+tc3kHYAuZW
rUe4Ri0+l7io+mAXiwjK4Z0a5eugFZzxP9PckrIh6by/Qhza/8/qZ5x4Bl9xzeJ4
EuZN+H9RGg6sScHgNnM9PqKSd6861nkE1X2B96OKBwss9sk/fGt+B12lpoeVbNNC
L9fN3RkCycIy3RGg63dBoVEjVmThmuGAtL+R1f02aQYkNnSY8lncCAAkQUjWu70p
301zba8PdB7Zy5VPHrqT+azJ4t+GANinXb0hpQHZyvsUNvVjd5D9SkR6w4MAj9sq
3mUB8QToaoF75zyHj4px8pBASBEa+lJXQckGNTqVasDqzZb0Qu2wfhgMpuP17xsk
D39oM/vWSn+SdgzWg3L9Rxax8KTiKWXRbgTK7jDMpzHOjEPZMNlVeJuIXg9HlQO0
Rc6C5S+6bfgPWQUp+PAFWStogaxNZ2OUSfjJWI2AYNuTqgmEF11VtGNk2DeBkrU6
NV9GUeWEsM1j2NuZ/lM+7ICh9CVxa3jVN0twobFTDV7SzFh/axRtK6cFFknNxFKQ
c4thOWvlUaXs6l+DfZ4P4aqYOLtd4z0fa3dTfmZvWY7ZbFGKQ46Rq494gxMaH3IC
nX5lY+CQ09A7j913M3tonJjvd239ocvl7s3rFBhM/QZIaflM0DgJTY98C0aLq9D0
xQzp8UpYPnDb8lk9ldCdgePTLOijItg0yhkGkCNCtE4MA8o1+fiuI4MjZmRdNZ5O
uNqL5DiJTrdRF1x+4rEIRsQqyBUpMoaCLaoJHnJRzMmfvxtod03l4fWBevmugYLN
jp2hEegaYJl285rlqQ9cDoZfPWElv9KaClIim2zaSygajzAsiB2iyOuVvp7ype6a
HCb5E+R6qmd7MkkT1tw9cZ9W2XwB7PjSn4RLWDeluWjLBs+c5hcg7kAVdJReW6ZY
0tmU0I9jVf6erBXtZleE9MPW8oXGccq/kw61cxeFkuzxtjlAhWab9K9szQhb5D5f
AnKoD1gdn0F/avVqg8jQXJanUNRnULF+GpuWNmSRnAcybENTe8YjRc1S5b9/KPuq
/8bWIC8ZFyHVjz8QL+m+GkUSvPbnv/zWtPzg0Fjkrjfn2nBykux/kFRCu2QZ7kYk
g+jp+HtI3dpWnVp/9Lrhr7GzEYCcr83msxTtL6ITQJt3a46CkfaDBU7z4wXqchoA
Y9YO3hHclzQDOv2pz7xWVLyCvkD4oz+P1oveO/xffm7I9LBUUYWbp/OkU4rmmmhz
pyYv+DzcaKmef48RyL653Y+nKemim9utwQKBFk65SiUiMghAvoFPBHI8u4HR56jQ
uMYc/71/mw+j4geYEAl3XAQvMBlHzA2y9VCl+3/iockP/COB0eS/W5e+cYOdLtah
+BxYN0je5CfGSeGbR40mVh3MNP+Ok0rirnema7lED5S8QARKdkJupshoACyueUlr
DOVRy1S4Ztd5Az7tiZcu0NQ6v3BZv7LQIZDFL5vbSaTSyY+ewB/XrPg2N/VWAX9x
HMek8FcoGR2gV5qLb6bADy5ePvwYxJ7O7m7+mS3kldybNDcopi208gYjvMYIopIQ
oP1R616Xx8+VtzX6JKuqxCsQWm55rtb5AwwQ9OODKWKU+TiMZUPwvgvqkvwnTjl3
XJgba8gePibnAycxtG9ItZLNH0y4As4VqrNaFSiLzDhwzeybW1p6iPmtWvU8ZzpR
8XO2rDPRjnftU0doyLLxYZsuOUt2LNYkr7vvlaTohQro5ihnEP28SCF4QgEz2yDU
O4csMDfI4dvbWDJcHrQS/92THZZvFDHbPUDGvFsf8d4t3R9UmTmVW7zps8duv46j
dbHihWzI7gRcnz4pq/o9BInAf8CUhCPhrW/bpscVw2uD3qUGbpEabaaJyJu4k7Z4
3k3tbgcNp39lPT5+0C4KeNAQ1iEOujixYsIRfwkcoqVO/98R1bqqQXKa4Jr6xjhE
7HvylSAjphA/iqSOHEUaVQdMU98uaURciS7nvszEoQMntp6jjAMT63Q0biwF03L/
Fm7WGz3vRVxkJMqL/F1oVYHRFggRz/EdooFA3ngIywE/LcAAT2EHncqLS3vJ/T3L
XclFionFMvPTK2jQ+A7heEb7/pJN0WfQilsPQrS37yqS2yglTQ0oO/r/KhA6V/X7
n3WgOahwSrHWpju9K9QTj+yZvXjzS0023vM2pg2W8hVH5t/pK7g033kFQhtZhz/l
Ak59PGH57L2f2v4Bp35Hp+E+Tm9pN0vCYghpnMIfs3wDR29hXJoen9PeYWFL50OV
J+idU5jzif1k7fxmBNS1WMNv5+hbCJRFOpto3A2U4wdkCZuvzlLd/XQbr/UJZYlr
FhHoNpp9g98vvYw6KNnMV8VIdyEp6xcqEiBNiyhwsIMZMOayAIL6hwqwXzH1K/sR
qnB6O8AGKpmcYQFBaD9RqwHjr597TWhupkGbYYFmICzFt1RG//3Y2X5rBUsws8K0
PHOimxTqwUKJO8N3LzJ+vvvlwKLdpj5yX9FiXYBUrjeqaQ2pM5BjpFK36BEA8sVq
pIKyO7HORxvGku2ll71Eg+bjXSrKsqHg8O6Ao41YCY06O0tC52hu7eAtGGWljMSt
vFPmjQwm/p8QBPh/K7XChAF+O3wy3e90THTRbht3NI5EYNiqAKzNAygRL+Fxtc+2
6x9d5mDLu5blVsLpOqgbQk4KJRtAoqPO4ZAfwaIaoq7R1YI0KdBA56juFD70w4Ke
Daq8wGcvPeq/2n+EMkoKMruQCC3m496xnS01IXiWsz3E+aCA5G7FIA2U1YntYvVJ
g6ZZ7Ledn/gXxcYyGws/m8bZFMefVtHzBqze8l2A4ksKOg+B487CEMFXcKyoovJW
dLwh7iarSmKTyQYcIwZxM2PW1Vq11Ofc51PpAN26f1H89jkmznpQfS+owmmaSCKe
6YddATsHi6dbyoUlb9i7H2GOBRp6JpOGn0Ek1gyJVjg02lhDL2mIlagIQJuxKqzK
qu53EBpOTEkScwl/rtjZCEAa3ZGk67NprG0xn7kgJA+J/4RrSkDRimb3/5DdWKqv
tBCxDfHwHEFXDAW38b91tm9KPVEno6nEX43sO85ZpMH/hog0zhyF5EiSvdNfX1Qr
pWi6cmwowz80hTWJAYxVGWlCieaJkZfHNgy0Awar0PeU3yO4nq2yiaYsstr1IoG4
v/BzaVDlQsH0Ln4d5kNFTIacqV+IIs54CLK3QjbIg4DaK9ekYUoR+Z+XQLrP05GC
v3P8LKcqdlp3ln8rGGOdbkb1ZbV2nBPqfnsG+SmgtgpArQtlG3wwjBa1o7Te/14u
UB8DlUGSxDK+7sJv918e6a1nu8MRNHzGulf3GcEmTycxtz/gVm1Mv9kx8L51Qhnu
KZmm1RQo5hpmdVIGpEhsEV015NdsN0/ApRVJxAG3qVUVoJuJB4F5af2TmNSsxobX
+AvZcJ8Hzy+YsscgcVeuhtkA9TIgh11Er2+GWFk/tlNvzfgkZEYK0EmZkdk4MFCk
Z06b/csXScNQE4tQb7Qjvocce1tckug5pcdQvle90qL5DLc15ySmt4rVPK+neON4
n2lExP+mNyyoEmufoBeneXMTslgicuhF3BISon+j6mKc2Ly27+Bd2CDtdg+keKCZ
fiNFt9PG16tun+V8D/QDYxgvDIp3cqapp99uMYnBykynKsRkKJBFdSZVqfPRrCGj
G9luCAKBqnFXxSHw3XzZBFiTyZh5YaD7xi4RwvMN4cI1A8nsJhzWzE//EJC4IovB
gQSM229UN7L39pggSRuqDcVbFa9uMYBPaNjP9UFCwQn/+u+i6/lOJt1tH4n7pS56
+E0CTuCXRexLfsN5rRV+lqIBgCvmvYiTilqCTYN2czibXAQq+SjqTn+eTivcpDZs
9z20bx31ZncebscUXeq7epUPbn/J/Z4k03/bZkOT1NCOf0y3iI4G78d+5rYsols1
MK0fnBLliLyu1wb5Mfek+qgSdfKn+XZZasrDJigxiyq8SRDM4kD16NyLTRuljWKG
u/DApIOBNoHnsdEZhwMkYJRkgwE7iWrVy+LMaHqB+V5adI+LW/lStpJp1frSjCPq
AY+PNwKL3qCoBI2KxKRgZgmnoZ1/NrhqgdKLsqbxnFUGec2Hly+OXndF3R+BHq7M
c0bwrAQq75bdHwSpiomfeTOk57j45EjHpNggKJ/KDTPrKf8AZ8ZzavsHRD4SP7A8
ye+IgBira76Y5UqJXKSMBQv9sXRqAz0cUcqQ5ZK/pE/KPSmCxR7oi6nlR/gc0zkz
ThMKTdlTQo2wFlhrBiydCnxQnsBE6G8mfYAiz9DH5AQN2VqGg6vVjxzbMuhYRRIK
HDSQIFs5zdQB7r1uq+ka/ULyEFZj3QGBbhmUzkzO0r/6ZWHZu3F4vTZoj4okew2q
VM3B3N8sL8F3VshgiHzIWJOcpRrFCBYZOxmFwMP9uqLno6Bx1VawAMXV7g2Sp+zt
UiH4Sy1lqXhJBmbGr1PvO5AE3m7FSYbbXZwGuunH749D5Z4uB0uMGLKLR4TFow5C
4Qs1HTF+Z6flqETGFoXzkaWuDPw1s118nES9oc3Iak79rVJWSCswK+5MsjLW0NAT
Efi8DUVm/5olS3dXX1rcb8Kg0kEDA+HM0wVZkvhkZhq08ew3UOwx9nH6WPKRwmV8
eUi0veIE0JwA3Xdj5fmQyYKm9yhxgSzOJiJL1kytQjoS/qhSPGKvNtrzpcN1AIUu
mVfemjT4sLjrUH70vQeoVduu9cGr2ZOGwWLb3nj1iLzSRW0GwDLlsuy6s+PBRxUw
Nd6snonsmbVarzhy6XVOCU5YYoJIQwGEJYKgk4TD6A0OR8Pad59hChrawP+Fz+il
XlENLNXLGjnWXTwhE7a2MLTZ9ZA8KKev705bA7+g3GR+5NA8xx5ry72o9GpceCLV
avLz83kxFJFPnCrMgJIEu3tirjZO4C1h3FVbITsH33yJhDoBsFOSFJV2Z75gnB4+
ejX20he+QaPffMslDEmHrDKG7hWHTjsS13J4fEgjSi5eGM4iVfUpd2HxF2s+voEc
3mzjqS/Kl5jWbvIlMe3eR78mmAxsA38AooiDSuxBDwW21t08c7BtBqGDp9++Z4r2
fPmfBxxRTEBDBs51vzBvWgCniVDp380lkyI0xfx1xg+DbzJ6/RpO/taJlcz3pgA0
+UZQciLqejUXkZW74QKUtaciTXRz1THgAloWRVcdVoHtrGYyj3jwt4xLe+7hPs/3
f4zeV7ixrrhfmlPwdDEL1Nrpe1IhAsknlQ6yrM0vG9nkDTPESTVRqk7M+xTQbvyW
9wed27PMDZXBXb18oJCciOXepk7UkXiDWuQxaeQSDgDXYhSXtiUEQjZyX9RXFaok
ipkwZjDARDqJ9KleIkScQ2t2Grn6XYwHYslRRwITouVRqvmh459LilSrBK3Jd5JS
qPQOOae5cECWJkp+QQy3QTrEZnULUCKM5FFKtQZAKafOFONPpmZIw7oU73qiDK82
u2ZBDqcSiOEX7VH6vHT+AXR4uwJ08K9Qe2oFupilGzN4d4OZesLIqOcVtjxi/nif
RDx4gZpb9yjNtlgmCe2EbPIcePbKjW4M+hxGbguaHEH5lYJGY2pjW2fhk7g7VaL2
mbUjDwfTBkm1TTg5cGbJYYk6A94Lja81/ke1+AioGmGYuNB5cUvjKlkho1vbU8UO
UkrCwUMiIPAWyrzFuezlkFTGiIl6tH93+4BV5iscMUXNQynXfUf0CdDbAmf+fFu/
oc5AK2IZW2SLeDFPye0svhOCWYCapf0nL552uDUm//OpAUufPolBctzlZJdPlBdt
CupxhmkK+uUDzUzCUKuVUpnv23XAJkjUAOqZ5AVdn4xqaoiy+4wVARVagQAjEO2L
RfeyeqbOlTuRqAnn1TwVOl9MNFG6+O+ztayd1CS6MvFR+OU5mFXzRJsa0FkJ/vkX
FD3Z8psRlL1HHqvtjfOF5YCdJcaFBDJzNJxwuF1uqodIFzkTVCBsOUvym5K+aI6w
07HxlvlY+FlKHlD1+ndrCLjxhyohN0+VrhLba08JKtmzXjuYt5W3QM5JeEcikp1I
aCiAc/yl7t5CKcdTnSkWu2Cx/cfWKTYo4A7BNlhHvnrH/mH/5Nyf5vFz2ZSK+s5V
1joajPzOUXfYCKySt5bYlfruawnPwKz18TRTFTx0jY7nqIixhhHJQ3A6/11X5Fm0
kh2j3erKrNU+w+/mhtNwKhEwtUI+PQtc64E2RUpSN1qj6Ypm6Bh8+bNDeJbj+BPZ
WaEcYgoGX9fZx6V5ermx4pSRXnWSDaUwMYAauXZbwf5QgpDxasRu+2j9lK3X4gNo
diiS9yFVQ5A64FSuiFUdcc2Q8PxcgfNfVgv/v0pDkhuG4dWm5nUD4gxMcLMzmflR
oKlH18aKXXwMk4QKZoIHU7tED09YJ+YzeHuqAZAfVOvm+qLmK9H0big6iRlPqKMh
gZYm8Kt/AoPgXz+rTrQSBT6arGWfYzDM+Iewjh5ZQWsCUcZmxqn6kYISQFUX9feI
I7gyoFVYgxt/CuJaX+ZuJHHVRzrPn628gNGy2QL3qYfP5wQ/LP0epiqe2yTPcoCm
Inc2NV25NdAgO8CdjbL6RebZewK3IcuSdV3+cUu9S+p4Y2P7iDolipC1nCpwkKGE
/OO8zNRj3rQqWLkaP31SHkmhhOI8QHHke6FP5CZPD7A3IbCLVmThf/16JLJrRojj
VBa+dl0jlLN9Fnpd4kZ9ffeRyag9QNtkmFQlv26ZcV3PtuVshx3/5uFCwx7bIvBk
tXYvXLe1glu050nXvxmzh9DdsXmsWY2x8ZvmkRoVbl8T9sH6WJa76fcqCi4MlKD7
ZaO7xhW4dtPjZz9I4pRkBZb2ah+KMwHws+nygcAjgW2qRZNCCynRS3cDL4Ric1iW
o0EDGjTitCjCFf/baKL3CtAIC3D4s8DMNCetWpr6Vg7+kERPesC050OtpAl09W+M
MWrmd/IXMfclBdjgHFx5PtLN7gx/qCATE1brJcQ16WBN5dEEUjeAxHZywWTSpDld
ya0PSZtYWpiZhzguuWyx8EjJQa43tX/XZ0DcKGzVHh7C+s0a3VzmY2wzN/XbQi+s
M3Nk+7H49T9E5Sxq0cOeBFn4TGfI65hCpVjzDoEiU/sUp0cEEXKuYmPQGmQX3Bnq
7NDXVwBQTmrQMBYer45pFslT12xRTzwkQpC0fRX7edBqQ2LZP5jf1bgnbVqVrl6m
LvOkpTIxA89C4Z36upnjqmi6c/CSHfI/ODUpSMM3EUU3SNle8SmmYzgoQYnNylXQ
/NgiUWMvFLTvhEyadWQMJ+Tlk62CRDIGwtXYfx2s6is2hKvxFVes5ZmJ/yPhd7Yz
vTNj5WY/kT/UOWHL+H8q0UnebzDLc1b8Ib8HADqe9av1OoLSmlVSRP6oWNB60OMI
NTpC38iLVosXOoVp57LhvoaVo/UxsCMo0huWi6rx/GyTz50Svpne2eC9y/tq8xWD
iiJmHuPR1cJPU+FCAg7wpUVyVFGO6h383xzlsdikagcV+JrMugpC92U/DWPbIdQ7
mV45Jf+SC9O9FR7ACaeEL8cIXW2vfjzGVKuVMpl6XQYBcgP+77seuya6Lldv3pIB
HLLdB5OmnEYo2JKIcYJHZFLW0R0BMxQ8LepAGMfWo2YtUQAavPhgj+nAnpZ+4HQx
C8QyosIBtKcOsb/8CLMxfFaKWpbgvvfDsj0TR7CCbNLghr5XzcwyPtqB7MgCyMhh
0UQV9oVe47W5rwXpQpW6IQLkUJsyR8ZMN9aKx+W77afT585KlX/dluMYt4/drgoR
DXvuwaLzGSbhB+wQUV4zSoCO/BwZ7w8J5TDcq/RzF12DcrY+I4dVAjA+w7Rog/sL
STzVaKB7KakGvfVlatSctYgaSbLrshR57uM+Z1t0SP4D2pnz99xO39OOmMgu9BUb
47dBOrpqawES9JeqBd0GKO4fbQTsJlZk8Magb+oVEmHY3H8vmzHd/0cJn3wE/EHb
bEzk6oEZ8X32fLBCVjxp+YM0Q0C1mjus+RmPcBRY18Y1lzzlyccda/gXRmvZUeRj
8np9bO0PIs6kG0x9zQFLne9B8IWo+QBt2sTe91dxLNZ0beY8JzpNXOuhdKmXDI2/
/yyJn9KU2pKKgNNLZF42AHhyhHhMaVUX2p1OcA7BioL607n1a1mjallETf3tRwhb
RMgVDhyRybEoYE3FQlr2rKXnmW6Uhw1EtVwt3UL8ZToK212MKAzw8Kc4M5CysVrM
dzCfiA+pCBPtrv5ZkBHvU81tFEHLCrYV5uaJ6yzlVOwfnx8qXCOwkqv7HDLSImsH
RzYCuvW8SYcgZO9oacmhjPfULxasGpsHiMfPXO/KPCi1BarauAcFv3hu0R4uDDvW
pSqeeT5SoVRd6eRIoxPLpnA594T+0lk8FcCTLmiwfP+W7WJ1M9PpWBMJqGBA6xkQ
9N5c+t6Cilx2YjXshpG9ecCq+ZsNcGPGzK6S9cSWHG/taRvhkLzdhT0wgyUanyly
PC9T116wTmRvioVUdIi10kT2/tCah0DeCH0NSski0UZmC850SlplVx/NcIbXoJUx
RdmrRx7kwPELcd8yn8xidfVQhX+jr9eyBOQ4jHnab5LCBIRLIBxhxMbUhVHMI/0J
BzBhcjhtlMPn9HDfqHsmtSi0AKzgvLks4E+Wn0cvHBS0ln1jfh1lXPAUtFAmmHiV
P1OlGlLsxYLxOioTAZGSwlzx6L5W9EgSGxNRXlDSCa4MHPa8C9Xw93AIr7g0fTTN
fFFQr7cOm7ZDE1iF8mo0+0l44QU6P5N5SZRK0FbnUoh9YVV20lqoZBT0mNmHd9V8
/XYpxIdEuQII4aMU/qUs/erWhx4sj4GDWNC8BlQc1tGesW+rOeWG0eVXPnSgHMkY
Tz0vVZ8W8m+1zF8GtOHkXZ90csfoF30Z550H9ZNKctNmlzK5zwa18+24gVUrqTOK
PjzL5MCf1uBehbpgWMSdkxt2MbN3JgDNBomXM2FJn1NwFKVQHwM4PQUKSqGXcrN0
NaTdbtY3yf5RQUJyCee3EL+3fsbaH0uo4NB4ZmfUjJkoDBVl5WkykR74d/xNVGq2
PHyRaLH8DEJKBFqmcFIw0AtYeABAaNXmzTXvNw+1hmo6nXmOJVKLcaboEyhbeIDW
tzdeYqMKO35VooDir+9tBs7M2T8q4Biwrw1Plku2BZRTMw31kIBpbO2XAFwaZV/G
0zkcAbWxsApngMdExWGVJsuRMnfNsXnwDIP2zbyHglDtf5u09AwhMiFV4sZnjlnX
NrXnfFNHMXAlLQJ57OSU+GVomGgNSHQVNWinQ0jTG9r2nYC+WXmo6Gv20F6u6CdB
IzerUcJm+eDMZei4IqUca+/wvVyLF5A+Jbk/GMalwtIU1l2UuqPP4NaMK+KSMx80
bbbHtGMBZaqOLiVwkEwE0q/bkItwz0qugn2jxAPMoaZISe2STren24+QkmtEyLLM
5m/GKwVrtCF9ZM+6qxOelFwz5JAkhHgGAci4uWHTtheZZmosLOyswcD0esBa/QGx
Zo5WKZNaaHlyNSXr42FWaHgXAHY3TSQ1h/tkCIIKO2AKAh7UDbAyGNkpXTBeHvdw
jq0Dpt8Ayd/XPa3Y3ocnPkXp1+FeG6YtfFg9qpqoJa2koRmZWSOJGw/4d79U6+Mx
IntTd62oug/C9rOld4QWc19eZUy6Qjd0V1jZyPozyRDy8bwJ+mM78KrBQcvI94Xs
GK8Af6jBlV/jgWvQq2O9IESeL6ucFUHCeGk8ffCPHizVRoOU3ZZkbgR/xqURhJBF
VJ/nKJFOmRrc6hMmajt0G5jpzbaNCC5f5K67Sj+kmi78FwXddWD1MsYSmQfCzu0l
qxUKkjdItfhF188u6fRrVH2bLO3BlGOsPAH5hG5+zgGh6v6q/eW2BOHAs0WmiWv0
ZdYTwF6W4QgxYpKBWlEHn9lFZQyajRJqQy/GLNSSGu6fhWgYnKbS6I7TUo4pKoh3
qX2SnQJi3eTHMOInEC5hyDZXnZeoDv7zKyXAwYKgF9sdTFmZ9zc3kvgj/HFKdNdT
F56ChKmAthiI7nkrGft2KAFdhuzstAvM9xV1XAJpPs5EHFZDdydq34+LvYKoUFrE
s9oa+4Dz2DWN1YjP0wB/RjSJ4b42Vo+bb7ag5UR6c+m382e3LuBtbXTdVTw6CX4S
RfX03Cv08355b+y0lfeB5vcdIdmLD13BN5E/xpj82zvup6qo8oZnzfoOdk8wQ0iq
l5dXLbOHskpR6TZV/kf6d2y1R5FOCiQr/ZdUM5VTHT2XBXfG6tWft8AHnDXQvOFx
7hkaumuDlSMM5n0cKPL/rPcrbMCfaRzW0g1HXveJPAZcoLkuTIx71cGY3Zq9iHLD
cEmV/b5DACwdzFXpeV66+Fp1p6KNItmnw2uTvmKwnMhob4nbVnAgs8nK/U9OdxeM
VYsWD81qDTvohDCo9vAwaW1Qu8nWHwL0UM11d7MgDJyEzKZySzY9NhgVUEHmfBlI
VRTbd1ysfilptNjCzQLqugkeQwqN0xD4dfdixFDyYh769rqkDxH3WcNVxuspifEO
c9gSroa1Y7Ekh4/BgMY6Vd50aXHzlndmSTd8Jl9bdJTJfzl2L58x+y3jp4bAaKmo
9TnRbWKyeyQpieiqLnrkM7qQ+AaG7pZ1ZYWkQ+IhlN7GNcXsFscK6/0ArQTf0hk7
267Q8UuwyZ8or3O5GC9zSods9bSGp2ZUiS7nYoeP6kfhFr19OQtjF1Ea90CsyBAv
BDDTGrzQjYNzl7rFqKRZ52FITOPEtTQaUY7qengB50CvrkpAVZ/q6HXUG45wKJII
FAzaOukgHOL9cBT84bRrgucA28OSPL4gRAjUfFgO0h0nF2UJ4iOy/zXs4IQtrZ/I
ppvlD9rXgIdd37bPg4f7NKZdfHMsvRltfuU72q/BBs2Nzn/mOeWZhXAVwyxpFYRT
z2PnI249UQn7shnrbQcE4KrxkzuFYPx5lSNjvj5NGpzqCC4hzW1eFSuYVHgbwLFs
nz/w9WnsiYWmIIfqE9y0eRp2p+pEnO7PamQvbUWqhEshBTEk6B4rAd8gNzfmcK8s
PVLO6QqG/w3Cn35P4dpvFUP6XbJC8R0IVfH6ulu311aiKHiqXwvgAgvKzM9zMp/q
HJf66sIypHXpwcsc5uCSMWOxJHg9rTNKgMx5K2apKaDSTWI8cKCtEAEQSfZQBggp
PXUXUBqSeYyhNCoDAMOF1HexAms4nTlWGYmiL4dYjiFzpjHJfInndutxHEAHqevy
7dASsa1J1WCDxXQojc6m5XjFdxIEGY6yUtNIs12l8HZCGpaIIvnFlWUzh7L+UO0f
aBfVZ8TrHlYAu0SBcuS+/fCGwU8HKSYevVKJOGMml5TZ5VYxbpIlgfFgp9SSvFZ+
ifUNGZ8LRQ1THBIQHLMqpGKxvL8J9ddxq4iYTEpyRa/xemZGPgfQEA72ZplVL6OG
mar3ikrnSKiJKD8daQ+WFQgzaMKVnNsVIOaoSdl1O7wBOjGT8SwWa0q+i+aAVrHd
VoPi9mITbyUNZceqf9hucpA2owFt3j3e73Xm6/w3EPx00fxCDn7A6x/lAEAnFpZ4
yX+QTQ+lGkzV/IuvUPsc0/tbEAMNZjYadetopkKgGYsVfw/LfGJsumdh5UOpSZfk
GzT7gJ0MhBe5XGoAjTWfMIy9AEOhMNiVbEzNSEH/3bplJ7XxfiG4EZBZRTKi/yBf
rAtB48Xx8e42AvWOFJBBp7JtPKIBIQUFd4/GXxJveZKEJKGnFEFOVoIImA5BHUtG
7v1BpIZaWhzSIKj1Pxb7Or/hh25H/GqkOeVEyWfHeyyOTkb6ekcXSDtgF/4DD7uq
mKScjPAMKqPxxVb2aeFn6xhWEtGJA2VL7t5DwUWUmTdHbF7T+oZi/jimP7E11pIS
Z/fBk7ewCGBBoKvnGpBERuk13QqVpavTtvEn2B0vTM3EJTl98ziivZTSsCky/c96
PyLLSm3Y3M2y8N15lQ+MFmNJVCIcq6wRX8KnS81jOewVXNeqN6I9NxdfZP7pw2Xn
T2VacE8vkVJNSx8r1AtIAWYVkROraXKvgb+/5+Z4hSKbAgPTLjqOzLpWxQaR92FR
fTqGBOJ+sBnaeQAqI6FtOopTmmOyxUcc7kvZCysw1Ypk8HTLeOREAaXX5jRAulO2
JM7iYAe3pIo++5uglOSIHTlx4njpM49uCsXf8pcKW/UL8TiCbpso2U7mOqifUtwj
4ZPOcU3+buyDickDmbARA97CPPMEl3HvmfFOF9QDJlbZecLoh10ElfhyQZ0x9uy3
kGawc5eogiTnenEfFloTAuDDv3RfvnlXkHkOtGRw5Im5DeJ7azwm+UxO8BtM/2PH
76REGA8DRST1AqX3qb9ct52Gx7jKioK0wqyJNKJwFFKcf4VZrDLWECKBVagBGTGK
EHPJ0Ig9C5k+ZUdnQXSskqvOVBsJuswbTsJNiKJCouwU/CZ8En13TMjEaf06kihP
r+IJdkfO7Y6pWwlysO+8cPakEjleltkPkG4e69OU92oQgojg4ngOWUlxfw48Xibf
t5qJTNqgqcqbiuUH+ap0xEfa/b9bfomBk/E09mT8zrNNm+cXr8eQGvCnVhTssRku
zFPtbQIkv/juNqlBbuD/ficAG0kDwphk8bGAgM3E0EA4cLTWxoPZEe31AATKd8kF
2H6Vi1IHqtTDOPDWF0DIJA+ZvWEtIEw9LcLMKnjdrKEi9l3dyR0oL9BKqEIL1yCk
JMO81uIP2q4LsZMPNhrfg81jUiHy62UbkfBQAFWHTBOtbsB1TJnLmHc1wCHu3X0l
C35ob2WPvRrup2L5K/xyRRT5vzLmdbqI4DRdBqKnjf7Z+YlSjRlu0/6lnKoV4ztl
UenNX1UXKTMn5yfvmDZKIIDEwy+6rRaqkmTrM4hIs1S2AwWo8/6SWMCI1HnIQcN/
YrpAsSFDk2QPTTb3Dfp7LNp+6k0RMxZH2/7Nt7S80ojlrHuHwEWZG5o2G8mJGHts
OEb7x+4ZG8OVSBge5hlNY1zy7fgfWTSgR7M61sGIRzOZqrUrtukwwVqDN2NMQReV
z1rA4ECQq/ISV5HxEaUSNEWuyL4w+5Np0qPfUB6+Zj9CtN6gg7C2JLDZcUC+wJm5
rBH338VTyi2g769xSZxLVbAxBDQL/IIS+2dA6uhUUgtpqs5hDKCCR5ma8a0EAGr/
GQZ5Kt6wEcpqyXH5P3Pu/PDFdTEGySauA6OYIjWoPXXaf8bozD/pkScjRni3X1jh
LLoZcs4hnh4Ycm+pONaC1N5XwDSkZHnK0gluV+vYqZT9nKS+CnKIWo5f1/KucCT3
KBR72EgK0t+NYbKtGdavS2us21ScD1KnXZqvNRp+EfxCTStlNEh+I/74SojpR1eT
s3wn6TEvtKIVjYp6FMfnviPrNoKPV/8cZ72AsDGfvHh0rPHAhVN1qL4O/Nav9OIr
xnq4oYjkjRpDjqoxfVErAYUEvhpvPTaJZt5G59LjyaZ72E1vq55ovVtIjbCOTXW+
dYjhfkqhelgD7EC9/tpg9uWv7Bpf/PD7Lh/Dc3h/HdmHddVsWCbV7yzfNJq11qrq
SQKmnIT+EaWY5/GHPsGs0vMvLb8/MNuJT+/jTg+DrioYjoVMwbOhY0pEQw/2BRsz
Txe1dZfg95cxnAXha31SBuULKNcmzifUpPE/eO0JSWLUu/f/sVTBfQSUgU6FCW3g
M0j0wf1buFyTYRkdDod5TtjlMnFlEGYPDruTBXVfvQ6zBJtVKP1jwrTw4rBuL0Hu
F/28sctEAK5mK9KcZyoB59PbK6nizXI4NcINwLDLVP9VAbXHdsmrYtvcSpRedVgc
73wmt3EvpAk/fm/pmC2UwhVfLu2nXh5uEgkv6yGdkEWU6kLT5gcmZhmmrQkIGu5e
FjHE5pp8NHuXyWdnq6RDi8YPg/ALUhQu5n1oqNTuPxw1WG5PO0WGC7pG5eMP/3JS
Q/nKtXXDPAscvMl8htIovReOKZmv4ingddrEQGRvk8ek6rRQwV/T7fx3W1GLubgt
HzxCWP5uSyPuW2A8rj7TVsS77LQMUNZ0b2Oz8JSTVwprudOoXT1nY+2V2UxtNL4B
rtmFSiRPkLxi8dg3YQfu1rGtqwxW4NPe0uiz5KvtXVgkouI1aSAua6t9E9/0wMhv
xv9y8Fg5gtq2GG3CMzQp6ZViYeY3sN/0NfhSgMnXTKSb6feY+EeH8tkbMX3JtlUZ
0+gswEtO/GLS1Eoo8yO3R2Jwgj1E1xC/mOamE5x9tucTXBKmzOCUAIIDmt+SBpxo
hytmFauzK/dpm1REBsH6A5FsaosWXPhGNjb5lBKXM6DByq7JNPCuPjjxl8vPmmAQ
QU8v2od0qk5/JKi+KmvUVry8RBkUcgwAQKpJd+zxwewgJNfU7KHm8o2WFpaPM2yd
07s0EG8yi4rOZqx6BhUDlYQNjYYcBcaGbZxcU6TKN7za+2ODs9K9HiZdg3P0d5ol
Bs8AiQIQ0a9pMFlSK3e1+OzCJuPNOg59/u2NH9VqS/fKjAlp8/qm2fm4FEEBcbs+
BfUHRyOA0LNXAxlCoDIA72NRr7Guout5HWKUhySc7VlQ6i89t2v8RHeXEmZDSFjG
qfbNdg37jiErj/jnT0dJyTyOrNdhsgwj1YhMLOeVw4FBDqC878NVRZSmMerTDNRI
ENQUeVA3eV2SSnbdM8DU45WYxsmep7Oijd0Qmjm4gNExKhosiHJfsC8sp7LiiZiX
WIMYDbqARdD1C04ryWCwdYeVNslTEtIaGweUUi7zU20Iox3IymfgCYDxltXbFFVh
25+hV76MFeyLQYKaWifQqNwL05oTh6jU/KPMdzwdvKIZivlvmB9Vr+ATI4g/SDzi
/Fr+deqGOwXyds6ExP6D8tDltVno8fXn1usAv62MJ97If9QSyj++LHHkfK73o7Wd
+PT2QcumjrFi+1id8FuyIgoqz9Qi6zAyzthCs1qX1Dcx2V6l9O5LHvzp9132Ycby
nW/kzMoLrgNzp26+K0LYtEOlMujH1lVsALCX1FynXEh1PJU5WQtJ1WF/HR4qyOI8
ramBlobMU8YfuVdBDcnbbD+9RBaVZcU8KCNlN8/Ezu6ynOnZyaiku9N9sjZCag+u
IYBCirSralIvHnDWd+le0clyjQDbkWPXz0ByIGQfFTNhtZ7lsKGQzR5UN9Ar3pSK
bpMsbIgtdxXlWfAEpDsqqe0bnCQZx/FRQCz8JT7fK7jlH/qSWTDJVXO+L5sU65AZ
NZbpz0xI02VUeqjPUiH/sIHQWgza+L9iYMQG+gu3IlJnVJnZsBXCOJTMJOeKey30
hBBCXFv7lYERl4RKQ+q0SI6oB/uGGG829A0evITYaONUlTEjieSzVPqP158rhsnc
36HychVHLT4btuEr+d/IhSpmMSZdMr1EnxFZrzCO4mKVY/0SiBdnypYc8ocHso3Y
sWiZC/Y6BOy+g76xSFbn+Nm0yC90AFvsA313QYy0l1NIX5Oqm5rjxc5y6upHtdDC
cV7zhGh50zVakLsZ3+xXj7wOb0g5kWHeIZ5bge0FlnBMcUUZowUnv1KdmicEpd+r
ZQp36elLWwEC15TOp2UXmF5P/RfRMOHTGpI5wHx0wl3M15+XSbxUi9U6EqQQ7qWk
bUPWCvkd5/VpXdSg54KNDBd+QF9dbCa6wVM0s66HJi1I6B7kuFUyHrUYeTAGMHVW
bWKXYBlSraxUE6fZ1PUSMkQzQA7XHf86hD6lIRfYPdYii3Jdx+i9xzl60T0hwwhT
I/PDDA2gkiYGQ08FazkLRqhxsOyZ5uBcbbRDV8J5lY7d3x1IJrKEnRtC0SyOZmUJ
N1ToQbS+aZd4YtWRam9wzu2Mk8CG8SmUzEsJ8BgPIYaiE4d4al9q14c2QICKH6Jz
R/Q9/yzZ8AzVb24NGyEmQ/honE6KAVObHP8BqPwEcMqJ+ij6SAIee/GqlDNJdFhR
0yLF2MVitN8erH0sQmqAhUB5mjWdcO1VlCGT2U9Bc6SJFvmpcc8F9MAU9W9U3pbK
N60egtPOOKQtfLprXHnzrlZdx11Bkf7tL6YO14dOQiDs0zmArHtwZNdylx2Na2Ub
DRNl6IllE2HwAXJNyNwdwrpAbXmRAFdGQAyhnTV4AtGWw/t84aBkXfs4Rl7nVE/A
SDV9tyGirHn2NivOHtTmiMVbvaMQHIL7cFLKQs30St4ARqA7cOCdXFeAnQuS1G0B
tZ1XwWA4rnDtPaVcYRs3UmELxdq9Bx9M3tiJHKLzjP1dBbRppeCuKV84gGDmj4Gq
jQethHT4bF4TRShuEWBWYNgBom6el7yPaSIII0jAYDByTpnqTKz7gzjCldT0MVG9
0bqakh1KuvpyUvCU+KvIFu38J57wxcxAcV6rlfAj+WZyyDqZh7k7g42/9f4ZSzfj
6wEmp5cR+DAb6bhTAL9013o6RzoA4Ig6+buis405CVuAZNIPF8e5FiPjflWKERvR
+K+IMa+BUF6Kp3MQ7Och602FUAFFR+0u5evfPQnihELk8d9KVtfsfnl/lyDTDlxX
qvef3ngQcETxV8cubvhG01WT5w1Rfp/AL0gNbZb5wjsS5AR1C8ZKcFWe1MCbpO+a
taM9qu8MUoqpGYvrnqIDW7x9YLznzWUXmEvI4CLlyi9K24p9eDEOIGWAPJeRJQNG
pxiOt6xtHegOIy8UN4P4ocTlLxzD9wNUmNlz8cIlM+88an0P1QKel0A9Lzsb792W
qAkfaPGerXQex7tnJal+wZGz7TRfY+yOwsFSv0Gvq9PTe5hrUrwGuLKUkDdq49sf
IJ6KyBj/jwFbl/qr/x3Er3JgwJOzpEuu9UIu4UkiodbP+Ek8qNvYsJH3K3W0o47V
xZ8br4IeMnmRrFfu//1rgFBJ29Q/wr145JSo8QlP3WNwn8M0N8OQT92eDjBd9Plk
5nWTe5WC3fADhiQNIURv1QoLxOlqEX+8rBzODzOXVnvpyjb1eDthdKl6kWPRVwaV
7d1jy/PZTx8iOhzU53oTeZXPG2bin5ymC5LgMTGuNttpBh/tWaGC/VJXz8wJ8c9r
QHGXbx3LqArj6LErc2kHI3DDHNSlio3BDF8VZHdYvaiHdf0dV/+1M4Eu4BTKJrX1
AnaqXtsJm1KQN/OCILNtj7bEZ34f3PDOQSjrhYF18tGSePc5Vro3hMrphKaNe3W1
BWewJORg82NIjmUh0RSI8PyaxiV7duyXJys5A9PdqSpjm893ilAdpDIny0p6bjhr
S80sARzPskNSa262g+9VidP168fipWXpX3uspyJiOUr0kWEn/mEiPx+H3YpmFvIt
oJnFzfwOewhIHjzn3ghJIyRxFduikpNVb7+yWMJGhhwmuxzaTs7Rx9CbbugL3hUA
RoeODYGUs96I6FMvZMVeQa5sdbdYsRjVwqFWImlXPmnDO6CislVTDI27IZ+H7Qwk
na4fnY2BKrOPw/jsoz5XNcmgA+PcAZ+WwQbdCvwV4buCvsPYZlfLPEDKvvgDKxZ0
P7L2THTP2eUehRV7wK+rAGBEDH47zErVcftjIRXHyjvJolrfhcTRxZ0t/idkCSFb
NJmvq6LnO17AVW96YLkrkw/CnWDcxEG8rDgupRwpR5+0X0CKPZCP67yzO72hm70W
LZdvMbKSIPl2WDfWe7CCFn0fE/HZwtB9haLNqYxfIXdXm1IBQdrzYVHkYz1TAEkm
1FaWhBbTJ3g/KlTxyCvaGy6kGA/7Sv73K5OhkN24jbBOtSryn7sxP8hjZ7nsP1QX
efliVqElvLRPFq9/kSJNtywHSLfaG/xDwWYsQXDKkW40+/D+TcNja8ERO5zHVPnU
9cIRq1JKze8Ss6uChXnS7WfuYFbMaVLEF88ZCoSS1L2IQ4EhgKlOVxjwgbz+ORcB
ELBsSJ0eaMjVbm7amRYB9KfF3VQyx21FOPVL03EB6EMqP3dIjGwdXdeJjExcDop2
5C1UfPkfweX88xwcaCW7SL+1KtPRh5PEzJmIs/cs/2pg8Me6pSubAPQO/PuxtMrT
fYQ4QBsieYwceimw9zHjNbjMDgL9QDhH6vv4oy3YzIJ+c9wBcyN1JXumuOsUbowz
KPkTinypwdDPo8LcqqsVya13iNCB/cVwdl7FU0XmU3gkjaMjBFA4KXCc54TBVUYG
mtHCCm7kHYs5P7XSGvsJByaiaL/Xjca26PEKqBouSGWPf+cCU+pg/XuzEQPa0LTh
smwYyQZu8YPqDIpBh3yrKQLPfnu+WNbWlDewxt1ahF02IRPCZfg4kMHwjeyKDzg9
yhuDpdI5pjdtfh/j+kTYmNnoJJL4cnCHkgbB+9yBMA/0a49g4daxNfwm2DfzfrIE
49uEjZnAnxJr6Q/VlSAy1tDDrtJEDlO2TXfSt72Sd18+SFL6KQxVZ6z6MiQvgDH8
x6GCi2+yFFwRMAmCl1Rm3W1dl3Mq1EXE+78yU36Qa+VQmijPrW39IMbKjLD5pLfN
j6JjidIix/WjWNm7pBHNsESXARUZ+ahwjxWxa5tmtU+Zl9sb+sFVLPEaGWzxrhPi
sWqd3B6GTHI+U4kd1cSOnVLedTe95OSS2oMndgubLSHgaDVyhakYgVmbNBe3XVmM
WmwMMx6SccfIVtGFtvma0zze4SIiot0X8aw2vTPdqB8UHeSMBr64ZxTFBb9o2Ndt
9A19DxGqdnWv9FClUgKUJYveS97oVhQ3lvsotjB14kvRd9R4p76eNMUbeX/UrpwA
S+gm1ozSk0c5+Okata/9+z5V+3VHjxXIVQE1bLVjOzmp8mWf5wVfez6aJHQjX0kr
eXUza0EEBkls79odpQlv+uc9FveWOnz0Vwl1ZBZZfVpxj5lioJwZzrsFItBn8prl
7HzUMcuY5OLNQ1E/wScRNaXmV9ogwMvgBt0Wk37hfvluxl6u0XaSs/P83vlpbQc1
DFT0LuuBsztDL5Ib8Lulc5TeNuTDbREWyG9ceRJmR2rjmrdAhwZ0odsHIQku3xz0
kmyeWQYeI5nSPwjdbP11uK/W2Ox2d8sb+y6eyPk7g+wtRY5LVX15jXfpvuR0l+ku
4ZXU8Pc1YrPZQvSCGkFIx3qNBg+WiopbaJXmsgqHfJMy+I+Xlo/XGy+USWPRQxcY
kaosg848EIJg5MSjUjuZeHICCEhjh5iqHREhPsm0k9y2oZZhR8074AsvHxG/yhR1
GJzDygBrK5AqBwU6jYJ+lrLzV2iT7dUF1LYvc0cvl7ZKcektOpuqBrdFG6lukaUu
zT/4R9VZCgRDbW++z80mdfLALbAOxlZ0/REpPRIME3YVZerhUx61vdYwbfrJN769
/xkdyewlJhG5jwlJFD35rti2B4R2I+BoNxVpKuF8tfp3Q5iaVHVcAVcFq4OsIg2+
c/fZcQ02VDML7X2o2OU2qBd0rJJbGFmJ7yuS8y5YTA6G1t1l2TwvRJqHXTya8aCb
zsNDZljqYRb0zQw1iy+1Tv+8omMCfp81DkPEIiU1KQCFh1XzkTJoaHpbQ23uqKwx
RpHfIQLaVdZLupskqm/NiJgipLCIxkfXbr1DrMkDQUus79KsZ2E2/3B2/VZPY1hY
yzinAdlSNIBAxc6z8ec7HmEmbKuS39hkau0e62oT9XH3CD+vCZoC/GFuaVbomC49
k5D9DPkGwf+r2APRf4NjCwQDRKfM9GzzOzaNcT4d6CRDdM19B2BL0XFr/3LkY3ue
zzNXHsbKqkXEIrjRwRpWEZoDM3sjoxEbDfl3ildysXrTTQFGic+RI3mGnk0akgFK
Vku7JXd9vFsW12NeTnvL4dv+tee2rzkn7lbrY50+CqmXZmJRKnWvQF/uub7hG6At
8qe1hHBCNx/OZIMB/lAre4YtS1ZlGz+/KEy2hwgsmOdrxQoWjQhd+rcicQiEl2pQ
L0fHYF8MlRy6hlVVWt6dzLxBvdTTnb7MRJ/TK31mKazwALddItMFEIRsATjDE/Ar
zRyeT0dL4KR8j6NNOBmPFaajtgy7w5tLcPUzG4kFGARJTryvTowrnCMRfMuDkZxY
xEyki3IaVEmSZ5W1aUhObHNW+cAO2TiFYsJitmOPThp6u24xa/Pq6ApY2tS1okJx
yTVYDQMQ+YBRjPD1+AKex6dpNzW89SQwRlmus2Vuie3LFpqcX9dtDzQAkW64Ur6t
VMZIC+5f/HOk3JY4RGrBGbkhZcdXHBdB38PU9bQ4oiIcVDDEWGB8FTbG1GN6urpw
TRz9MprYJLxWREYVAZ3rU47rKiZtWa909S8Xehs6NtHKFGWBFNSkvcSQmOk3Gvgx
kfXu8dRCCvWKwZ8hezjcI3wiIc1i2WZ0x2IeCsceny8kcVvPPFX9Oi8FQ7R8eXuT
GHZlJpPplhN0o2TGBGe1q2D6fZoE0PD7L/EfpxhtF3/RMzp6MYtwxKcfJZKz+Nts
ZYtQW53ufxQ1ZE8lMPoWYrI5FJg+st0ilQ3q6rUqXqt8QsPSvjRQwM7T8UZHs0LU
WTTN3SFS2POYd0ZmkEZsO2CNmY0CTHPIl/Z/gHjK6ACIBo0OVXxd1szTQVsyhEW5
d0qLJCwB53XzR7+mO0xil7t6cShWhGmNq6gHQHhF2vSm1vQIePTG2+fFBBbyhKeY
JjY2fZptq2IOITDRUFa41HT6ll/CX/M86ZF5tJUDwNJDVnjPMTv1W7rJp654HD+W
3p3wUsOXHWoeWCLasrdfqqSlaHsd6aeKA+ALI/0ydRuhC65FBnVNM4p7P8msjAeH
A3SPHacbkmUS1lQQ1aVK1bmaVWF2e/lH0LHQ8MqXA7oSWCxsS6ODOshQNEclHMh5
UkGUrpX4dQKJPdhuTiiSVyQpMXHk/pt+Pqj07qTQZa0z6BckIzhcfoPlfvf8RK5b
GgSQiPWCC4XTNNVv6s5zD4IimzfejmYskAVWJbstucc07QtApqFDabOszvKJgth3
dOXhfdVAN4dM/cNmv4HI111Z1b6Z/Kjb2JXhMz+TxzE3nGrCU3YuL4HXryKSU5yc
v3p+iTkAyvTeji9k0LsqbbM2hwxGg340e6jKofr2rOC4i7k9HvGMCnI4K9Gil1Oc
tGg23JMFjZgiM964zkcLuBAYDHQU4dg5m9OoOackSUddkDQyPmAewnd86TdWz9D+
f61NoXehz9hmcisaWkYXYC3fw7lDo+03+QvUjUphjaGokErSFN9dYh75svO5KAZY
M+/+3AZirPC1xQOiGI6r/ogl10EmYeRrrB44NYIj37HLdnUml0dInRhk0yQH7Q8t
WWeSD8Y9a6iwy/sgCFDhXCFORMNTjTE736RxwJ1Qw+yN+fdhptskqw/63BJsXcCD
zyeypc83RxOn3OorgNEDT2Ett5Eoh25rGtFUXFxHCLM1SIhrF9kBhDOxDdg+I7zD
EY10nni0fmq/LLEOgz0jfOXFCwp1dAUpdMUeXw2GvGX/sb6j7VHg+XBFC+btdKDE
uVtJn1m6jIrF1xxqEWHMHezWmVwSP38+LPKsdIFv5R460bzl5lBx79OBQBER5EcQ
+zcTIez580NpbPpLhpnFxCWWrhLpqjUenHWn7dLQd9S+WBHqreMt2gkkrWmDGli6
IY+v6fKJshBumyLws/G6d0bGUzJxdgH6M6E8jOwTySp5mlFaP3V1MVX05Bl+BBee
tDUfoVyYM9zDHh3Xt9BkpMgS/VBP3cQ7OPu9carpSRfsMnjDeayA7rMxvBhlyTb7
wvY7JyZChcKGgPz6jGEJ5d+U9S1IM+GZHZbS+FPCsp8sNJRI9sFbYNtUnVJR8UFq
AVhSf5+CzfznTWmOFAfCVawoeHS2jfNNW/heCGPdpgME3xhM6Uime/0aO0PQHPVA
YS8pJK6OPw2/PSCvAVqBtA1ibPigX5keY4TrI/0SXW746l8qZMv6/R5vuRWSE0FE
foBA05DtnLCQHbdskVoZXopH4atWN53QsW2LqiiJkQjfKPr5ygpVosRzMGk+yozI
Fc8WadbUW7PmPsJGzd0+V6g2fQpxsRWL7cYZHSQS/UvnROZJ+uvWHu3ZTc8u3D3k
aCnGk+D9CvUtIXwQPrlmCkhmpoBwY1d0q5ydyQhzR2OBaYNbD8nsW0wl0ItlKPgq
ANIfPY0LaZrTl1MZUC9WvVzspk66NI+AMpk1EGY8wIs/UkG4hGTNIryhJcAkbjTw
fyfQNCbjEyTkLeXtpSQluDhSoz4Q+Bv7Hy/B4gYmN4ap2mhwByC/Hw4ceBJjeTEY
e0HS0WyOapiBRD3ls5YLI4+PWOaZX8z0iX1spvbPssmDqm65ot5IKHJjwqLyJPkR
ChKiLscQzcYqCd23SBMtqnmc8f2js/hOhPtwUN5CNQHwbI0Fj6E/pol9JMrGqJ51
TGVxq2R3yrd0sONkiNwxozLZ7mpnhYXhxGpqXZiHlNQQjpF7Fz7d8trPnaOtUF6e
4HhPHAPkepDDiyGhrlmEhNEeW9iSHLR1Z+Iupflydzo93ps4meN7ZBo2sDmJzVzP
br0/hw6kx/FS+K9/13/eRH1znsx+eSKQtiOTAsvDpSPhBMlOIcmoqPg1dGXkHqKD
gpF0iaLs4wFYn9bGXEnorPwc46rkEjnKdh0OUR7eDtWrKMYAQuJ0FAwOg9FUqrjy
Oin3rnV/5pk+JkUgBEkl1+9uYVT7lkj7fgzoUOCm1EU6zPduAPnqzmk6n4Tjd8OY
oByaAlSd+P3VRh13tIb8OdEHBMLx1qcrc1WP23VEH1U0+MMVtH+gzIkfPziFFLcw
sLs3ZmfJ7KSr19+XSyymGYDO9/yRFs6DFp5OUkPPqd2iYtIrdxY3ZTaW5rXNNrnH
cKoTpVM5u8ZScgvnHwIZYpyDAGKN8RLcQtM3xSxTZ/fhhAUmcdA9Tx9zuyUrc20u
LM2Hg/oMMxIZhMz9Jg3cRvwc9GaANmdo/VM+PPo1vo52Nd/QMkA2cmsTajQFtItI
27HiK/a7BgaoXWaziAKDRVkCwUl+0O6g/JwyQfUHI3QyQc5N5SdyTC7XhtkIiwve
m0oSItqZ7tzbeBfHwBdD6BdX4VBYnLu9xyHUBPYvT6f+zH6/f883M1PSqoytmuDn
qnbXy72ypJ4DSCLopCFD48RgS67HPf1q/e+90+2EagpRL1VktQ0iaIMmxNOPR+j6
hSHZzhNQ2KOAH6ZNZna7NQcRTyvm3crQg+avj/7U5S6xCLFivkynrby7bN9i4cql
2yKHth1NU29bOQUTOxG/afx85erR1VIXF/obNGBAifLPselA6vsPzzQRi1hW/v1d
ap7YhHt6h1hfx4dUBlb4cVNVwhlBBFulLYXnvVvA2den2li/eygUg9A1ioMhroCz
mX0DUaSOtoBJR+t/BF1/7aL13ZczoLV8Bober8O76f1eg90xUKFhuK6QJ//ihoLq
EzPLFVyiYXehp4exmxZ8TB4LVU4Kr/UeGNZMR1E/BXpe5V3FaQx/dTqVBxWp8m0u
607AgE4QlftMFWL5DucSijIOWF9Lc9VErPXBbhdzS0UcOLxgrvH/XSMHMdGcmJ6F
6pEFwmXBeNeAMmOH10LMnzUg8XCpuoQ9mHNlBj3OaZIZAwofz0elzgFJPe8ffeFw
01rEkTH4pNljfA0rSBtQQnfmrJJVET/BKNJHc/9bJlt0CW+L53/tE8t9W72/y6v+
hHGw7JyNXBjtpqAFm9Ntt9KdQPaUX1MJwx4x9p160es3Ndz9Bqp2po31MDGcsrAT
A1s2928dZAf3hgEyk5pTobCH1E6+aB/1Kirbfv4zdjya1RxgBDb8Dj6ggmUVIzZN
BMXuDwsCth2EoIfkyETgFOWDX8HF9YhdBu/Eq8hEqS5o7iChzgyI4FHXOdbND1OA
wo2V7RxyxYePwfUudpuPiTJdV60Cfna/p/n9StL9fYtrLeqpyRGiI6fl0PfKYD0I
LuMJWM2OFkJVHOqCGwbiTU2Psfw8WZ21GyKif4XxQkNd0ZsE9mVWzD6tB50ZP6e4
2T7XQkRsN7QW2p6Pp/0NZIThJJaPO4d4b0Jb0bEoEHEJQE0CBDwpYgKUoVnk/N1q
hxGEwqi/QQfF5CfTsk77IJA3kj0NfRgBwjkdQy9l+QGzjy7iGTHiVeTurPMoWeld
4+rrUvHocJUEoLrYvmxG36sNcmR0wNzH2Hk6/Hxpq0nxBlYPgzLFL9ZBPAawF+RD
Fc69tICQOdRZuxxnPIFbwxHDkVNCKZNg4uKdg8lXfX9lHGpPv0JbMyMgRK0Fca6z
u9COYwvAxOHLtsZqQf1KjXyhXAt1yMDp8xlkUWTKcmdmqkEfTwcgWPBI3h7piTAo
ca7KydXDKQMc4mW42XNQt1UHtaSM10bPS7Butz07blUlJXmhaemfZT9x+yn7CiuV
9NiQY7GHwM/b2nebzXAXSrKY0lLPzuFfkrTpgHFzTgQD9jeRZVf7zPDYE7u7RlLW
bseQdjYTbmncNg+CL4VbdROKMomQox7IlbLQ/gTgANoALNepzy/46WZyZRdhrI0Q
okijKoFnkl7EaaoCbl1XyjZEoObgq5Q9YSr6UctH/kpw1yzbhADohoLlLubxipP/
S+NkTb4u+PM7SiYn2o0Whx6B+JbUld8YGUozbYjuO0JMIU24q4yQOv2sdd9lHc62
VAk9VciaOFj+HjcHDgpD15C93Zw4WOKt8x2Gc5xS+FVtpxxJNOXJR3or13Ksb6Sn
SdHeUpSS9rURQrQ4lrOM5E5KMA8VzewD73/dpUUL07Ovip1ligHnyfkqWlsp4CjR
dH8E64WKmZEQ2pqPyBLBwRwj9jVGaIvT7laER60hSL2pxJYIWbgZaXP8zFHQfsIs
3njvddOb93BDJ4M0dH8AAxIs0G66WzLafwETahdJBfjwTmkIc3MAmIxjT50JZa3H
1SxQMMz2x4jvL/8Mg69uAo2YJeHtw4XrrGSq+8vPwuMrrsSwArhtHz+tAgjJoHQq
wr0A9WISu1B84ZEvkzOmN6/LgoSCxgHuV8MfWv/uq5cK1Bwek2WSFjT3d1OZMS8X
ZCv6c5v+rVTvbLz9lzAMUCmHzE1px+P1L45l5ylmNpeJbEvyc65QbtNNJkHfxQg8
2mIFXBSCw15UfQN/LafES3xYwZdlgEw8ZdTdCdUHzUG9w1aPkU5TgBG1ngXmgRPW
8MVKRkTOYmhT+zr157qstqAcau2nuPrOQVARbQ0Jpzy9MRJoez0SULus883UaMDp
jQXfmRoXiFPfvQkVt/m+VussaVc1w8pVqOCvXto82nlssigfmSPS3DlciSkfPOBT
1VQZA2CSye1aIFxa84GbPy7GfrIjXJMySIBVNrBWQgYWkAaJc0R3QUpTjvq21Cbv
fBpK12zUnABjPi2PGvgtYnE25HqhKGLhGiqcarCaerqZ2qbJ2irshBska1PFnEH3
O4zmPHtKND5753/nSPqm9O2XZONr9Mb8tOXrdSjzDVo031s6Rq+JkbBgsc0ygIK/
NZylGokx9C3QwZLZ2mtkXZWSE38kAZYjQTGC0FAEo27LZxmnjgl36YCVyQJLTnS3
ZsvVcCboT8hJREUdaA0gfWGLJafS5dXsPGJsWMQ455NMUl1kmtebx6iU3pfQCUwk
W1RfZqTTdlvR6tTwB7W3d8lCbsUIWRibC5LVZLtXEta+DCFzYEeJcb1jWAzJoqBa
NUvVgWCVkFkeExZGlaguGhQ058kMJ0zqVXRKoN/9zwMLdE8F+AteISWC0LYASanx
jwIAfsWk0/21toMgXxxwDedr9xr6tIOq9lfklXwMc4zobOr6RwGF9TwkEXNr2g1o
lSeIteb4UUeD2PXguQQvDVance+TgqnvUkDTN40qHRt6WdqhUqBgxaeOk3EGi7Bx
OSe10vuuFZl7ziJ71mHK5Gd7N9s1KUw7KMGqjdJrTzeRy07oE0FBKjcJvTrxf/Xx
MQ8IQOxH79uBcmBqiQqXpqMZuRk7PFhvlFY2VWFQ7SKIB3CJ+QuAVAFcVdoYnM9q
T3d26yexA+L1MpK4VMtPOYRsjIhQp1uWW7DTTlKi/9fdIJXzEiNKFAjAcvh0DgHu
4mW7FBsIzNvGA5cCK2AlgOwaRm4mBOYW/viDKoah8kH79w79o4FXANQDcLN6Hw9i
W6RqllRfhNfj7kZnO58FKgW3UzMhQdFReEhcRl5wONajvDs1UDrCHx1wfzxqshK/
X9qwE3sXq7Gh2MKBT3kuRgAqnajXVWu6g3zsTrp70AHqw4BvqcYuGTbw5zHVRbF7
y5idvPX+ONuRfZHszBo0CPr/s+SrDZgkLrjCYgMxuc4+eoYcyPPubqdi6WvxAzdF
QBRtLVoImJx/3gfMqK1xQgAn5ZxZgqK0/NN+EEG0JlJsFVcRXvaxqvnDsF+vyTxS
lcDgc+9h2AuCPSOaRTeEMCG0ihJaNEwAaihwr2QAJi7BZfeTTO0yTlSns8PNTbQI
XwWnXBl+edVsDePpxwfFjWGZLSMNnuGWo+W/tmhSfOS6Et+3g0QZMvooRmBwUv1X
WI5ntMw91MIo/tfwbkc0chtuN/1qpT/yqP94uoGI8HeON0heJoUL3rT7gBtQo8Lz
gPMolBh3F5iAYnwhEuUCMhv0hTrxLKKANkPZPghe/kCEwdFFc7V1pwmHX+dHAOtM
mUca12dvoUAUPOKsu3jqBayaaWKCtbcjKfxQSHRd1kopXxaRPg7lhGGQJqff4ylg
CrAk5R96nO5SJIFtLKvyo+eSNBCjFYcEU/GVx3ONS3CPu3UN4WQioSvAQQytHQqs
BxiJ8YRrtOPCV4DPc3H/JBhccqkmJ+CHpeix2zUYLVrGFPVmxue9T8Sw9r9YsBdP
bE6IJ2hmaGXweYRlByXCSTPhdU3iFPII+QcxUqFWF4vmWnTTlIdBsbSqrPHPjF8f
39ny/tAoRTJQUt6Qm+zqwDq8s9v21s/qPcvgBfQ+UD3oMhFYtbNRq/wOr4491Q/g
qrHSN5woGv2BMDwfk4osMrjdoZvocoQKln9J3zxFh0H3NXklx218dyoNjj3VC4o+
E84b8x5PlsYhZ3MklzjDLXyJhzFO81yi1CrWU7rI5A7dT+kLuqvMLRNRiLzTdBgc
T0gZkaduc+jwURkrBqQcvd2Ep/fE27iqmRoEYpINBAjQSIkms5Iht3tPkSBSME+v
yUAlR87SLV5zJ2+ziXVm2eIwAI8mY8KmYTKWV8MmeFbFLqW/EYctS/z35fi5srbp
+XLZnx+v6yS+WBmFPpVIjwfP0N5nngubcmy9viJSHOQW2T8NR/1KObDy9xe8u9La
0ZgU2wwt/yLlNfFp+GoBqAyKyygzGAWrMD47W64jh8W1jcUfvUBhP1z23+Lp2ivM
1WrJgHAf2LOAiGXwVSRCidJtFvJ8fzPHTrpdBiT97Cd9bDhKmysZR0miC8zthc9u
SktCaGMHiPWfzO22PyiQ5agWLFw1YyEQ8PwvLewF4dp+ME06BRE0KpsG4tl5Z790
Uq6Vcs69RXg5grfaVqpR3lZB3jcH4nMxlgxrG/sWP8lA7280mT67YBxand/TlrsV
flYBgWXLJ6yLnIcQvObVhg4HY+gcNEY9hNxi3dV3gZLb5YQpCUiIR0+vn39SCNXY
i7P5FUvqCCj4ErOPrCbSWDTCvzWKfSVdCY96LiaaPlkdsRI6cGLURAcEhmukKPXp
yEGVPONOUfB+jF/JfVJKbCVpP6i0TH9T83ttSSHHeZdUUdelcbDmz4mCAV4JHa8+
Xq8bIBcUYUwultxgEO7BXw4byUSr4qbM1BNGFTY4buPJFHKundTaoxVv6jBNkSlN
Q/NfeuZahcNEnNCPbHa17omIf+r5Y/QQp/T9S3HbKFWye4m9SZQnUFO92dCUp+32
vNxnPdDSfB1Sn3NChSlR+3pTIzgDtK+hZFwCN8gbWFKOagtLmnxeKDqryipoqpkq
eY6+0lNglXhqoVByZLclQCAC2PW349ndB8xVT2MOKmYxGlvnCQfY6AAHCydGTxn8
xFzoV6CtU6XgpagqBW3sAuYaX9xBvsIgWk2rW0JDayMhFZo3L+EkXrVAGjdGaObh
bWj+8qAIICFXk5oDA+yNRV4KFrAqp+k4sj2CkKBjg4g6thcoN43NbKgseaKdPS6Q
BRz0quG36zGmy/Hw+d/5WtzijWuGhrIZLk6d5J1A2O8Pp/2iq50YbTPMdvMrhSMS
3ndcpPAd/4XLm+4K+NAOAwlSC0jpvmyyCZ7BCt9hTm6ORanX02c761oiVcyiUiJR
8Nd5nZCY02y0gG/71wd6OQjnsoM0DpBQRthaEI9lfLQ/c28+TFBctjycyMr5udOP
WhJ4Qjlm+yNem0+CwY+nUrROBu0K+6fT6xuwPIwrhM3jmArJWrSfVP0q0MqlUdV4
UsM4sT8B9lHXA4S/UT6V2NuOvOfKkL3vo3IYDBilLqMl2GY1B1Dxd4I5tC3gF5vp
zRYP7VWwCELBNOfQP8R+NaPiRM+MupD8bvu4JEEi0zmSds6Ey84gucREHHhFiovl
f5baUdtNglnrTjHsHsojEHDhP8jiUFHD3A+8uQsrMxKozOH2MWHj2y9fY+oq3Nif
O2GAgboKKmUqPFc8pFOtDfdeVzyVifJYPB7Sy3bdBjYyR01/fBHCMzLXMHelzCyq
h4hYQF9RfrRFExPjMo97xD8P7Wfgif1caZbzPPMHnVhnPjJj+0EFdJL5Ib8VKS87
JwHoDKZT6T5hxsheKBH5fO8Bhe4JrLKlGTHwj38qqLTFyo3quWQ5b7dYf7BTXknv
a2zhEQpEjeGMOYfn7fssIJ5CXG+GWmflk3yD6tNnNrvswlXZ4J2Xxbat3Dsv5ny9
U5DpqYNiJ0lzQdLPmj2cu1c9+p8ht+JFiuZC1P4rybsTTUYS83HR8uwxATygFYeU
s9mB1FW+wmNX6vGvL9ozCp2MWTtq07pIEAMLNB0D5n5mjjmoHszgs8iiYy2lkpCq
4msj5TK5Q2Ey9e1OBD7hxlbkbBK48IHlt0Xn5Y8WAhZIJGpvDb8oh8oEi3lKL3YD
no1x3roh45NvxyLicSgwK+Ckt1C1YxssEgOYjFXK8yQKy1bwyV8/Cnk7Z30YWG3c
pcWmzY0TcZlaeu0cLgWclGUZh2nDTWPR/qT7i77uxUEHQHP7HMNJZZbsYZNHtskh
CmTRTjZpdz58EM90eIy9WJvzIhk7h6p7mEURch1bPfdneLFXkYFK69LhHgpu7bwY
7uOT6eDZ21E1nh3wiVKJxcfVxAvRekXmR2Xp+qnmTQzrOpjcPk9k5TFE2MxDHjEU
JnQSz2fyHbRiZ7vqr7tg0bkSlVuCc0XYyZPqGHOZA6ZXAlGVvsiE2cJQQ1V4CYX5
FI4srnkKSVlFPtyBcG38x38cn2miiclwoMeDhWahFL5MilEqKOFbU30THGuB+nJX
N/5mWbBx0snIBAF9Xmg0QwBQwvcFs3fRpqHrat7M4d8HTtP5TlkdjCbqMq0qLBIg
n/sOaaEdZLlCpyC0Kf+BJ55udcFA9UnbItmew7qObBB1729jEHnuDmsTSExUz669
O0DQ+FNTR+TKPOrIR+ibd+zGlAsziKax7E6PEUGK0+JYXv+tagwHXRTdK69xUIJR
asmOKUrfmgB2V/nRJ9E3DDAUQa5zRGiKPmf2z+cWbFpt52nOduAWPH9fmBa+3uk5
zrJwTXXFl4L6KH7BurNEZ+sr6My/48VZIP+43vzXCAc3QK93NA3q6lRC5O2PEolP
4sNwQDqhb05TLyNW3ssziXe+Dy1IxP7l4nICKWNhjMn7giSzcTcsK+yr6AxRZeiK
sGoaQOtVecwMhjhkiTpk1eEWrrDav26r2fU6U91A6neaApgcEM2hhjXV8CN7iX96
YmyyPK0/K3YtO6Noya0wYDVg8Aj3u2WCPGF4Kt3RqTIDK01iz9pwHSaVjzF8+obF
Src2AW7Kwco954ZO856PU//dYmH5vTVmGoek7pzBFnucCJBqcl103hIkUI78xQaM
90utpKrrf0k0mQoUzya4RX4xrJ3dlGtLj3CJYHmNZW7cP97UdsXd1nasX89BQDJl
FJSgAfU5v09j+3qo9bT9Qbl4t/X54TPEtJrkwRfgLil1yCO3YKdvdOeXFiY1Tctv
d1N4+9Ic9be8yt7QkyDbdiAtA5bFJX8oJsDe9iDEm7vShlOCAWcGbZF6m3ESbgYl
c1CWCkOLdKCYQYGEhWJczCAbaUgpVfRnJNJKPhOyaSdKBznCsFDftLZG8GCmUKRB
vYadEX25qor8XggjFk6y/9BJ7YgI4DUHDxKPrlnj8TZ0XlZfxJwKp/yO7TrZYprl
ZTIpq1OODSA0A/Z/m9QBgbAAzw9nfjDd3Kh5PAnBOTPNiXx0dIudgj5apkZVCTS6
ITWuyAR/CSQUEQvywr0U3beS5JJtQD46YdF4RoQpYwpU40+9hVKBxI1MqN6yIuN7
oxU/tvatH28Pz1iZJKDzctiy2HZ1luYIbUsionLYGG5wQO6EGGSQc4m/Mv5aqCl/
Sslqs3bAHn/nvl6N4+quvCyUIgaI32iNMIpCDqakOaRz4PETWJHcy+cWuUgCrzzi
gFsfTlCmGyfhKnSufNzoXOrwmyDtwhztGpiogPnS/Nw3YkAv16JKZAR7PXRCvjo9
GzZnSsIca05N37K8M6HhVkwGZyuYO8xVRUltUJU11JSQo+gM7nUZ43OyzGn/WhkT
fvZnEd7+k1AF+55zMTYEln7tf4Z7Kdu9luS+DryJvDLCK2tuLm7js1tmBqYEUpsx
xN3+OpGaGUx1y+yIUPI7USIi4QiXyKeM2wUX838Z/79bijHnSLWP87wjFb6yZ9yO
li9PJajk5VhVD1U4/vt9AI5CFwiJOmDL4+dz5OvKFPCTgUpXAkVjA6aBTIoVAJDk
cukSZxTDcN5znFYhthBydO2YWZsz/WcSvs6rIuGt9AC0AX5gL1RlCuSIfx9Ez/Rg
AaI5yijrujbPM1Uvf5eENPKUIVj332FgvdbjtM0JH3kjS78gH8fZZoP4P1MgPy0b
SjFEyc0Z412dNucnXrvjfpBBs3e78jYivsJVMTtLc4y5tWzQrf40P6ZdEqVqXyOp
3g58M+HcXSPWcyYgzPsXANS6MUSF1O+ZQxb3tV3yoWWef2vc5NRpDUtFUc73jdp7
MxZEhoPRXuQcVsVCD2W0ugjzHoEOxhQWo8em11GrHJ6tNcKqSAWeEBim8JADXaWG
8HUrttfT/H9ARkjki6TZjY/WbmgjsStPorWFQFS+IbwPvstf2puXKvE7ojlvw7EK
po4NTMXYTsCqcE6Q0Gh4qgFdO47ovenEfqiJMCE9OgEtBv531vKXQ3XGh626lv6n
nPOFLdsnpOByqLOr8uKhgg6uleJm2Pn7yEzfFimImQKbNOCGtQcUG56bqz6qPuud
FkDe294AzdF7Ldo4mtDFbBfQVoFt5pNmwEiNXVYB125lx3Lz4VdUkxP8bd+UedsV
0SQ1qG0WQqAS3GVgp7Wng/0pE5g5OuwPlLgT22f7kUqipOUqEqAJWfZcAg8U8X0b
+ZvMcaQ6X42fKaH9CYgMq0+4/wYUqStFPwM+ToI4JDiZrkEx+kYaTzuXYA9Br5zP
TdEylcigaQUk4rIOJV3XkXNKRlQnQ7fHqUGEQ+4LHiD1EiL026dsHhsbN/C0tPTe
2On7H05t4kYM1HtrPkEGZpVfFZknWr5FK/g03lIZqJlEi3ZK3kj0fHdOZ1YDiCFR
UfQlwGKLK2KdJiXPcMLI+6KyvInzUbGe6OemQecI2kFMFl7wky5oXI+WVDiOulQX
AA9zclju8M+ZLwVRP35gc+WoO0/9W7u9NsPf8JQgzNNSzvRH8PPdh2Q+Dz4aNzhO
m+UjvsVF5UirblEbJpjLwNvFd/K3V1knRmf+ZD3wXBPPL/fe4i2LMYah+DY/LxNj
AdHVceV15C/0b9Ulh13k3OjpBlc3PdhDqMMN/V3i81piYib4lpgMwjEQCVDhVytY
V8PIZHNuiPnvBeldmdc3nySAAioXDyyO/H1Y2rVXPhinQW1Ok2vaqURL0Rg6Fwic
9g54/ExOZMicuWEOYfydozQR3cp14xeZoRf3F65XzNY8zzA1rODLJDdrImLDIO4x
sFu9fcIs0heQA91QzssOx8jMKFM0uYnXsCS0UJLrfJptFSGdF/eWqnJOy7UeuqIX
2bmOHG18AZNcRla7giUInB9lWBAYHk/AMP3nopHO5aRUJOjoi8JWxubKfm1mawG5
gFfdydR9FvkCCMg80CZzMZKQemtaIWa7mpTABG7Uz2aP/cbEME+YaThujZfeVb/i
Wey1Mm3bmULSuqvPQ9629dQalvqavmO7LOjsWO4zWfNoyIypnPGcgwKxAsrxzAgB
iD8tiLLqi/NhTb+7t75dM/dccbcLXbG7Cect8MSKlcyA5rQ/0QK6RsEehGvESoGU
+glsSAnWMv/XB7ykbPvZyfws+EBwPiuC0hopziV2q8eYxYfjNUoqJs0FjYlaQN88
EXJigbe2LoRts+BQuxqH/QLYOBmUQgx+erRLyoSKaWWSQsSYDzc+EKc886mqbp2Z
cx1a+9GW70EWXlUC3yitTuj3vXnAkBHXb49QwuZ72JWCEwhDwgdfKE/fI9NUps0K
RgxydYYADmAH6XeXkxHBeaDs6uBSb6cGobCoylG/01wLpmlPc4A4D9u84wZXyMeN
cT4nD0vbL6mk5FT6tQQ0ZdzrjUR9Tgr8fTn8imf0dZ3/vTc4c4sfjm7PemRpIn9T
YSSkT9EEj+BkTdDnkYP3zpYxC46Rn42KOVgkWVPWx4CGCDa/ZB+AXgLltasSUbGn
mKiCWeNa/vRhWI1z20vZGyMXRYanzHIoJybHm/EKeWrn1CXGDvGww7qmjvRGMv4i
h2Rd6vSynoIN0OMYVfz7AU3gR/yDhQRnw/Qw9j/WmM+njPBYMm3zuTHqAPuhEEbp
7C3FsyaFu7pzFPq8hNCg6hX29sIpyc8f3HYc1mx/SzcYCRkCuHM6wTigWKQu/WWF
s6rugcYJG2i7XTv0nEoADC8MXwFHk629gGH6bep1Eg03r98xpoTM3Pps+Vkfba5s
HNF8t2WFUJqmetGGwVxOq+u4iZSx4k5S/gwUBKpFsorhH/Ybba2GLA9JDrCx4x1E
rLD8iP5QrNmUWmurwYaEoX0crcpplOGfynDAJwZLH3TMQsyOTun7uovsHw+Y01ic
2eA8QOdX2ZVFhSJE9xtbhFvQBPrWoEwPDtA9Ac9obmI4k9VTBlFWnOae/g+71QI8
ncIwbucO9We39GlSMaWrCAhgEM9uzAq3aawswoaNUupZ61BiM75gxM/4aGYRIG0B
fEBBEuNa3Fzl3uI2E1lBHdvkipAA6TTFh9eDV5YqV5KFBrSyE9B7wlNj65euYo3K
RjBWifYbCZMm2xcuDnqpjlkNrKwCd09MtdJ5rhbQkSZTVZ9hTTlr/AQqY8cbDhLK
+PrXdjtp43Mf1ARyisVO9bb8KwzETgzyczBcx0HVjxCPqlY4nc9zxOgDB+iuxwrk
wQ2OWLYguwFXIpvTPppbAy9iisALjdVI/Wl8Vo/uTtTpizecp8kr+MiP13kYMj/h
NZNo1nzAR49coS+wsSh1+viSAQjloGAh3L+771drvY2pDQv2NVpf4ujAO1CvyKvD
KQvpwXPwzZyizfhzuVE5HF6tm0xBIwG7eSOEu3Q/YaW2Wdwm2skDJKM4RsDmutVw
/0WcOkP4F3GA0Vkvr7PK5RxcCsjM8N6fcHKDE7PDM9VtYn5Nvh9jUBqQO+TbcXyf
BH2OIuS1Ux4FTct/qlZkkvT8y7+dfF89KBA0/FzvtZA/SV3e/6Cs1OfEarqLOera
irSW5+29YMxVBubeBUytezrRLe7SWVKaxbpI4gdVwuiGMpnPCyu+Jm0PW2KOl4pK
wi78YDlE4s4kXaxwCZ0pZhNIe7KWhjZktmY/97/4hYJMS02R+2MUBbP1A87GlCrx
UKsUZytF3qVuabF/YFUO4uc/vNLy/otgbwkP6tLwZH5jimKocP5D2S6XE6Zibqx4
T+xqf2q49mYfdMSb5/qlglISHxTjHvaCtclIa2BZ/JLpTqqvd+VrWn2pVvuiAD9p
o8h+UBCWj+uLrWKmzzDft/+MVnJzEIfRXTg+jNOr2MCipirNzH8p5zHVg7dMtBBk
nQqxb9tx5INRJ9QUTWlbznGeymHCDddRh4HVg9PgOSqcTp6REb97PjwB+GztmSeX
NG8jS+IFp4JqqP+guSb5auz+KBRqhq3E3jedBvIzXfMWxjuaxqHcbMf/b2POoSTN
RxAXJWfIrWszZ1ieGlNwjcEAEDalPxYXmNx9BvtgONrrPTEtUIdR1nv9uSorKHDp
xqcGo+nKJwEn4meb7WIwH+XGc5aVWxdpOF3v2hldpIhE/RH+Tahma+eesz44ZHYv
E2oYWf3nEltlGCFRns7ri1/b3JaxBIu732UKnx6xkkapJXGNhzXh6k02DcZhkk6Q
/Z+lK5bzcA3COCztrnPBLfBbU4maIxvQT4bxp81zprVlro7CmxmXLB19wcqqH0AB
0hG9UjbICTgGtKbvlC2Q7GVp+SIkvyoVpKAXKEENB7v/f9eYn4VPOWDXP0lQqetk
9zRt1hxVJP6ZOEvGFbD828bFLWKYtDuny0jVHN3TYOCXs1oJMQFg/kAd01RfqiJc
0h5nKq1iCZMAFWlskgBlLvm45ImBYPip7QWMz65nq+U/Mkcq8yUL6momvhwDYLMs
XQyylZnwiCILaePL+HN/qEePP8uNW3NJNfImUQWB3SoTBx80ESRM9Ne/XwX6UiHQ
ku9v0LiZSYH98MjSC5JPht2v3xaKQg6bmpX2ci91qc7RlzLH7CGPLnPuWsn2cL6m
Vv/1iEctURI3IDDnaJqx0YjJa5TZeu9SWp6b70KrwJZKDyKSC1qFXrErhtOia/Kd
dpVlPSdpk3DXJKg0ZkMGZhs5XjNXZjp3GPBg8Y1hsPJN3DR/QskWJrNK+jgrUh+l
PrbGPvJFXda2bEUMv7JV3WVJEtbOOaMsm7Hm97to9gMKh4tPR14BdDSiG3Ta8PGN
rby8FqwHAQI07GHp6cLT6acb6C3Hn0wIdci8WMu4yVyKVlz/wPr2CVvgswQdSLui
xc/ib1Vrv79CG/7pVTyUOMvH+VofIt/WHEZ905nXJMEZMmN3wOAIlVKYtHhxqnsY
SvKPDDIrRr0YkJt69N/lSWaPmtB8gjMJjVmiCTjsITkSS9M3+NI+iUNsMZ/zQL1q
EmSePt1iXLMIDZRbpikGBKKm/2WoFng1/xXDZ9WYGJDexLTB2XK8SXsja/5AP6Gj
2uVNEQaggJ9BqdRFPsEYd40CfQDcuGmhKvA53L1hxT8/FV/rsxRn5Qp6sFo8vXN4
xt7tDgAIQH0aMh3GHiX58B5LJ06QoK3syS+WuhZH9BVYyzB6maYxHLr48nqP7rR2
iQZl3Rm8xokeMRjI4dxTNVmNUvndX6WT41qNX45aWCHOd6w1zXDXXEAHZ92ASZ6e
wvGMRLkXC+va8BBSMVxRPIdQ2W5LvhjzR7OB8CjNVRT4lHumrrrvba1GL/YOJdYx
CgTcyeHdcv2SAHHAKYqGss/UYPQbYAEzw+l8ShK3Y8R5NZBlU7M1MKbO57FYYkFK
t0uDQFUsxTZFCPhnRrMFkFTXbvJCdsnJj2OViaAywiFyZWi9G2fUpOUqxPycNrr3
dWjXeppa70Hyc8k2PeIcNuvjM24whE4kbsyKgzmUzgpX7sjN/3ibcms2K28Kvfk5
RD6epjqkaz33qsvnmJliDBk8jZ3ffmUEMOltDZkBIDBNEjuTqYYPKlvilvB2po2Y
pwWCsKmdH8SDl0KyQaqNRXFAjCVKSQX1EAHQGzSJWItxtnDDl1gI1RYZ08p4voPq
csB1CrQ0+Fcvul5hSclwThGVyr3KMwF5Ubgc2fHn5pH1m2RSFFDULdse3T0woLNz
lhXi1u/VqdO0QOoPcuolP/9kpnrLLw+FRQde1Jgt9+V2onHJjwmrAv1U8kvJRqyC
DDJdkkcAmJLWMhqAA4oEa/+jlmVvaWhP/uWHW2h1hxPBUSjqw7rm0Uk9A1tcMAsb
z2ApfFpR4iYCq+jqJFtZzVbN9szXRLRRo0TVWrifhoxewEYCj9e6FqVgEFmgq7c/
sO4Nwb1BVdxNqh6Yr04jIU0bKgLTMQS5HFPWMV3hLnPxsyPMtIfuKdvSSnUAURTB
a1yF/u/NX+ylq2vHzxqmejs5lwA8PIrNYabn84lqoT+ZQ968825O8ElpUvZMuXxL
RFOnZKP/hPLVlnRlJOaUSL7DTXD7/00wKUhv2qdCCKl7SVc5NH8OyiRDn2tBztGQ
YUSRf3p3wvY2bdDuS+b7z90CVBL3p8WXqZVn4S4APL40FftSveVPM0ExmyY0zTiy
VfpCpDG9Jk2wI3JQ6gbn2CIA7UsdhteoxoMQHIVY0EII8BUC/+UjgHapSKDSxK1K
t+YTIbE88/R/T2RsJTPYJnHg2jhhjIwL6X5i5K52zdqjErC+oCSysOWxXLvY5pYJ
XcRvAYO7C1JcRU57Nlt6ozJEtIJo1lclODJp7C8//14pd1Z3lNZQ6leFqy4p9yV7
991/mw6PyyIXnv1KDmrv3uw2ZaY0RaB7fsLkqJLf73ShhOMddNp/eKJp0n8HN6ij
SWsUV8a2oZwaVb9T1dNLpP2P0hNHjBl1K2xAbdPCzDn/wSboJpGRDOVjIzUQg9+V
FGiuovcR9aFbl1sxKXyrlUR28DahpO33LowHq+R9HPMSGs0/qxihYUFvv+ZErKo4
vWGupHSkDNIyjQEzXz4osds4dc7J/Sjbw8OwaHUR0WIZTdL3ickCwTp25Iy0klgu
uApqotgywo2qfNmF+t/eWtY/fl2uSv0VX9zfy5yg+UaWNvaD0AIAD3lTOVRUtdle
v4W5/gOS8Nw/hl7phh8x2k03ne+iQCsGERaoJY1KSlB90M2xY/a9Q5PKC9GJvb+s
RjdE1goAaOWcXUWRjCvwr+DkCiTWElxSHNiuLBBUr0AeXqxmkVQnZD7j99NfjQ3o
REDTXbCDqelbYek5KOdnZ+LEfed6x/9be4R3lnU/yHQl92hSg+lJAdpA1wREjWj3
au0seB4IUGxcYwW044Im9eJOsncmToHKfwdLsHvrwtzxIMM5Mr6Ci+nvWRbyHSPy
K0qb8m9SYqdWqN7ntD4w2aBZJT5j6YtWhqbOOTy+7PWWQtm1uPaDt06vIHFHTWAq
4j59j4oMlXYD/LzfTn5t9jPpYXa3truwvSnV1cMEZjo4mPd3up1gjwZamJa19UxB
J4MFFPvaITaElx8tPj/TzcewJztOvIkmfSfnEBZ/Sk2D6HuXnzvvlTBLWKp2xs91
z0BBrXbRFrIvlmQyooRmOWNAZvcCoPE9zFBeZkuRKqjrFaH7CDGcyQMrk7dD8IGr
A9Mw4qChfZhMQZMleoW1IJ8aHQosSokGNXtQ5bnxnRdkGb0UzdkLW7qq+Hcg1G0U
vrqweutnCqZk87/36k5NcROin5iUygy2TfC0k+xJwsJanGtTvsCkshGRR6Pkzaj3
iJWs4vP378dYm1CIw5rHax9iUU8wA1Cckv2hu8ybpERgawtvguFlPro6KHhgXcqo
EkC0oNBWp9lCs+T5MlZGxxkzBZnYOobufvEk33X6CUapCe7m7oJ/m79WN0ZAnIqD
lKMd3X9BCiLVyh7pAR9EJSb+wPXvnIbrkzoy9YpNJHTHzlDpq4caI2qMNVGL7cin
woBwtGhQS2X/4/syyoP+4IPw1ok0PvghmLG0ZnLVA3AIULKNZ94ZkNhM150eLaJs
R/EmtwIoR8XJzhN67/h95X3REmg2rhsVfFuxFUPZhIVLKMOowCUMGNJ60Z5I9efh
+g8lze8BcyKtN3qPPxPTVWtMa/XsDUfmROIka990WECKZ+W8bIlOnt+yXyVu1bb3
+bUsUNduMlMQ7IfHXrsI9EvkVxlh9V/5ZWl6JzGjWtfWoDIFaN0dleBso+xODM9h
ZBs4WxcXUpiVT/X852MkgNsKtQvfqDifZy/2LI4fcpAG2OQbs2z/q2tXOOXRvLIi
+EYof3J0rz42kRtvWA/jOr2BI31am74Zf7v9gXlRDqx0cKGTWFg6m6r9q3dIofL4
SpdK7ASKMmbdfJUaQAPnQdbaVfYQv+e31DnY/17vZUl39Tr1+q3Yjc7lT3WyL+Q8
X1jZcgfz5Jc+ktSx0l6oviFySozwFeHUkk0vFgj86x54uIAm96vdVf7mMOtkFP3/
N+A3rqg4rE7HFgUrvvpcuzSI90dOp0QTYcU1dBgS9gnKRuTp3x3CnFA/7fNEUL4X
QSDgdbgQpIxu85Z+skBzoYuWivLK8/Fom0lPXZXnHlr3NJPg6CECoCSUE3Fzi8ML
yOov0wSOZIliVCNJi4Q+kiv32dbsAL5792h86mX5bnnQfQhO1ptefweYYWamRcL2
oGeMDBy0WsUR2HFao7NLMsQYAXhhUPmg9gY5NK+zel7DIDpNE6h2JHs/poHUwAbD
AI6yaIQRSJUbJuqm9LjnShkJRwG0ScFjvGr9jrvCYUGNe30DnRWLs0d80E23s/s9
2RMj1lhmaUiF/FwS26Nhg1NdJFugtf7BOaZgWtkXZmwDUF68Ff23f+WhtFHPv/hx
O/v9t/qCzMu5z6co0PAA+7e/byhqB23BgKgufJ9Hv7Dv6ZGIGemgeV4gMxUcInYf
wk9ZaAfR6u+97uGRs2/nm80PLy1PdnGJrcvNs+LIHGTZwaBG12AHlXOJLg1eaKTo
kC6El3Ai2NEdCrYulO3dQMS94x2TN+84B+qogG9LPIbJ5WKzT/YL+6NfGUA/FZDi
IPWsmTZdXEYjLzKY7WelvZwaC60Yo5mtCIePDXUzxt4kGR9EoP7B5HKjrNfyOYQd
5dLBzyTofucds0ILd2YD3oNDHKKl+MKR2SZPZVoebLribya5OJ+pLKC8xSGx3RJL
HsQ1kcr79X/BQ7WOhPBWEkWldXqnztnJGgPjzP5IBJxd7ajoQgM2y0JQu95hRkvN
Jc92DCORdP9Dd98Js50mxaD08U/yJ28vZdsUFgD8uT9t/jULSZSt9LlgbQXfm0/s
rL0asbapsyiMGRfru4MvEbGxpvoZk+wdKOPppDGO227+AQnzIEcYCUkg8YCIDGVm
X4GxxMLZzAytvGNX/72jDqlurLanTAEc4MKheVT5MWv6cp/BW8ij1SNiM8nmm0rC
JtkSSwxGlLzXZA82iilWpfPkoqQ7iDT5jGcoOgbkyHSoRU81dziPMyE66hlZtwgT
vDFl/iGJeY5m4BJqImUqN35NAeaN7dO6nCH+9UtngmfvyaNn4HdRGdYI8vHyjsDg
P3nlAE7msP8Z1vXeOHR8WBxEpQ5/I1T/PX+si718CNXZtzoggCSbEIG0BoYoLehy
nzMLkMhy/nyHXvGyS2naei1+usdSR9/oYB+ECHds/WIfdyO9aMyy62Ni4FXRUFA+
u8ZNwp86etKEatQop7etiRPJXfIC3HO42F9B6wBGnoDczx5D3ej9YMUybq0trBsu
X90dlboQM/oMpanLL0jRONd05LfrX2tyIXfANXoAYBHWx+ktEPFJ7IJYMyho4eNy
OfB84r0dcceFbNwJ6kEhTa47ImMHZvbxRDrCws6KM5Ss3ZudH366MXLWr8PMnJ8g
Xsv46Q3+wJY9djpwfCVNa9n4iyQPkpoXQQ7dcREHSQ5Ro96iv58hzGkYIH+DEapW
HwStIQYK18jy87p++IZCXKteIXMVGn2OZYF/TdSvBH+9TwZxcMxG8/cH2DT/D3y3
xAIrGFuQZT5G78LDjhiZjaTDK3avnch+FdcP9EhIwZwSf2OvrsDLClz9pXgwnEnq
QlgqXfA8p/V2jt5uA4IpihmSdYYVNIxlI0/asG5BU5W2w8nJU3b6bjrISRmgKT32
qVLzG0j7Ru48OxTiHDLZ3j9DeKHy+qq5dA2JAGae4l72RSNfrpCU0keTgQcLve1B
Z7vlrTz7IQ0iL/1H6T7RqRDLU3Kmn8zcU+pS7OlfUbQ+sx9CvJbXWGGPtlRTBA+j
SjVFNk2IGGg+JtXpEE/5AFKxMNkKZzEfwqmElwcqZznzhRJUgHcBLywFJpRjIeVJ
/WkzuxPCCL9+bOZco1xcuMq036XXYwVfd2VwkaZDZuQPDyqzrCdRrHgz1tFSwn/4
nCx1T65W9XmBJGoRRXoa/+d+D4GxgoTlBX0fwk6GCZ110dBVVtT9/R+FM4+zp6LG
HeiMWUIfNdkX6XKXPUyQYk4FdF/A84qN0lymd71KkSE9Z1OgJ4LVJg1B2c7UEyEL
QqHbjJPzCeTQz8yhd9N6cqA9CER3vF8fnnp23iCTvjiMK3ZjK/LpSPJHPJMlwyK7
R7D4Dmt0HKXg+G32VNRkWrl9mtk1ooPcOtt4o6a7TsdKfjMOsu5o+8onXqnPJ05l
RoUZ6DAfRAgD8rANEjsFjOC2u/7nvsu/O4OWIxUaByjsiencKTRwV33GZ22l7OOv
cT+Qki0xFOAAvekzBIP4mKuQnnKbYk3FVzadtHRziGQ3KCV9gnhbAt2SNkVGVIf/
T1kGMKPo5V6ar+RG4nPODtxbMnCPdasbDOBKhEBSEi3/rCRyDUd0/jF266vmnzKN
m4EUTwBTZGD8EhPIefUDsNHBnL6Cy84nqpGEogPcfbMYbBZU/95GEh2KdY3+YDmf
MIUqTbIt4I38qj0FQ+KMMP4ixpYZJ7CLFaGSuGMzPVqLhxWHcMksY/NE5CqYOdTC
FCVXwIM8MilR14rovPoOAclQFbcVFAG4IPde7b1vb3QWa8GFMMBXNyoyI7yLbNeJ
bGBX3OaikEYDnCLuBwH4E1WBJA7oxb8i8GTE6mh1QvvwODocmy8e4f0VHvrycsiY
/pdaqs47NAnzOT3mCjTKLdr+6GiRV7j5UkuxPbSKfilS+j1a8+9+VcYtrbgmAC12
KfBYiYfNbHhA4Nz7vJYTs5W3QxA14+csmTdoHgBA65E0KUq4VkmilSyuhrb9lX4o
P9h6XM7AaIVU6QTs8WfDWFLGUZhSw+ynWVarPwmoWU13McfD496xVkaPUJCohDH/
4SDDxOMM+Nu5n6ARzvpH7/0fjCF8vwGT3idWzAibCKDH2o2e7o8YRiV54eKyh6bS
RloQQn6yOlUUb68Sx/YHHNCfIZjYcJbaddi1f2LsfLiOVqGDzKWZ1Y3lwDh5pFv9
eDRvYmNk4njyGXAz4/Jgs0HhbOi7QUfa4MwDthnCI9phooV8zKzFIWjA8XFBmXXi
tEWqtG7Qg3qxzicdRizNROB3hqMmpX9vt48LwzgvYxVPjVM2gWXVm3G94EU/MAfi
YhNCvEqzRBhAb1RIQmGHRmxOfoDore9sET5GtO4E60kbpUUaoAOXaI65ZcflPT+A
6Gxi5XTv0GxqlhsSBF7YjBk493JCK/evVzw9MxBEg1q4nSQiq1KRqhTO9DGyRQxv
a9n5IsqoopPQosoq3eC5PJxx6cak648pIE10IC4t7UPkEaeb/eNrJYYipq7OIULR
LzH6K3RdpF2MxC0YvseQajyttxp4F833eXKc8i9XD4NlxJVQpeXH1pmWVPAIfP/o
7cHaDgMvG3SDKGPYIlL4qGpr+LrrXag9arl9OzvVNXdsEm4QPtnq+zLNgvNt/AaL
v7Zkpz6kCOIF1+e9XJP0OKDxOjKH2GzS9SwosdxpvGRgaUB4myDvIRPRjZsKczUt
xAzxXVK5zJ3P9balq6eGn76/hbVwOPmJNQ7TflKsodpGRu0Rq8ZB8S4l3f9mMfiw
tT4fLu/BypqCbLvK2Rng3fiQTp69Rc4+DpPh5wDnPhkmZr10BclJcto8LwsU0try
RN5haHw2xcwlF82GpApymn17WJQCwWM4UjZds/goNBNRlCxhZjr26tuQm3yVCczJ
yIwLOg96p9aJgbgQpXVT4nE0kYdkGesBweYX/T1iflRfpSQRSP2orCAmOyXSLz0t
CvZx32PNIcPNlzqFtsQ0/xmyXV/ZIXwHAJiS8CgeAj70pMzsF/884akkTJwiDGp8
rFLlutd4hTkRDiPPPl2M4ynEBgKIyukV+xccKWgjqtrvV31GxT80S9UneNRxVvKE
bru3SintoDJuCqY0xETkVgsj/LFxUceSSiWrC+GqPfJ9KXjDVxHGaQ1aEUR2k1a4
u3crm2Q9SbjNe2hF+N8utn58ngLRvZhNlFSaIihuMPJkm/L/lbC90MbkB13jZ1uX
6olTW44dqDtyxidRoErRxj3HE9xWKfqTjY2wH72BxEq5lBxySZFqE3vFg82jQthm
MarAx6RfRKTSOOU+eaHYuKkAfU06eXvXDEH0tzIjB0Z63PlZaTkiAEOR6cz1tXXd
2SAdg7gTOu2SZ1CnGY7we7T9aL72uwiPySAOahXqZgfxcZhHPkXHgEWtD0E32ksb
Hpcq8X4rlAr+lFdZVsIrY6z3VIJHcIfcQAzqfagaHjElYpQJHfZ/wfloFcH3U9Cu
gcaJXsYP44phfysMmOAZhf+Vim23PCyqUWJKqbE0LFNDCBlMAlDrBls3OCI++tSU
/NROvt+jU2/ZLYOh9Fiu8l6OqExM5RJDDBdlXKrAw9igBtBAmOmpIRlepgO1W2CA
FERwKMPcC2Ye9YzTUiLHuNUG6J3+AJzOgXc8n4ySI2dohsY9xDFKrWlP8j8eil+f
D3rNu1WAcsydY7cfd3xk+455ow3fpPteNTiM3gyHeYba8ohgJg1BVF0nx6DFstkM
07IyzV2gLJc4w3hg9XH4NHPGkCMKxqagv2v6YqJBMvccCJjFhFJY1qxSiSTtc2wN
WjQq+EkDcjtvFjs2PUY6O561oW27NLn5Dtfyk55/Lt+aQsr5hDc9AtifpGC0JK2e
u904WD1yZn7LKFZ/UdhqbgQG/LkzKWW7mltVim2thxaSsOvGxYo5A0vzdZ7p3yUE
SIb+tzZLxlrylT6K2tq7dQk9xjV1pFyY3UiM+2OqEnsHCrSG/W5p5Co1wHCqa0+P
fuAan+dHyPLJyunmRqmKxp2Narl8hMcx838QDcuSOw7l0SbsbxaZ3gBUxNsWctyc
k+W1Ey1UNdJeCCObVIKzZNtE9P850G7iylVJBDOVVihVZ42nSZKVH2yO2081CG+E
owE8EjpKJWIWrSyRMkN+UXld5nDr5/yvKW7XfnxVVrplB7moVW8JGPglxUs6XT/7
0IMVwnByOyz8zKMLYKG+TyAYwB5z+oohdsWENAz875ieCR5n7eKhgAYZ8jWDQQda
gCjNiNYHDRzMVScs7LQ84ZNB6TwEupvKOM29yoraSBFSHw+uLWziMRcGRzvVzCWD
INPiGvS+D+tkhtNn8+cxgVHNZFy0QTR5pQyMIqqslH7vLR3l/UxRYY0DZqJqWUkF
P9JXrVqIwCtxcu+CmTgRYwt9x1H+Udp/a06BPInv1sgzJtDhiDmILwYnJqcFaw4A
4ayk3aDlCjmFq/YhZc95vGg85A7iU0bE0iIksH03zTT/pkPiW/GoOUt810rquZ26
39Y5JUst4dy0Etqzr1pXfzuNOO6NSMs7V9mmI2Y9akmHMuzoo+MW2LaqBMMGhW0I
6pmLb8RUATyqCzBVVXnFB0KMfCD7ClDCeHB2eu00hhafUk4iMNfJImU5AsawickU
KtKSpw7rM3SvzSY0mh0hqlY5Sylr13n1aANWrSc9oE0L/J7tiONRwfmUF0vYHRk3
cZYnojU9nJgXaJDAKnHquIxs7eOXrIjFXl4E5AsHeWdA60TlkDjzAWncnqBuEBqf
hfeCPeEexoD4n2E7ytxZe4SwktKnB/2+jMjrNxYCV2UXLXAOwx1f8I82CLw+qwry
ysVivc1EShyXayIqA8R6mJzO55c5sJC7N1uLTBW/WZN5pJ+BVuQghld+8arYGIQe
fLj3eo0vBFqlH44JJV98u6vEnVfnh3fHw3CADhzXBzZzM+xu5rw9VUy4GfbyEgMg
Tk13vCByDV567QnPqSyYorYd4I2eB82AUl8zLMrN6Qty9vP5nrPFcz8X/MyJ38IJ
80BF1DZwjhwNRdWyHh5p/VORQR58DWvlDBLfPUNTaSwxtGJ9tjZ3MWWskxjXsG3t
L1sE1ew1zcCl7LIFoHvZ6AxJimwnZvcHLLY0Cvbw0AEitR43v56YhabeQX2JZvFi
U/OLe6IOXFw4LE/qpbdTll89R4DXFj0LrNrWU0v3tWuuyK32hkGd8dBek2m7h9hF
jn+1vAiLc7q1Dgag5Bo0GV+nj9T+DKScy9BB2S9vkbdmuNwfSitJ/5wPMf9xF2x6
73b36cmwpevGdkw3SXd1UxlvJHMvPiZql0QDBcjUEAm92zzDoUYggbonqJ621ZQ5
wSvZG+1NkunrM8DGICBUEy3PQYA9lBBqf0j80krFPPLohOCe7HEd3N9kiSJ2HaxV
z7RXHQ/c8iz+djRBFrAolebNdBc9VpH05dOy8Yvb3m1IDqoqtgne5fBmgdKEZiof
G0FBiwsphFCy1RbiAU4FYxxuyFSkLUrjbrwqpABCO2IB0ySzN3hCDTttVOg8X4ve
Htxto0u5MFAYv8E3Vy9D+3eHoSt7eKSsZFz4axrvVnAtgIxhic16O2j7W8KOPTEn
+qOZ7I3bIVuGsuItINmEG7NcfVjc4BaM7C2VJWR+gCdV+RuybTSv2+0Yuwl1sONl
Yn9Ey2o5IcRdAxpBmw5aWS+OtKKZ/MmDUEXwwsmPJdfnIGildzE/rXR//10hAV/7
xFidYrSMPCFGQWvTgEdFh9F+yUXrkhyLZOBwoO/Dxqv4UaVpIJJtGJE7WybVf0v9
gofs+QIWCXUy9Z1FQ4mm9tIqMvaEUBo8Hmw1XJZwB6AkmGW4x0yd2APFHQnzeU99
zfVsNUFFu2blwpj9pYR4DU2LH6t+XhtmHQRgc1GXThiAuufAB3eSpDOyaQ+E0UQV
wSQkzxNjEFGkGbDpC7x3AUh4NevSGyeUtVzPRICMWruI7wcdmd3p8Syp5gGmCn9c
IL1XwzNJdg+hDT93mi/DDu75O7/SAtuTPaXLaGPGHseeL1LgTuKi8gFsmJoRhqz0
ilAZbYXWDdlG56bTavTrQU6cVZOG6hXDg5+oj7BKoRPKipwO6cxvOy6wfxDXDDmG
RM1/5gG0jynWYAaICzDTHzFjioFoyjPAvT7CeS0EXaSCDZrc9LA3vXVo55bUvJJk
EBPUpGSBtvMo1ld8fGHZTjC19GoUKA2Khze6sf17MeFemI63S3PNzk2luHNzWUUg
g6+KUIt7rUFIG4GLF8XOqEC5bjJ7poLoxAl7AjNpKKn3nXuV8LZYSiyscaybIiDo
t1zrGdK2nLPk+2qjR8NpH6t/WFAke1RkvMorivEbIAdGiRzOriR8r2mKbPUyRa6f
rkNr4TIrMF9s6Ns3NYHXT1cCB14vFgvj4L4flSf2b0zxwPRwN8ZrputvVwqlZnsU
y3W8uc/3G87PDd0pq/a7N+MU6QoRjWy3vrTq8EQVs+HrJrEB5P1w16y1Vr7QnZFq
pSFgg6Utl3yPMx134v+8Edx8GDrjsa0xiKpnu8Ti5LSZ/wClT1y8MxydlMkkOYEw
VLZ66GrI4Y7dzaP1EFfX01vW67d7N6iSxcOq+vGpvl/z5NqPhFslccqLcAJVn4Ch
VlzqfgS/wxk+q0NuJo/D549wPMkvvmaqdOqfLbvdAVvSPdf9+WWWsVa2I43w9qG3
qhQOyR/KQOO1mMrrP6VSM2fBFyg4vCj1Be+QNiTy+uIbRHqgd8/16c5ZjBXt59Wn
dqTLDE7AeYdt1b++7zX7nEoEyVVpCj7+cs6Z6AJItkKYHE+q7hJ/tI8Xr3t905/U
IX+bvhPOzqbc+Gvknxqah47gTXYctkg54tn1hPRV552iFxaDIbxLFqqdqZMCQNVv
4g8j6qyp8BNhm0f0yLJaXX70dp0ryfZDEzob8I1CfsXObqkJY5xbY5rrSJELUZEH
0vgtKU1qQslkEKiYorMAZESDzQTxdCsX2hHu66G/xVjbDZuldx1L250PcHJpoNEE
6YLmdPs68DxFo+/2zLii6hAh78w7iiAN+iM5NUZi//6kSR3nr/SqvkJNBLHLSWm3
HgxET/EKwyiM3UcwWJZoyh53aSvJLmYYCfmT6fAdemmd6uLB926qUgU7n+NrK8od
9UaupEbdAFcY0wKkkIkj9gpB0Q66BA7NXiNSVa0TyAe66kF5UD/FQGDzQqOQetam
c9NJPiH6x9dh0D+sEn+hKiUBCSbJx4JL3ODvYcqhHLrX+lbZBy3ntIvTBp/+u6y/
u4W7FASgB+GtYZVVqfBPfeXIjqwuM6/nr+BKLDBK6YplHYkMES0XQZGApjg2Tfqy
Duk5PJ5ipIJPu3MP0hNLAy4kjZT2MFaVcr0Q65lgBrWC1g+heC/fw7IhG/PLn7ZU
+mYbo1Pty3F/NefwBXIPl5MJRQylwsmF25M0QLvsUb8pJnAs2f1Ccfz29roWdFbG
oeq1qyOgtqrj8K0K3fuWe6Qnuq58LGfr1Rul586qYNjz8/tjkx8IxUuRz8UKnZQz
jit9LqVcdBIWFSJXgjrBVUy+zr7Wwr4oB79tlVJnTLpLQOhTMl2J09B//dBqL5Cr
q266TuOuGldQhTn3L6HbuQLNdh5a1Tq52T+nobsK2eWklIIBOA86CnYmagUQp1V7
7uPcZDDSiUBQEcsaLC5ybMiAMwrTsupipfjSIw4+IV8H5NmWIDKS4COdzYHUXxTF
7MDmU4QtRmbiQM4sAwWaxAtbOKpaxJ4v853zoCsYav8e6XPU6w7JtrWk8rUFaaxl
4Azyi2MIvIfBN6o8D95Iq7LbQ/uJtqkeYrTtcToD1V6ljbjS9BUM51whUhkiCfqZ
nCW+WExe3skBiBq19m2hdOgP3EWpLYDOMzwd9yTOR5I2kBrXe98XkhqhAGmAl58W
9+1Y+dhc95ere5bCq5efxLn6OIGzjzl718rd+nl4qnF4hwNny+93KbjvT7+1cQvY
EozyapJqPafvk9eUPsuO+zTz08Rnu7uxJIth/GHO0elS+q9YK53kaHLNgvDWOF2G
QWygRwpbFQvw8a/xdDD/z2SPZExbfe5trA/8r8hg27No+OGd8ldPcq9pmh1tF18m
f56UGO35aj9dPg+LzZfluquSaKiB/MYXKxcxRjwJvGGCGe3Kztf4moI4MqGTo3iV
fPxrioJ1N0QcvzM0XD3SG69heIJlkokaeDQN68Ts0bfWB1UaP/NqpL1cP5MMhUv2
o+2mjLe7I8JDZZZmB/UiWHTvFswyArQn1Z+fUA6HnvgHn2VDI4yO5pIxVykBgoTu
gkGcrXenpJB3ceAqJqqO+oyPRCfpnp6SoYOxjOBXs8T1l5HI52AZX5Q5TkVzMDTU
lNKqCWsPKRmKJJnkC8nOHOfg1QxJJpY+t4lha/1yZ4eEqYEcfhajG59RSjvNh1wz
KX8azwV7LiGf3BARW/83G41Jm7zJTl9hHuq68JhHFAqFAbuKV/v40hwef+sWRjWs
k4UcrYKQeIVByN5ImVtWELDNyla+oECkjejb/HHneV+QVMgP618FbXLdoKHx2tpY
v/3Z9qSgnuWVLnXdOttRZsBOMFx+MSRQXNibVIx610FuH+e3131GnqNJi3Hbtcc0
qtRAa0y42WfDH8PkfkPnOMvuPSQ5XPvKTVGm0nUE1Cxpnxnym1M60eDhcviUsPVQ
KW5IgDSPvpq/wN3yNQ8HXMqTMkyH0EJQs7+ThnqKNRXFKYGxdQ15Wm7kB2oAttah
ZxyHtvtDLIRujz6y2lfKdUielqD4BnjTEe16TBwnrWt+Tf/ZNSynk5SF+E1QXUks
xATlaw9b0EYoHpwTkUMAR4ImALgBe5AYLt6oLBt84k8coCB12fV4i9GEnZWYJ+uQ
pPVSo+ff4K8EN7yW17AL7akQ79LHy5qoU6CtRcd1erRD/aUKp/K2059ROOLAeLEX
yAWJBULDQk178iza4TMQ+UbUFJLDIeWI718TCkHmzp6qsr3eE+kRkDQZyAXX0cWo
+yoPBpOoS2p0N2VaHKtYDM04+StgSw4h8AvWDqDQZvMhguN2TcAioDF3j75NOGMi
1lhsBhjl9Pe75azdRGkOzRQ3C5JtA618WIG/LdP/HUOBpi48ekVQmnBDGkvu+lo2
TAWVRkyiAhWUmgw5ESUv6cpRLvMqPAEl0lGnSW9LtfU6yqIYTj3qpvigp23hgtwj
IlNL3/bx41OJYQ3OlbbQcemHqA55iw9yUAzStWtXY4o/G2LWCf+55/poqKpe/N5k
33IBEBwjN+ACqv6zgh72cCtJ5RWq1UvUa7A6FMiF1EYqSGw0MbLjz9GvjPWwIYbB
PEYZ360dJXfXw45QIxOaq/oiy8mM5/swCmHXhOS15LY0LEA1Ewnh3FGUW9CfVNj4
9nbe5fFmGS7ws0CKT8y63U2sj8OD/b0OsqHx6qw86/6LNVXwZ467GIK8XewF1gsA
90uQuUH6eHX818cTCl0aiaxxSMDb7g0e31Iv4B0hbiOmyI+aKjgPxRcT5+C+mF7X
7QMsH1XYwdtfd8q0JEDZ24NGjdlQCddg0vDicXWI4Q62QAAPB0DQIl1gMgRKyXVI
FMZmcIR4pA8dEAnt9Lhh60Kx2PTpL8tKQqISTKKGQGkBIdnImPHPpxIw0W0Vn4VI
KYWfP2Z2aK3DUaq/bXwWBW480+TEqBNhNt9azpc8WDcAspkKGh4sPEsaWi3iv216
HIzUrkAvpMFbwrbI6LzGJ2vbtJzNiIV1wEZLt/exnfS4whOZnYTOjdrljJrrnGlR
V3rvYv9uhGTijhHx+zJG6pIQ7xJck/26p+ZfTB6Mb80CfsXGbVTPMkXnq6YW5Gag
uXccXe5gb9ZbPh5Hy0FTbu6zmIF3K1Zs+dDzyQ2QxLB3xjP9MTZ3HMXoAqUinGEa
g3+Quw1hYlOrQBzh4B7LyxWG3NMhNaCk6blaNRbN2B0taPcTbFx2HLs1ecbV6FUm
gGtDQ4CU9NKE8Pm3mqV64E3xh3L53Z8Kjn1LPYQv09htP2XGrSSf97nTVun9848m
0iCCc+KXUFnNj+3b8362e2ksVfgwJJE5itoKYJG3qdUXu1XZ7vjfoJh5HcwoIr9v
tCfUBxCCVzxX+vLtF1iA46KT9lbgYqMcaUbmKojGiTuWBvcUi8fTO+oEjnlgnZO/
h9twSEcLFiiHwM2DPcgGF/A4vQjJcKfNnUJPKS1PrTJXRJ18RgqYBwdYpU2JYZkm
YQfZBiTYBa4ZAT6Mjt32ICz3mZJu7DYUhDIr4znq8/zFcqzfaS+sa0ayuuNtobSu
G69cppitgbqja28bL8Mtu/lh1ARZxLU3bwhhBfdZ8P7gnJVeFyg/gMXKN4DbJDiG
/ILwZNWS7236FSUYMdRXFH+C43BEd/WJnA+oCAKO12yDe2Tx5EoJ3jigK4disV4r
lKBNmrn28Qyd2LHkRXVf3qSDXoID1ap03MMpzHWRPQ8Qy8/wh0/heqSs2uFUeBY1
/OtnPeqxw5g4kLIBkieiJRJvKEUcOT+7/RlY3E7gfM9khzilrLIP0gVZX/8Ow7CJ
W0JpcbwfnxIU6puEWymNMQLbe3hNqOC08ursm/SU1IvWHY2k0iE6FmrlwH7uRTJT
r8Ca3Eiv3ccNOpVIDY4QmV9S+jDEBIkhn8B6nChvXKIO2roNlpmHSFLsXlb+I24C
r27g1achE26bGyuTASieI5QTjc9VPVI8X+NorAJ5nM4v9Zd53jo1zRPWlKH3weLZ
erft8Jr8UthJCiOVW7kKpi+dTgT5Tn71ky8EuFaQcGtEwvuJh0Qm4W9r9IULoJ9G
FVZOpSFlsfUNBRqJQWQsFcrxzVkVrBshIjJ6Vc8cc/EKjaX/0pIK+XGlm7vj+JQY
+oJllABqfVHm8wGpunmez9C6uZyQ4iWfVZOwVnDyakw+HgTdiKpma1lyp785Y+xA
5V9jKfX8tjJHb1eaBHFd6kHRLfUEBVmQ59bjamgTxNuQUglfP1Jd/ybNnnPnafWz
dDEO9g8c3lq637CkOyeP594QZtr7XZoOWozdFhi4FQ1qn2eUnXFKcKH+EMCjcFrE
WA8rU3fn0RWVGAN9x8ggET+x6yUE8r7LRbw3bRwtPRE6EtfR40atdm71vSX0KSpV
8tgLDS8ph9oqIsmMihr9cyISJXqfF90d+vSi6OU5Wph8X79GFMc1+DRWtC+Tfh8F
eTsSWORnhiz7hhfeoBqqlXm5djL6ezFe0G97j+fBBh1fo4G4z3TQk+6Twem3TlYB
pd/fNexI7qjCuI9QvCaA/sV6cyEiBwFav5nfodipZFPCYVevYSTDwd9xb+2R6AqQ
U+KczTtGqHPaCgxpFs6FZVgYdIJzV7bJ9ivOq0OtqjsTwo9zPADtMfDRJNbYntpf
f98eg29ofBymX5LV4RJ2w0IXtUUcCJPHWDoIccgdSdYVdT0XMyHdjjlOFWomd6RU
z+6TD/pm3k5kAdV2StLRBAgYfqyR4njJ7aJzXciYKHaHBMO4cX3TrEZNfYTVSi9f
U52c7tvntSWtZWJJLWZtCMfXvT1kWmnycOkHl8wvRSJcPuk9qhxes7LU08iDiU5u
Br7nOW63LB2oabqb8NHQrXSn0G4VhIvRted0giDpdy3JkJcBjcnRNy3W4kCNLPbs
p/18PLAQFOCOlasE0cRh1TYscSMocN6c4Th32Ll/ACjkcbLAbDMaScOVvH6Xwa9N
WlzgWI8q/WugxoG6tMSCpOwzfEn8zv1l8JsBjiMUBatSnelu/j46Ui/lKrL4i68Q
U/XeRE3K/woyRABRJLkHpeFL0e/DUBuHX/y/h+Bi1LqSeKjrkb1YlgFE406IL+RH
nPpTjBzARo3N4cu/8Xz0wpU+4PkGoylqsHR17iTuCzp/MSn0U9vDLAJ9cuNPEE0R
mCp+uTGjEKcrXY0MnpU6YWSTXqAnhmJ4a2ia/8GPm9fh/OTjAkR5+pWS0QxdMjnM
/jKf/w+OMy1rcYyE8YhSOUGM9pa5K/U6psN0LwZbKVWB0icn8/VetJXV+a80HjbQ
4CGJmsXV/uucghj6tcn+++uoUa3uYvzW+oIBGpi7Uz5tF+Vr9pPWT/lVZ3eZUovm
MVZO7dCzNmWI82HJfVrNrc8lR3HnHGft9W9+qYwIcQTYERqiWHq33fy53k61CNHC
lvA8J0YsDROq7Twd68mGywzJ46AazHFkHvdYIfhkXSCeF8ndnlRv2mB/IhJ8rAac
8HcCEggekvGmJl9No+29f7SJifUHaO7Q6dkeiheXIiBUqj73hVqmU+NFcHScSmLQ
guz8HUFWuexBOwrpkWmYIFpBecyu1gIVqa8v3SkY9Kmq7f9A2Rx7SjeFtbHX8b1O
C5Dnk9O7eqHrC/A2+UEfmZEFKJXsnznpAwwHL/1uUtbhWT1JbMFpC0w0a8lmLsbl
PaoSn75aTHNt+9MYYXtkcsANtnvUMDlSlLGv7hK8bqWl8/3Ryv3dUILSpeWSZ1Fn
Repk758Tb97JoeHy7Mo6t1VaL+tz7Gco1f22udq4q58UswVsO512NaNeNh8YdhdM
d6WLjg2j68U6v01KINYXrAIjXFosYjAhpEnSQWEqw5l7zsuARAckVfJm0Rq1+hPc
EetjKnUIxpZkxoWrwJZ7wyB/HOlT96DRZLBlt70JUikF4vKtzPGjg9V4bInqBvNG
dpvhFZ3LT+UUZv2yqVMLQC3pIlz2zbcvi/IQWbUppaRyUosEIzRBE9rXIbpe8xiU
6J0qdGem0WwRI06C562mwtInOxao6sZ/g90b1b6cMlZ5DQ4Aa4N4461CqR/m1VRS
GEypjbDMpDWzP80ILf0zIC3or4Wvvraab7G9DqmcvUiVc3vaKZAs+X4wZNTdKl7A
05FLDKTIGZFmrJoQaSYsUAne2L7+ZUEzFbgdbgXM5RVFmSRCPX/gDcLnlNYnbnBH
v6MTXDkRtMrEbpQyfiSiVCdeZZshLG2CxPlhm1KnDBwETDXUkNXpxRrRziRCmCoQ
xgB/4lBaDilk091p/YumEgPe9bavBgNzcz1K+RHYKPCFN//gqMy5Y/PA2MFcJ+/K
3fW2j6uBenwnr9lcIDCbCI4XkLaoirwuLjzo53jAxShPPcgTs+OIN4PIgy/FFS99
SPC+XV484VtPjakpSWXoUxrcxpoubGgo3LDkty8sXFwqEfN//MBldz/Eemx9rLXw
SYZsNBYOt6eGzpcKTVxFEPHROBlv5i1I3V7RjgpAQcvW87Mpu1WrWn8A3Mq0rO5/
vAwlO6NHq7BWtmO8epekH0bogCXaEr0oKeCTLTrmRctiaZGzoMLl15Q5rIyBLnbB
Ul9OxPJ6aOWrEuzQ11mKEsDPIUHzCPtbbKtmPNUt8rOB/XGpghAeifNX1NY3vXS9
y1Vuq7KTVTzagq6WFpIrlyyz1o7/avYibdKC4h1L7zOz/6X/9Ej2eaDLjn8uayKV
C/zLfE81hER2mvEz9tzF3wM0b1F+K9XCBMONZBUKF3YkK3ouiQRhRT48P96L68VR
bOCOGagFt7XOFNQj/0TEoZTxPLvQY2ypck84Qmo+JlDd8sz+BrcD+HQVNg+HajUZ
v5QV59Okokm+4u0Eq5+aK0s8etJcR9xbbH+LUC+1Qe+c7n3eixtW68UikHgNTsFq
h6bPi8e+knkSlN76hc7qr9lX4r3A9PTIHO2fJBiwiXFIb9a+rdZDnPGeTRfaEoPK
mv6HavQAEzmsvjneCJ6YZG43sPoYQPLdwiCV/ozxDbol6yn2xCTn6F/020gw96Wa
zSk52w1AupUc65JuBM93wo91+8SnyzFces4ndmqAhKTYDEMR6qf++vPdkhf3IhFU
NyMeJPso6AIIGmgI4WpoyOFgI0hlFYt2UUwPV9JKlfYa0u2/jiImC3+CZI6k9ymz
TpsQNlcoNXg8oSqCp5gG5sf7oPHJ2kQvX/Dn+YyzBOTHvV+NtYTlTAl6bkmtzYa1
vGdqvkfBOaIDNXyJDVRfzsS8jfJk9mrDxMYfGw6EdlSAzjNLAmAe3wolHHwQWfiX
008dPrVjID22vgEBELCczlW/o0qstOXXbeUU5ShvyKfIUdZ62dX1knV4cddepMNX
24sdAeCu1SwiCY5d3pzRma1gTmafqPdu0Uf3zm7M6KWCoJeMF1hIPbPO3N07OR8k
MKzq/7utFTaaIUjBSzl2RQYDCtL9iv5nmsYfBzRGI+CZkEHs9BLtmwDrXubWkmuH
uyklu7LkC4wcxcEVt6XUDS0nNWu5qIWde1aWOz60YJYdE5HVMxh2vsfPI6Z44cYU
Ht7+7gkjuTRbgkueGK3tlP4wtDF/FulK/5skOssDFvHKDK9HQ7WtCeiIvp29swG6
JJ89XdGGCEhsswPmdz2zEYi6okBDWd2kk4Injv2/0uj867Mf8UgEPuXYJnBHqCm9
I2LFF89SVcJDJ9QRJWGpCUlrk3MPndKrOLBIBuwcEVJM9QX8ssWDpNWzhMAs4Ysz
NjncEfutrwD8jnz0mOzjZk/gZp2J59l6kLqQ3est0kXG5Hu1QTgTSvOczF+OQWih
i1YkIMtnIMF0lkrBxmf2lARNGacOmMEdsyNXgdZRKFVEdpHNZ1h4G5OSYA+uUJH2
juT6EREhNAd1KUhMBgp8VPMlDm/tuQGKhz7Zn6CUC1A/jSsXI7JLapd6q2+3W+lV
Mwsd60giio2yOK8NDnRQRe2GqlYi2KzhKdISSbCda6tebMQ0WF1CCkv4d/Gd16nH
pHV/8xUtjp5J04HOmvstMxoaAsGNWfGpD+rFaPxFvi/PAZdTJROLzSn1WDSW7OmS
9URaw+qmIoHgQeaQ2j9/yCJKQYqxV0BC3+MZJ1kw8nBTSEq/xXHZCVUxWxnalSd1
BMG4S5FkJJyQ4WyGhu8M0fmbN/TPQcKKTgrxmCCJtnjozPKqT80D5y3QkNNPYoit
Ry+UIAWJgRj9qKPgxq8GywfoRATW77R0bgtJ7Ztm5da7bLxUOB11ce4Mrh0WYyfX
oYkEJOn1WhxSq5ekPNxwFUEGbIPKPmTmZ6aIvNhBWCGwqwJv7jsPsmiPSfGsbbAr
UNLWWdxAehQh9h3C5ZXMz3y5AuYK+2QX9efbtHYv51It70xvWVDylMCDe5Ho+eDh
okJwWAjlJ0h1fQn8yhHanlZiBShFgFTdYWXmaliRmVSO38/Jzf2Xwdu2hkzO6kdN
4vFUQgRQ+h4PDZ7nxKUePPzITy8oNXieG399UDrV7/Q//XKPY9x9C8aGEHjLVZQb
nNOpr0JS5NapKWZIlKmfj3xvDMwZEK0bszPNbI8Yuia7Ghv0NLaE3mfEfYMFOznA
DkWFE2yUBAsgaVG28P0CphMeuj/QvUeql/ppVLK3aCr9BFOdC476upZnL/AiKaJB
i0Ln7Bcuj+dXOoQ6hqvlQrjV++gt4/iUDLDGN7uYA7/fTDZu6nuvZ8cWWgG0gcdu
c/kXvX4cKRTRkCL687T5GZOQSV2wzdeeehYZtzMwueDCMPXi6I0v5XXYL7SC30KV
evGgkyJqKSkv8ULcwsZPQOB36ekzOPmweF8GZEcJrCdGXd3qO4KETi7Hi0eLsDCq
SVn7FCHyRHIiH+bJIeiWmX4zZCu1pNbzyQ7q4JnSYfW0D5Hcr3v3aNiTkSPlTacw
AXGF6ZulPEUQVYWLYIKQsfxY7cvy3frfuYJXJSGrIF7st/7KCcbdupL5QnerHcX2
k/JJLPsKyEUP1ulfokYNEzesybmrUHpyfaauXB/fpk0mAgvCB83bdKykd5L6Yllq
yIlvEc1EKl5TFjCkoFnQ3m+jd7BoF1xwkoQxP/5xQIVWBTxJCStOQWmPpk/k+uVf
bvvO3kIj+t0U+NXr26hT9p6RAJpy4xtw6QWtCdLmiUEpQum0Qqz122s3iVMuhh09
Ke4mLYjrHJ70be7ODMGrPFxEVVUldjmQeDuEvBLNugNp0iG9IhbOscEkSH770XCm
fwej0Avcr3zAVZe7LD6xzKE7tMguW7VyaLRU51ANLi6s6c2mEx3Ii8WR3QHIW5tw
10rJjBLh0vjEf8vSPrAPzgpHQ+MZRizPgv6WinZZ+VErPMu0rWJFO/aAcHpY2i4l
sV03vP5eAiBIF0keZbAvSG/cBuzIVrpPsUdrWWLycTyVVVV/+d1KIhAZMrjOrvj0
AbnuRDt8X4SUU8Nzn9qrtm5KaUQtZaM7wIAo84X7/B3rySCI9cqQTw5aI3zx75Zx
XN+U/kYiZQpWGm1RJUi3SJhINsQjAPLKaMT+VGO5RdsrskCsQBTZWI1Naj1OgbLB
NPG75J6kBaS5Cgul28SlpC2fCwNsE4rr5jxMsgAlGrkgH7Y/rjJXDcXi483QuTT2
xqNi2QKd92yaMADbcKXZzhv3VXTN1y0Uw7yD/+i1C9vhGxYZnNuk+o/MQtSW4uWV
XGTH2OwYpLcOR1d2BPkNtg1wc42eaSJI0LX34lOrHgunPpjoIYxzxflrLMnhQkZn
9ij71wPEgPKf/4fjGFbcesk4pyYZZN46jOHmgJ4ec5Yt5I+Nyy8r/m/Y4cpxe1/T
B5J6FIlAxTUt1a1s62I784meEDUabVPA0d/fNiCPoJO09TcJ0h1rSLrKloyLZWzO
L1XCtCAV8JxLFqGTnoebJudUrIXEukw474+NpZQ8RKCllgqQgWfBfiSBhNgf1Voh
0xxtPPvAy010KGorIVjWfuz2AY8QuIJFRobxLfLmeQzSKnSPSvfVvCc4bR4vBLHO
UTbLnBIVH5VWeZFOrFh0buJ8w5pCGk5P6Ktb6N+R5okcYyWKWulwxs1SZe/eX7LP
JD7Zf6svLm1A3NvVgcz+HzO3GRnfQ4YtfARQfr33Vj2Y5zhXU+2VJqdQnp+jjU5N
2krCojx0MwUkBS6ytuAhObfmGHpkiP66lE72YlDpaJVSPC2heqmSed38Xk+Wb99e
kn9Zftlpk5E6HlNSysoQAouJ7959w6NOOQqfFKjIC8DpuPF8SQ949XnZUGXyyJNc
oUhZzJYDZc9R+M3FZhFrkoHFt5YyvAPG7j2jvYIw/QuAZ0cWGVK34dbiapF24oJu
syJ/T5EO668WbiXkg0GlkVna2xQbDtFFd2ROJVX7VHcrLonqZuytghRFx87TN654
WkPpMfMjdp6G6OnbUlHQPa/1Mgx0hGrZhyIReDr28FDwE+kbsBUXS9dXFLWm7ktE
dK2VnLiB0eK545C/fSsx3bAl0+x4Ha6KVM317+emTlbgezz4YnFR4X2Kwq42H5Uk
SpBVgQehB7D/G4c5v6++hayoKtRO6dNTjcGBuEtAb9uoJPGolE7bAaRzj6mw6VvG
4wXr3RNPHZkXaz+TkFPwXGstE2Uf5u7AaJ5o+WQyAP9JtdOmbb3cy/kkpCkd+K3z
EVxEqiDFmaTG9Q9VOFb7CMzZfd65azL/8bh20H5DtAYbBRTO+5ABhn5sOrxu50Ge
gPf0nASd1gDKoT5Wbd32VzLu5ZuwBnnjjYpExNEg5ww2k9Z7/3348275fjafiDFh
cPEqd/XSPoQgiKxOfEdJfnnbUMe5l6Sbk7WtU4WQIFTCiNrBsxZED+HUl7BUpyhM
/0/EkQr1gHBy4ojYf7a1oi3WZdQ27sJw2MD1udMMCVIn23pBTW/PXO3BYoCfgQpP
mwwZ3f+s01rUZR4JWcEU+fQ2n4KX2ONzwjhf+/Lwfz1q3KUc1NqODvLV/25cAKdj
xVFcx7J1bbtbu/VcDo/kXJGrNLH2zWAFdEwzcUOOzLwQi67x7ZP0mYQztkZT6C55
y1MiR4Wdo79v2XEiKbrWVS2d+zAEbP3r1lOjUA/K5AsyzGb3tKnklzNOGodqx5rT
07goJ1cO57R6v0xUDnscXyXxLAdoe+3kb7iIYVAPJtscL+iCTzBHz2LgJUiMsd+2
7aekr30tzZjvCmFj0CvR98+1IFAYnR+uJMskOmJ040A/BoWw3t8mLKZH33/B4I+A
7eyRjbCC558r6cHQgnc8oaWxOrXXufyCdzpB7D9gDQTv62M9e0cqbf9E6hhhPHN9
ppVDa+9RJUuXz4u6IpfCMzyHAhtYPNeFqxos5u3Ds/y7Mrgd87y9tOe64ijcyd6K
tzLqLKnR/n2Q9FK4KovsB/0Ksg4VI0xuyW1T0zunOfnR143ZnDN9pdlS13vZrQtr
x8/GPND6b/JrRJxbQnkgGDIfUF6Ys/pTX3di6uKu/ub57xuloRfjNp64dxoX1ZG0
JFoziVE1mHMX2D701I1fkr4WupD5dJ9iGD7HLWm4NxrPTyZ/JuszvVa++eVVOxWF
zj27LSIZG4gBDuzFCz1JcBPDSwNOffXLzmfDCpuxNJcS8VFnk3vd2/+dCEPJjw4C
xmD2XTTtlCaF34Mve5/nA5AsdtjsvHU7iOgEqL64TSLPUZBDa0ofEJFS2BpN7GGa
yynnYKr95+qWz8I5871RT+8bogY0+Jo65dxc0TDfz/ncjDqzl2V4avSNLihp/A26
9wd6chjucRVHDtbDfA52TnlgwxTLYTsbuv5e3pjs+c2fXZtU34pwPXEFA+E7t6Gp
VFBaQg/zmuj3Kn0aHqhfRUf7i0+sMSJWOgZ+l/wHjpAUqByAJUlsO4H4i9czDbGB
6O0VGu0g3zwqH0qr7FaghgznuvAIKXkA1hyPR58Oj5CAB0/D03SvbleOUiBueEDn
7CAwIebnXai80HFUI3hnd9r3z99cdt5EGexZpkzwattY+9upcniT4zrUWbG7hXMX
4pMrAZDaVk/lhKqoNH238YCo/wdZhdtofFkRY8NClxko7Aqr8Mi0qgLGfSHF/kvc
oztd/vCrlk1rrOfAAgWvAHX0fYzclvMs7s3dqQtonuE5SuuIal3BxFI34zL9T/Jn
wHfCCAtO9+0pz5Ombyyf4vZa4SyF0X/0S3DoXz+xfMDH1A1yFZIu/qdQVCZ8+Gv5
Ifwex7KgTCgg7EtoPqm4yENhm6huBatDt76+fXuVAyWWwoI3QODME1BFB3tFoUYS
ueoaCevCJ+Za4GbAt+IsOPN9vnrJQyd6Ty9JnPXZ0x8tvulcVbgG0FNYXzTjQu2P
ikwQ3O+8t9IYY89VHBMFGm1JWXsjBrvP+S8raifxZ00dVHb/sPe3CDYShZpXngts
/XeGXTtWb7bVRvz04WPKzwCqCix25z3krqsORzSaCD5HUIkMq5Hd+nQgMFULVNdr
Ednc/QnFbgM92fSK+ONgNM770B2Ap2X+lTbOCrAoYXg9agm+Fxans6+TXtYiICSn
19DGyTeeX+OR+MGi7sMSvy/H/BlV+8s4Ckdv4rVtYuPJYBNFqFsdJPktR2d5YdQe
4A6cykSBPIP/9a2B0/5SbtRiH8yS5D8sW//yK9dszoYRGGOMUnPIWyxNU7fzGpdl
G6o4wpZ0trzNla2WKBrd/vY59s5Twk4GWVHuEjw12YaoRNggmORJYZ6/tFKToTOY
1TCByIo/GQ+NoRAydBEPp9NmqRSY+b7X7uscUcas5VbE830t2wj39JZpGvGIxNUO
CaiINnv7K5/N+VaxI+UY+8PWNuRiRB/YhGfDfNeb1PUOMdgQnRTes0LWvd5Xi3zn
VygJF8BnHOczK3grBqQJnOwCSYWEKPt+Ey8vdd3GWK2+ACL7vKcfmejGA/VU2dOz
ILbLyZVz9WN2SKqhwDAyHIYKhf299/DyJjMkEs3vfJqxR3AdKDRW9w+gcfY226fu
xDUhsU1yai/Ln2SNtrOBh/ijBTAkOsTmzOsay/Sd1m57qbNchyrMtNk6pp3Z8YoO
rytuAkzub3XvVcp/xTLHhyzYY5Cx7SS/jFfX5hQq0scyzLjxN+F0vNj/Fwq6D3G2
Uhz5Li37RA7ZvVjrNVQdQBRhw+Mch/Cq9Fii/4K0Cyvzh44KNlP+9IuFwJBn2Rat
VXixzip3zlI6QjLjvlKgYO9H7BtAds1pOuCNjQ70GiqnjD10GQAJbptAv+ZRGrua
IZjPG97n85BTwfQdcLLByIFgfQnvjBv9NNEvKkTv2j/I0CxASeuV2le2yEF+Sf8D
1a+qfpuJECvt9oIG+2T6bWZNEdAMsaQ7UWwU/KkJuSDXJR52BsFyqaRgZr00tu1A
3WHZNG3BF4l53vRU8Uyn0egN3dJIg11jjb3V5eXiXmWX9aMKkNWUql+lzik5NURC
xyDTqV2hP98CYhk6KXfiQ4cpoIBDWKyyu/Cic/EuRIALTJwLL/FOBzVyPcl28K/+
fBY8uB46cAaS5ALW1rHEKSn1aiSmUPb8MefwbwB8WC5lV7I8JqXoncwry+EHUHI8
/jGG1CdyQw10zBHu6g9LDo94Uz7lG3SjmtonVHtbVwj524mStGdSav3ANDRndY3N
v8TLAlvZ0sLg0w5UKZ8zKzARDbFP4aLuUvesUyKqLQXmm053dr7s5WyTaT0zu0xp
3WsYz2xFrwdpZfv1nZRwVU1EMdjyUte4l/EvdJFMuTXsoFVIj+nR8VnRrn9Q5m/x
JMSVQJuqKqPS1g56fXQT2CQePCrVYjYNWVJOdbqbrQjQNtIXqqEancxhfVZZVPkK
0+QxYTi0VxmFPCP/vLLr7fuQIPWbzUdAtAzvxQGQx135mvXnr2yTt95Plx23hrvQ
RzI2QkjL6YGxcgM8vlKWI+cVsURUN7lovLwrKqUmUaYUWs3VEFMGhHyWZoM2y0k8
zX52h7bkVVc0IpcKV1Rq9bezKD84XPntjE8xzVHs4AYMiIpHPdTJH9J+0kw+dSAg
3o35xP66K8EnLHn+6Sm7NneUJ8iY7quqbkBOkdkzMBjHZX3k+dSTZEzkPNOh9tkG
gOKv3ZHWFY1sS5TFSzpKdwXfkPhi1hG9MmhRQzB0qpmYHtNep2wtzZZuG195W2yN
b16CMvCXNMcxXgeF22mx3r1tZOHz8OTotnwdapHGsWY9Ax7nhJ570vf1UG+IIUXN
AZ2LOlCEoXlPogDFw1uxwzt8ujjYelwB79vQM/eYHFdVN/Y08/Jrd1YSZFaMrwtP
GY+53cVQ2ip/D8L0if/YpHZntJ/5MpdsjkmJ8EYPTe7owqEVgSKNSF/I+IpXLKDe
Hr3IB36DUj5dRNTDFftluZZxLvy42h9WSBdIJUg+4z/cCrWaqpk3YKxQzdta3T9I
jA3qBW4IRKevriy0/cYFpOWdISCFW4J/kFCkxtrCXJpwDcBo1qyHvhWVBBRdkEyy
AWBr/iqygj0pK6H35q8tRpZc8Iet1eOJX0kwm1J7yR5QfE26tlQG8GkhVjHLg8+r
CET62HVv/4JMvvSN4WA0INVS8tmynZ1S6Dsy3YVhllK1HeGZothe+6DcJtiO8jgk
hNBv7+ZqrWSFzxHFZZGRyE/JTlhCLQPLNQP2Wo3SsaXQJUPFFzaAQD0V6tLF4BgB
dzWPdxFcsCVhzOJQopZZgTeDSbkzhhHTlIZ4BFUbDucyIJfvLb7kpGiIk+93Xo2l
/rRD5ccZ7P05YV5x3/4g0Qx3HoHvdhJXZ6oXKy6iO3aZVXtERdhgtxUmqV4gUUEu
zDszSwLo3ew44jyRtHlravF0+E/aYm1CG1ATwYSrF8ZCm+CXUqIA4URNdaOdsqNG
5626nZqv+1tphhxG5LPIWQNl5dwNXTS4LaPOKQNoKaF4FgEVYwdpzA8O0j+MEUAX
R+W5f6FBpeZrTVNTmoqmdJ5iAFzhLYuW2yvvZAaO8cplOp885reyrhqUkdHXh7H1
7qBtxBkh7jWOSbAGaZKzT4iY2ihxnEYkJN7EBD8T3SeRVBA25I/0SG/1JVl1C1uj
dAzdQeCx74WcQTum7iZmeC/6VWrfXgU4X5qi24nLYV6P/If2XZpWTgTelQz/Mkjd
ayRIEGNzghMLUjXwvJ8ldNPkYRy6IlJm1bUqJ3ZOpA5UlOiuTgiIgvBWjNYa8Hsj
TykcLBgHc4rrsw2J5J5kWQj7vKdefnOaFRFWIVYsXrWjtOFrLNxDuypdD0rq0WWz
CyIwZJ2+C22tTUGhw3EOUFkTEXpxBkhcx9pf2rTKP3S06i1l/HxypVBE4wb4D1so
Kqqvaib5zKlt/iQKwQ5ZQ8FlLmkWvaAqh6wmGsdTpQORHEYiffK9q2zYHbiBXYPv
alF6tvLAitu0TxjIt87hVCHLuTVWq/+EO35R4ZAGUmJRDWxOvmN1FSvMoLGuY/Ya
xjURHTvuCW09EhMvdq0es+DZXiV2XUXrv5MhmVFIs2fD38wUzm647J41aA00VSaL
7LPqRD6y3KoEXsvvbGxZeuC55qsMPOrStsibCWCu680wm4lSkx8zgKStiO54Ye82
7JylYkz0xtx39PeqIUo61ahRFwT83Mm6UcKVoZTvje831psiN7N2aueHGcqhN0cN
umryu8zFVwl6JxwzYOEchS8ZJZKNM2oIxhUSKM3pMWFy2h1IuG+Xo16aFXk2jmIO
MWAFKOz7k/v5JCy7nVEHkW+fCvA8pb4DbYtd2H3sq8mxhefNsK5E0uIXFpzsC/WY
W2W6u6Wb2Pz3KcTpxEoJMhTwylZCNuYhDPQukn92a23bc1ZNZ4a3fEttDeMGCXEA
/itNfgRmd4awE+srGjO5kJgyax/DQtX7YapIkjCJNMEyFi2d5sULNmwoMqWrPh0u
QlVw/EZkaVAGXZSdZ2LtUu74MTXU5/QSQGxiWkG14zqRKZi2s7BBL+l9bO2SCRaS
CNovpHSAR+N1qWda04baBDGpuMovfVwT3qlv2JD+Lpl3Aw55RAowGKUzJFyoBw5h
3dEK9I9gz+QI6J7JvlHa5Q/6bnwjNK+vdOpz6ORIZ6WgMk1q8IGVXYyTOg9z2ElM
UTCwkhwrFwDE+TznxMeXTxfXtxyKeuaf/d2Y3Xeo0wgE3wpAGQAnpAZMjac6rYP3
rxfWykzfmXJo/M5I/aqN4kPXCy0V/MoiCgBsWrOPYAhCR4YcPbZa04ay0mjxgXGG
EpkBMAsNqaNRSyzrcOAl20zh8K+1iBa1qhEna63Ce7FAWtnF6aLAfORoKaXunLt7
pCD6ir1SNtDFCB5VD7otpNVMLcw1nBeYnPUX71K855FfTiHkz+7efUDmsuajb8Wp
lc1oW4PeuE4IbEtl4DCjkpNLfEpmD0g8lvw+YDPa1ZTpjhV1bStkLgx609ARSp8d
CmQIX790358/q3c00uRTmWl1fqEzGxuKiHONYaxapih09XLhb7MThp4ZTyOpo853
vHxCm1qnXVxeTpltYLxyk80ovBAprXlQFT4C9OiY5zRjsW4swTe7UBSghuB3pGNn
5XjWE4aOi052U4SVvyL60Xf5QIQYX+gKGOBXCtBYdYxRlspXJmzWklkuP1uK696U
cqkhbpWeGyhS9zmjpztevi4ERTdvlcg85xzMxteqSmu8zT719sLRVMPZ131w/NYD
t3Qmie2s49ajsi9BzvjcQgCBUDvEXPx4rjawLbA1FzxbHfcjDM+wBLAhxQA/wJ0G
oLomZG30Kc1vbVbQPQZ5A9OiceuBw+hFpB666JgiAxUFFRhFzrH138YA1G7Q+Ae+
r3d/ctYYy1ifJDDe4jYSkHCmM2dX8xgb9Bx6MIXFSk7pval3JqD5+BA9oyRBmLtZ
wGkvcWyHvTApn61RzU4V+X4zydEXvwEHs7E53B8r8gbKc8Y9jWm6GkSvFye0tXxg
EGd0h+mLDJx/QtqGJ9QKEi9EqV+hrAtFr90fVFjGiHleoxhlFrunjkKVYc4pioBO
RFGQXAxqnM0NPsNCGz50MTIQTJhTyUCUJt/aDyxlzZc/nYNYGxiMDm/25Iv9lb5f
N8Ee9+/sJ516bp0Jd6intyqEBMdwxffwESvB2lYTFCOecL8m6EY92BrcoKb9hdXz
v2acwC9NZdRD8ZsKahTS51hxYFa+U4S/3pp5FkVi4Z7WRXHXkhBiMQmpB6c8rCw/
76ocYIDWOchpeRFe/Qt+Z5L7yEdPdSFCjjGCqtNJ14w0adZraLkaYy0raaLYa5EC
tdg5Q8Ax0CcPtgmq7yK73HMkidzMRpH4CsG69YLqongxc76G7tpEw1t8iLca60QY
/UfbOHdKopx1vNyQGEybCWswuOPD+4bIHUe737frPdDyvgRrQI+NA2EV/dTp6f2u
pLy6RrZPbPf7DXTgxEQaC46dvvlidzzSZQMcwbUEfWMFXGuhv2JBvZSxcl7bv+Z+
0xxb4U/Ei7Juiw8gL/m6E3JHCTc2hhdBf1Ea3HjLk/jyFpP7ymxxnLWk8sN17RtD
hOJCR8q/AKuBXR0pHBtgDaatI8n+qwHyCOzB71giNQVv5znZt8e01rV9rGRXf3Uy
DkZI/CrLCyOSzLd2P4wZD6x1BfQ0Wn+DMa25vzM/cZfhwdCuur4O9ozNYhERZTk0
DtB4MKTWCkhr3XvrhbQyjONf+RYR/vW8lfSpM5zQJHVv4WMqgLqdmMt11mWQzV2w
enpEcZQq+QjFPxhUo3y3eoZUHmDQfc0i6vAUZP6LyZPgL14we1WPa2F+glJl7qvR
KsmDOPhGGWKqQ8z8gTTvwluvY5VoAi2by6G9vKI3KhqWomXvlANwRvZ/HexGyJct
nEQsz4MNKLJ6b0G+La83rSx2hJdWH9U4Sd2KWyFmBycldOX8Da2GHqEUkBxxFrMI
+CaHLfsXIsfN1SrbXj8d9Sj5j/Qt2N/lDDzv6bN5X1nvGLKwT81JfUH2F0zEKTyP
A/P1QRQ8eMg2mebetMuzVstBA864l9fX6HzJfLUVCCIU6laDomyM+MAFxaCgxspp
O8Iy2ARHccQGpRmjZZmL1TDGVguAY0a27QyS+izTJ4OOrHOPWdyeE0kGkC0lvw69
2r7OLpZ7yeabZQGc6Bh3qywBszTsUeb3y38ncB6/wMeubduITMgaLy3NfGqsrDXU
ltxh6XPowjgbHAo399q7uYmOcVDYfS+TxaksJKzOM9Yox7U7eMEZcx7XnMFKCaU4
MOEwA9/vTd7ppx+CtB6bL/SKF9RmcHyvFUp4YjIzgjDuj7o17zdtrtFpza8RFkcW
+F2TzUAVYecWh2pGSx/tACPwAzWy0uLmsFSJdsn6FKDVLmcxdMsriPRoMCotC9N/
PoxBZhv6i/NppbQxnGkAY/7MtOekxmWyzvd4tNipkXXZ+D/2BfnfdT5VrfP6lJ4e
7Dr2s11RE9NMGfSW8ZWEdtVvc9N9o/Bl5aYyuhD1LCWL2H3JtwjBF9aLt9hsJN72
iapzn8HzE5IyUY+TomcJAD4NoKINN8cklAMLVBTiR7KBdaxteCuHjPN4emMl4OEE
u4lnaaeMgMAtwgdjZw52YiBhsk1JVre5J9BDUc5OiR3mWX6t7HMIt7t5+OgELnAl
G3u0TjFiSXxnz+4V6to6ssZBxL2mjCnMCau6OlyA3vaYrRZ5Z/Fv3YfySOy5fiLt
oKVecmyME4pOuRunXy/n6dvg7sDkCJoei7nsHvXfqW6dFrwTZ/bvl5BjQYJ2Xz/A
yO51aRPAYzDPKL1ufnElxm0kejtFJtkeusVQLXN2f0JYBJE9d+756nUBr8mHiP3B
r+ax7ErBrqbTHnp5JTLeMwHDhOpHEKfMOB3hlG9PYxHBsj2iucSl/NLfxkma747t
rnIsjuo7W88O1xlWaSgfVNC7uvwQXVK3r9SqfQlo69ys4UFLTddnWDRFnM2khDWi
pfaXnhBp3KW2CllfoaaXHL5gB3tP9XBhQi+eXh+yWMBEIbsuetIWja4wBv2edUtv
B0DQ0aBTAmealuyXi7DZOY6x7fQ8aOah0ojOHdRgoKcge/9zb3UUdztLQnK0SZde
KUTqHaeOwOlmk2qV/K+ZxCHc6GtF5LeqqbH9cLe6WgeV7kd4hyGvT/PTn3/VoIx4
aCNnLDM8DgNnvu+2HxX/+3hrbLci4CxcCPfQcXM6TNc5wH/CSN29q0EdrofVbZmz
E7gXuaRGFUhv87B4YcripAH77jeSRIegaxG09h8cBTZSJsz/fRaNW1T3dSl69jLz
hdb7D9tOzX2EKjsdEOrNznSD7SIyegH38stGDIy6W1bA2fnEwrKuNAci7etOWsrK
kamugpIazjGDWMRjBxt47DQDzKmOL3kG5MXz/iFrQm6ITPy6zbZb/Ku3RyYPBXcz
1EcEwufx/HTgnghiFZ83yHGY9XLb3jkk1L3CHYkl+y8iXNzrM+SZGqqwv7q3hTKH
hLY2lLp9m9SSHbJgNtDbEI7BvvZ/0id5xLaY7qke0Yf0b4gNGqOV6uIk1ouXRUeB
NlcotQHoBD+ijSyiLKAeGsP0mLl0m8d39NDSWnRXp/+YNO/U8b0BjflGrMtg99k3
LXQ49K9WVYXjQ2KZuIMDepfX4GbYaghYVEJ3zz6j9cHCn7MacJyeIuaKRRJp8q6P
C9T/zP/ZdOq3hJqXTURMteGzPG0dTsU8B2dqveBJyyMCchmiehCd3P0DyEUPDsMy
r2+0YjBfLXlKx9UWBMYK0/KO3na6NeEO1cytxQw40x43Zbdqn8dSMWYhkzkyIrB8
czTXmVnAH2HUQdos5rw3AR8z1YUpz63b4B9auhL9ibNNhTjc3VH1HMUi2V/nGBnY
nz21xMN44W4ycVv+jrHmwFsZaa/jmc3wUlZpI51zOOjarujz1PFyM0LT1Txs8AJu
SxwGunAnO3cWwxkmHJC7P2G0/ezIx+yRIgsSKC+4Z64Tj286PgqWGnaP+cZM/qA/
4Ep95q8OyK0SWg75CkVFP2tzv/e9w8BLlo6l2ThDXJkvJtx9Ij8d5kbxTjEuISht
TcOyqvjVN2NT3kUtUKtyoZ/DJEVnXbafqLuULkKPwKWQn4lT4JkiVq/SJNyFLb5q
s88ZhicF782mWrZEDkg326wc4Zp2U3lxG2lxU5nRXkaBePuUturTW+TeelUBlQ9w
D7mcPY+VWU05b7bqdWjaGdpwehN1A74EDjhaEiRCo+87g5rnwNpbUFbAsVCswWcv
+flwjIRgj3uIGO7CZtBLeBid2vWbVW85iRWmD/yTkXMe3VvLfVX6d05Fr5eRIuE9
wlVQslttRGHSr9r0+nJa1aJbka1e7s18zca3PzBEevYoxgUQFe2kzno6PmJ2xDCg
/HgvYB0z8VP8gvMMBsIE9r5IJ8vaWr+LdVvLt9IcZgBcBQwwmus79WQKqjr14Lrt
xkDHbgBFw84OsfX4r2h1KL4cBytY6sHkGKX9FpS7xqrCYsmucqXMsfN56LOFSiKC
bMFxI1YmGfUZZVJrUJ4i/ggU5pJdxWYxJnOXeGGFUer6suq/L0nA0yTtUdcR/XgC
ihVe3e/kQYKuxvUOqy/LZLkV++AO3asVkSyhI8dYLjz3HlKVZtM5xodhCVeIom+Y
bpIqpyahbUvD+qhhmpOeqpAUqT1h2Y4U0Gm3MVD1WZcUnJolwpHCusg6D8SVLyzI
Lv8TImJONAE7+1MhAhSzACGbQtWNeNnhFYFr/1ea6WBOZg3OiTmKcRWJLD9vAmN4
sdZdZ41cqsSR77UKyBi8ms0MDF7eRx3fKT1M4F2JqVG9lyT3b50wIxozYzmVxpQ9
aiEce1vtbaAU0f+WIFNuiLY3Xxv9bP6YGlta/XfhNPm3QQJv37fV+YGEPJrOUpeu
b/Ei64N/HLPMhV0khWL67V3OfcCZVTv0WsTZXSdsB+u/rCVg9LVimnb5BWF3pKP5
c/DKEY41GsURuWDIAA/eUMBsyGRbRL5qpm6HuPu0PeEd2MSaFz+o0mFtu+inZML0
jSCATf874SMzRYMXGbx0XVENJRt5ZSrKznA1dG19ou6SkKu5iEsGhTYXNSGpsDmm
i/NjHg8QdotcCIkeFDOdMOnSHdaj65m1xYypjae3onTWrWMBm97w344lnCWDXeHj
j01tsxoEcjvU3EodlCmUyeRTVZDYt15prhyBJ1UPzTS8ibKd5Nm4UaW7rJ38dg04
rBl5wGIECU3yA/Fq3tyJbmPQ5+KZQWcWxj7+7VC70Na/uB9wm0fokbeMCuWoiBhF
L7+9h4vrnTePf1KsWMWVGXsusiLhVcdrALZnT67crUcZzXMFKf8F0pLiZ8eQlfcy
7xrTJPv7PRfaiyqvPpLYiFtC0/yNFNqDudlxM5Lr+4QdRXEdx3PfdSCJk3cmPk+r
30mCi54HAYT+lxFAP2f0jizzeYYsB8KK9gbxcCstMoIVCYQsS3y/Qm0z1LupMw/z
WWmZ3y27kFMeSPScUHlp1bBLuykDAY0vnGXhpE0sFJCZa6q+vOR5KtOkUSkevV3K
fsodTVI57tpjLulAmdCvtoh17g7QaruojV2Q9u1fVgWKiU+fehJI/iQLO5jKfRZt
29bgWmoLeczU3lCNvYAWtpXQD/C7yZ7yZkHGQics8ByYKTXu6vmn22M2001Hk2+O
bIyDui+qep5zyrNlPS+RFYaKPsJkg/ioFSqFUT1x4SlVg07UR/JsCzlb1gpOPFKQ
NAKh8cenx4CDVPn/yEcZbIcLJkRoG0fBy38nxqeMspyrK78bxlt+HPI14pYYuANy
22Q5rdDyFh70TqWONLd5f3MbS/YH1bUPi+hVEF8J9E12I7AV1Xt4tyH3VMvq3aEg
3Eq39I1HUVKWN6WAWc2qnnnlhlRDyQ9oBZE8YiM/IjTpArK/UN8Mk4QDYKYl84l2
TpLgehrLmBm5LREItze/6ZVjXJkFD0SayCQbi0mUrW0+JGDatS5gYF58aPmdCwVs
iJyR3L61Rwq5crwW2YdEPWqFxood9VUnU0I8jCFldy8x4MDuiL/q1nPRTuW+ztm4
O0FgwEmSsOajpiJ7ETCY+EGqZhV/JetT9Sp+tdsTF+zbTSEzUEoh4l0aWkZqNQet
++Ff9WF2hBICMET7Hmq9sLGryo3gCJy8dJ8loNRhI96z+g0ikZRFGGhwIeiTXjzI
gn3Of3wqnDyWqOTwRZ84uwIcjm0gDi6YH89Zx1FMNGAZNq4SccrtweAB/R1AyWwZ
Uhe2OLjQnTyoA2vNhcG/16NEgoJp9CBG+4oJeW1/yUjopKkvtM4IhQR78c2AM9tB
4bp7YPPhbM25cU41HDI1PGAI1tJZp22T8ufk3SSxh+4K4w/tS0v3m/XgHYQjIWWr
OtvpUriY7PnbvwE6i9tCKF1MWAgnBL9BpoQ16yNQm77tA3z/4vG5bCFZLaW6Sk4L
MWGptxU5rEASM2Vc3L2dCNxzaACfx6a3hJu2OlALEG3zdy6lJYMGo4EYCEL+n6jT
v+9QJfM1Sk1UVl8eAF/30QNRYsuxreIcNR9tiLCSp7Uo0JNUQzbRzXrg8PvXa+Zq
C70ZwWlq8Q5NI+vs5wld3ehzT8SOuFsyub5NHFR/uCkIP1q6i7Fyd3U/7NAyYU21
BSnXcyCmob0Aqm2eY7fOtNLRTKW50o02Hg1Fc/meJLocvP/ZnRUx+VB+O5LJVtVH
dmGItFWk4u9dDb0OBuUjlRlu63N1RFZ7e0Z0OPuGWxEZ3jXyyCFctVItB9RuK1bI
prG04XyXtjpe2UpnE+24bxsRldgr/lTH+thh2xf8CsuZnOniNZgGoPpX1MF8a9DZ
J3KgLvJPNi4bVnB3yLkiO/p2LW9OGg8uaVLFMbaPTbhTcA7/0Wnv2WJS9iLuA+fI
LXBbDoAm2JZsZcvGiIJOwI6+widXL62CsobVu8KEOGr26N0olxD937ta2PTU0emo
8j1tETpA+iMVZ/HOqun2EYa+4SDdH+NGxOYPfuVmwHZmW7l4QjX8cr0rhmjWNEMz
V8rAgFONVA/9EPIg2Btr5VEa+WDsAwSUbHPk2fWWm95PBKlvVac7NeF7JCj21nY/
AxytC3Pbsy0nMlS+NjyXypySUjY8r+kZEiYcYNHZoDz/qPjiJcLwEkMtGFB9Pk7c
pSo7hLQP8MZcWMIuJxiulyTdQ/1Rb6oXmfZ7AY6AAqziUzKDRliztjIjIlNMnUEK
NwsiXvMbR1PTJ/fjeTxk/QMxjTyts46Qc5BufKqtulLHI7w/dVV5WDO3k2actUfQ
iuOF4j2N0O7+N3EfiMDJ0lfFjfD95LZWzS0PwyXuUBe022PA0/qehYDcPhQD8Rl/
mrB91aNL6kClxH0OJiS6Re6+ym1qBXP7DiGYf7lXiVKYdmsbq/ygN+1En1h+UFc5
EnQRzHkPQqL3obMO7eEvFwfOk3GfUHVMZcqmkAchV7nXavmZAOTy8Ewrabin2wpo
dO2xBsF0dmnuO5UsGWHUUcKEvVFChmhIgq1//h+6pC2a1/oWsWuaMI1pkOk92u3s
eiinTBfDNpI1ieo07BQJESIjA1x0dsqDtXMAbh1yfmOELRumBdadRZTfd4uerqWX
wFvrjLqwOtEmwL0I5Uiy37KsaqyVnxtZRS72otsP0oSm36cdALc0sz34yuxRCYoS
f7+5rlzGST/fkrMfVC9DbEXepEqj/5fxg7BygcDHB+oPT7QlOUfBNPtcNAFfFyWu
49TUXOGRkPLvrZOgNj/GTgf2E6rjZmxBltjDVfMadJmdfDr1suLuzkz+cOmXG7qZ
wFWcMoV87ILxr5BUSmW7HKtTisImbWlwLXkl5D05pkmEQdt0fi4YrZtKRrX3mouB
AvHs8D5VgTd8/qvdOcuiuUSdDFW35YsL1RH6tue5sVdqEWG2yi4XXe2Mm0r3rDiT
iYPq/y2YPZRkZoe32ELNAl184h9Fp5+Suo0rwYC8ALzK1gal9gCq2JyvbKPnjqL3
Qt364rHXJXKaNIT5h4Z8PG/VuMdXwr92va1IDGL3LXcweQkgzMc5edstLO6wsrXW
NuSk/k4L4lPxSqxouWcxrJ2GbG/2beOmXvZlJn1gYtFKnrP/XfE4CxKZx6zGVcDB
zA68Cug9AXEtJVYGteLGy+CzrUTsI+N/1mSdxZjG7nv/P0ZhThm2Ttoonci2TreL
P5pIHwiRRTbWpNrgrMgjeAox8taGkQs6eO8mzndqr0POtY/21jayWqb7LR8MGSOl
0GMCv5o42Ffag4vJBWWEeP7460vfQ7pc342okrGnWOLvEcaoLpcsKWYgVhit9qZ7
Ty1dhpO4xR9F6H+hNqxffd9ev5uNEwdb/EDfQ/tzh9NjLdqUk+6AYXS3LrTTEkgA
G7m6EcV4jfdMC1Q6VFid8/iMZJBdW/Gna8CYmZ7pRP+d4IsyjSQiLT50FVohQrJM
XzuzaRROx5m1kId1dQ0ciOWVCFrIKbUxuooXJpF8tU9oAMU3WKIS1A2f+p+Gfvpg
7efZsOtQIs2fH4muNLkb/JfVkLCJelRP9Yk6GD0jGHWnqxnUqiBZhP8DKpr/QIJf
Msuqc+CeXwy/j9bR9pr22WhVOttGKpWkMAgJY2/YBXu2mqAUoMBjSVLwT91M7oKm
mUVrWqLEWfCjMwEVa2Ovcflpz4yzUv8JCal1r7arLuMrPLUuQMDeVDMulJ070fu/
40uzNak03wzOFGwfURG8qH4fzAsigalQAyIZfuMW66Di2HuCWoxgtfw3iBhrAiAb
LVNTU7xFClAeUEQjeSDdCN5l09oTcqUQubvQBSJRCCoglu9sf44o5uFfHvnRAfI0
7a8nKkYchLAs1EgEfPv2dyCpZSuke3URjVQ+cVaIFbi7sE9CZxw9726Fy1NX1cvZ
/6etf/EZBiEr4H77/BhhWB44Y/2sG9QD3riRwOzYL8F19E48abTJpvclkVTjU4uZ
LHgntt3N0OGAZFxhKXa1HoaME/+mGG711ylYGXOFlTnb+RVVWiPUkfyDNwKy+bT9
K+iNPOeOiDEdt73GYCKqKWDUdu7GiTlN/BNBOIihq5OXuGo8vwOswbYgkkwyQU0u
X9UTatANyOXyg6CNV2kIFSJzl/36ztmym0g4cjts8dy7avvCna+bcQ/DS7r5osad
Dhzh7UeFd44vgNx5G1jiqG8bdrDyn3jJ5lkArDDVfRdBbgniCqo3bGqnlkz8lHXo
Ztb8+NR+kUidlL/CbvLB78n0YZSeowkXRJHcJ7DvUfYYMUi57vVc8OQVoum728gG
ryC4lldo7Shy/VsN6mouCuVXAZ/dgjCLcpmn+WpH2Cy+oOhzidT/f29JIqf4bO7/
BrHxKpew0DCns3g9DexcHMsLz1l5QxmqcOBoO0XL82zGCFdRH55+I2IUlsP6N0Cn
2tYKRvGT3mAOLtktO68x/aGGdsLLPxQyc0l1PJwHxZqvQs6uxyfJN7syrEiKYnCQ
82/LTJv0o5Fa6IgeDBti+OKs06SkOVclXqBNmYD5rgwqwJ6ZGE+JYdb0yG7SsXDJ
o4/tCx42hfq49GQzu+83hdC4Udugl9nevp9Dk9ky/YBZgYu5Gdjb+etdIhYhs6cG
QC01OVXaqUsw7sdD6J9GmCn8prtyPgejVpVvbHfxwfLtPVe0cwiEbuiJ7MtLZQXd
UDvE+5aR8KO57+wrTcgdhsu1PtLIVX2QV2S6wKiSlhEMX0aaeUfMv+i+r34dfUzp
Fcj9SGDpHCuse/FGmmiooRLUlU5SmyNQTD33uDJArjQMvzs2EZU8Ja0KNgyDfTtH
sEaCtUcpa0hrvDqtIFjo8oRxUthR8dt1m7UqfjXlE4UYB0fiOWPMEmyQRvlhVbkq
KEdRMpwWIil8w8mAKNSPNqy9+4gLwpJPa8tv+WD2Qj50W29lb2uWAbMoUXwzng/R
OKkHad96VTM4fRblcQpJpyONpT8T4PNc+pf2HAJK5evobXl5bTMT7mihjKGSPuMp
NZ1McoA3pa8bTepT0F5J+yC89xD3r5yxbDPo8I8xLH0YyfPd5dh3XT5m/L2Kle40
DMzGE/0PPedtAMMUlux40Oz+1QZ6Th81lkl8RSjcNK3PlWFkF83g/i1TDiUjeLcB
4BdhM1O6Qjhey9JLtVdjCjahlqgD80wSp/5hzuOjiLLoR0ASgXJWZAaPk99zA/yV
dEovgL5H8ieVVMkiaKUjt1XSVzdHM9E/v707htPs4gueMSjwpkw648s6qxeEPEgd
QWBZrH/X9J0E11OQzeFzs07EYdDYiOWrn3kHje9S/RtEjYwXD5eImLjUbnacQUEl
dl6rXvrYDEzlVI7b5Q23onASlQEvc8fFcegBxK6E+1WXSfqj1kX0DMHKBH/J2JEo
97RGKMNXwB6b9U6UxwFm04iktHukzfS/CGcknEJeEjcbezLo2wAOMo7PJvoIY5Hj
oip1agF+saIc0GVo0M/WKoUP/zi2ZDyvGFV/jvURuUScKAlzS76u4lDh9DkqpdEt
3iFhQd3dPu/ex0+E6NWYw4bhLdmGTvML5LSFvYfrGZK0vgfo4QF839tEjNyrZG0U
lsOixl1McN9iK3s6wJhOPI+iCZH1lkuVoG9T2J16lGqklcVs8eMpxE4l6Cm5hTNo
vFsGVQae3VIWXhs8tjL4HU4P1BDNY2dZPeZHZBVbyKtgZ4b+nvw35bTg1MTBlwAH
fD7U2uTK3duCxJEwIF0KfRWkxXSXZ5iQgzyPECzPsMM7gjG1JUxEPWWijg0kngIK
I0J24HTLwLS9wLazVcPkLzbcSJpaJ5qL5xzKfA8+osFIyTljacdiPggNg1fT/mjF
LWkNE8FPJZp95/fmbQfpLpo7yUSPmbhH/0ictutkVHtw5VLAOevCtw7/DSfONkm/
HuTsx/0GMqxYEocottNukemYLYuR9Shguwczidb+6gD+lWZOzfqD0utBgJ6d1rQZ
3ltIJAym8vcq18H8Jr3XKiwF836LDfkuEVXcmIUPBUxYkwi7COyvMeOfheOQP5i8
nqIFv3NBPQi/KtYTBiUuTH0gI4hMGyJ27U3E7nxau/eGuXzcpaohX0NTlCi1EF98
Stz3QiLFuyVD1k/r6sUkRioI3Pa+jXFUCFYRXtuU6+ZnJHrwqcwtl7/HwG/IqU45
DHe665Ovpj0EBMTKCpBauGG1EjQVp37z8stxNgZOvvh6L/MJcYcm242cCLhFlxPK
YBz1BAescGBXDmm/BXOTg9p7x5iJtlG0XC3ccTVLjhjs2mlMkUE0x2zZi/4pG4pB
vKkWIFodxYCsaxLatSZ0GfqpIhIRgiZjoTX3cU0B2kyQYKi/XZ6ys7edIbCYH8Gi
ZPJOCZCuUyK46xgnBgHzZVfFovzMdvgY2QtYU3H8ZLvN1pvGm375mv1rs16bNnQ2
ATz54uGr8Da+h2Pf2At1qLoH4InNHmOCQGpSXFpDDjUtpjl+VIqio9idXodj0Gv2
fkLWaF1u2I/lEWS9C2flfhDaQjTf3cRSsEdDBd4qf0bUmTddiY0ES8pljH8kiYcx
X+QJP4KZdP/fDpE4zYoKTVJ5hw3vQdzWZQiJxN9kar5pl3w6LAWnI7pbKd5NjpG2
AlUqPxfnzxsV2vOFm2Et73C/u+WYXPO81Seh0dlTCVN0tcasnaBSz7PoWcKHmivN
4Fvk69qBFW9supjX+cmM3XCtqX3bX2f71Vreah0Dox2oaVOpYSspjJyQIi5eSLez
PP3eZqgk0MB8wqvIrAZ4joa5VnXb4SDhy3Ilrorlizw/t9XdzJu3qMigiPMvAw1z
ik31kTWbX3D0UZZlZSnfITWFTnD6xAeAg9GFlJ08KHla02RBuwUZZEeF04RWPQJY
BSUJMzf4XGPGhjnC2khywMJ0fWed/uS64B2Iwk/plSDTft1hLxPyM5TgWSCx6+fY
iGLDl3jG5Ppw0dRx1x+PzVPNDFdJEKX8kGB+8RlDBZ1r3DhIjfGsQWft9CC1MwpC
U/WCQEfYQ9QuM5mGmeu7EEgnYgqtdbnh6Zh9VFne/gbadYOLRC19tF88BXuVMqx/
lNwjgSP3hd3E3KX3rY/JYfzkhM/bAKTyisNnCMF7O3LAZlWBZZ17nESroSp6kkK4
/lKkfMRaamgkKiXgI4MrZ1UZ1WZ/CVtVtsgULMvEgrMnHCcqfB0XzZcoseYt9H3g
mPP2sWUgK3jxwnF+hAuqYZ5wOLsOMHGHkNO2towrjXLgpm2ZLRGvWRjBrh8enOrB
dXF2BoI3TtqOsK5ZxRBFnpPnhbt9FKbUvMY7n02VZp2GVrgjV5Dxv3C6YGUpND8g
TFQtrVdd1aaf0Qn4ELenJ2cl/774BMGKoY4KZsUNW7iiaRpkA/ruoEKtKdpPfFSX
SB19SkU7P7EjnVb5OhoceDHRQX74Ik2IExCNSR1qG7gJZkKiUWqXOlHSm9Jgkacd
P+3QixsbOeVQjIoU6Iq3yuhGKCQG6vsiwJM3qwSELiAbdxAfzj3Q+LjERw5OQgRC
3tb2WqQfupVrwc7wiuroJVe7GNMZA8r/ue6rpHnL1MILa+JN9WGy5A2AKKZppux1
tQv6EgtSEt5OyUOtmCZqAcVwTTtA/arwM52FNoFiWL+tn9DKeOJIsgd85mSs8S5m
Exd7eu1kCwzloPy76jck/EI1zGfBnaNDh8SxPqsomYeDl+YbjlBsFk7CGNWCd7Qu
qfxbpdApAsPtJQxtlsdJ5J++5EGJ1eeRa4NTAasH+IXqe/wLxuEiqyQvrVQ5+uMN
k7diZs0UFxsuDwIlqdxHldlnuWkuSUgdDu69bK/cl2XDpIZXb6whVnSEt6TAqG0x
cyVG3lXVWNSMEuEn3zmvCIdAs8cB1TX+NrMrwXuSBDKKIb/bipw0ygwS7wSYeO0w
IadgB2ZUdRkodrdJl87IehkwkvxFfBsk9vej7Nr35hqAA0Ts8GZYDYrFNUtH6+ex
26MMCkvthq806lax3frAF2/3w52Lk7A6Xyo4qJBu/GoDdx2mMgJsqctY6k0zBE/p
BEUS/owwQF0XchrFIW4dF1azGvX1qochfAi4eCxK0lmdbIFalLAgkf+YhgL6O7a2
RxStVnuXSEce8ynVfRLQjCtnM/Oe+WXo+ERVOCUTQSY92SbD1Mz2ww8GeqF+p8Ph
p7cPSJbJpOknIHIc7e4tXKIifo+0+pD4wGTGb5izmmTUFbLcrw9LyltD4pMO1cxU
QlU4tlkvOAx2vSxQiJKCOmi2ICRI5TQ9GJbk43IH4I2O2AitrzdnkcepZtOBvtzz
UirzYtKg7FpNSU3k2hmP3IehAZ6n9c9M8tg792v8GnUsm6XRzC29ekiZWBlXYp0e
O1K/NmDDmLX00xdtJzASYR6efLyJnwHCZ+xFn8vLOuuqeUt23MCODd6o9UirByK4
Oa6j0D2/474hw6qYKf80mW74R+DHWJqLgw/mnAvAEP+lLneLsaP6JwwM/6qLo/6F
U8Q9Iw/5vw12VZ2b+ZXP4j1tif5akwLI+DFqLBHRLNJDPW1n0qooQ8qevfyOX/qo
bRSYpJk5oj3O2v101gXFaRtgy0INZnHIX3dqewXR4tMD5EWV7acHOL0syIQPmjhg
CpQpooWp43OO3P44z01XQ/XsZ87RxrOAoSpfSGQU/BUS1AzpeYunOtUpTVPaZB0M
RtoFiwn5o2HYhajXDPQwHyPs+QVVqkzhpV/YNytKxwdgnnQxXy51IE+fzxlvbPsx
oIYuUfUseAIFtBUWMPWjvUZFNL/kHniFDN/iu0N93JKAwxfG/Ncg9G8Nzgm3PvOe
GZXbbIoQqt3r7U2azfYPh5/WngDZ57XBjfYXoauRuFHO26MvxAk48+DqNJWBzYl4
kBJJ5KjQ7mHIhq9nmbHxMRutBzwePXppDJIIV7Dh1AAJMCc0Dsi8AshQcsO4nk/9
hxg0lAStKQGo6N3wMHVmWNnK8dubmbTaP1xkb0BALr//7jl5gm3sbt9N3JCrPQZm
hzU9eKGmE7lZhx/Gz8QZwfLl4h0CMjf9yIRFI7//JfC04/j0xgS5gd1mGV5gaatu
NSRJoZ9I8zxSbAh6PMaWoJOZbeHlH8Zcie6umPDVkSZptMEXqFvElApd5m3VVCee
h1oe/g5Afgf5HvEXOjd7jurmE6Q8Gz2hFQzJBR2sgH1OQRgH2rIzUVAI5HIWTC/A
3T+8CGpIsmbN0i8jveUdffowJZbOuaiZPCVjrbCHpUjIm0iBusOZEnGxdKC8tCn0
/egppZmBNMtdr5IHTwKsW69/+AeEw1fzX8PgvNBmhu8NgNpDWZlxjF/GIn0TiltL
MgErGV9S5A4RkVQMrQbt2VqZDEEQqCUJ8aeKDMhNrkiWde0h8TwhkJ7q+a3ayzWf
Ojy+e5340UeL2UH9odxytK2rCfNg9jGIF7NcngdBwl5H/qG/0ju1ZwNU6R9RhCWJ
vIZDZPUzoII7gMitmpwC1zrschzBc/SECMUD2oUsC0Dzt6bWrJdoLkYUTcCFNZyj
0/dFyjQJvqhYxSV0a7ixdHqFmj0ih0Xbg3M/z+NzcGqDMlbNz1auWxOmUkEQomqy
UxN/HxWdCfddf/02q7KeEE+pNf1Su7/XO8NY4twHegdYbKftVTy5fWexb6f7faAg
2+bbKqxj9qZs9wtoQteki8V1vLGfBR1IuOkI5qQw2LdQaW3MgehpsDIljYeEDxhI
H6vIu4Ux3WLdeibV+MLuFiCt13IlPefb+AE/qKRoRWGUf0jpwJl0bTN67tIfUUaL
m1e0uol1EIPX738WEbEX0gH+b6jdzdLGzw+Eff209TOGRDd3quGlBirVk5bJIHPr
u8HEZkSPHwavmySd2u/0iDN93INs6rl1dwwZdgX+cWCuz/T6u3wy9QIS2XwQVVI6
w4EWYc3V4hnlcTQcuXcgsBHTE5yfoyXoONYBIGpmaK3ZuvDE32rTYrxnn6qnPUXd
nQQ1TCkEqfz9G+t+7j6Y4KF9g+NQfk8QccDu//iNZXlzsoxJ8cH/+dT2CAJUu0Zy
1qVAbe9Y0JH5TqC0mpxEZ8eTHPi/SbQihEZOBwapYOf6fNYHXEJjGjolv6WOOcDJ
drkIKGGDvmqA6p54HoTXKNqYshXiosWD5FiMJ4M63Mur+484VmHKQKcGwH3HUmd6
+wwKDZlSuytVQXZE3myXZCKzXMXWzeCkCBW+mo20l8SA1Y7dpSZzdHIRwiriL8xf
PqhtQ7OeUT7f1wpU9FbbFPHP6DF7oUyGvGXfS1RNlqL4Q9BO/2ocVV3qvFYO2rUB
JnW/ZEt4ByHQex+JSAvL7mu2PP6vxcTy6HlVCBL/7eTMWDpqF6r4etkFnkMFjnho
f2v2ll2I/r04EEUSo92gIpeuqy/ndmH/XpVaeaL9e0WEvwCejjlejsbD5xvhG6bn
MVkL9I0MwoNFJx5OsgH6O8BF4McLMtQ5mjFPZpdHVwgFdHFz0kZw/NXMurtnDXqP
Xm5OOTGgrKyPp5wH/VdoXro28lZE5ddU/EUKZC0Xvqi9Lkvg9mKXMKJi7o38Fvdq
wCuVR6Lm41lWKNjaAwb4RLI27Qh7rCpu9kpz8TBiOB5eVeYFtC8flwoTXA6M8NQd
eD/lrjpYBennNsAYWxxzetAYNa6H6dx2dulx9oeNX9e98XCsayY56AJ/6hBMYxWl
JttpBGoLT60fZPqsb+7Y7gA75agsh1J1bibDdjp+j9OnOB5pSsySSd6QG87euCY1
/NPJzKqtU5HiCRA8cGr4elMhlCqmKYcRG5GKy+OtWW2tIPY6jyWSfpLx2+Vhlw0d
lTWt4sD0kFGwGxSx0/MvC+qi56mNxNv1a9YQGnMg/4xXJrP+6+8CROh/8fSTcVa3
yA9PWPoRyqRhz5qKV2MbDFR+kvthD8rhu3dkJQrPrfmi0xJfYP2NC/YYrewv4Yyj
UAxNC0MeM50ecfdnkpXp8SzJTvPBlC2MArnKlsJ7BHKPtBBxHNL3qz7UwPnRk2P6
EAK9HzGaXosXB6Z3Md4YqhHE/CywOn6VEG/QFBRVOT1goxsU35EStWB63HwcBtcy
nB3CFXWWQKZrHc6N+AYwuEtT6LY3GDApw2K3ePTpOPnfa12h4m5kLndAmKaUlFn6
SIBO0Em1NdL41wcaOMZQdl/HfwlIU5cSmlnvRH5SiNM51gCUFaKvLHN0pRe1aqRP
y4/VLPpis/alBNcA5k1nI5P5pcLgW1C9IAWntKEkG+1ddCi8n3ag3WFNTPq+Zf6N
Hyvnct1bAD5GahjJkXvnMj8zI1ga24/UBTrDe+wwtg/JZMSIT/CYqVhKKOTZfZHG
G7ZMwrZTBk+z9x7Igldq2JALkw6YBmxVSAHUGcmJhso7Oq1LyJEwlmRFnXoNbkeD
afHV16drcc7xdNSDzYKhwn2KNu7lqJiycMkYPTT1ElOZYqCxv5UYdvN/CHu3k11k
j+AQkyCAySeLlY/izTOz0Ha0v8g8sYKW8h4gTrQhkU88sdAWVSMvtXHFU/65svvy
w++ZpUmstirjaHnxHAemOfby6T4yXchQ7KCenJounKhOH8TNtEPlDzJnXqPAa8iK
+lb3I7vvbs/EhIZB3sCrVB1nmAJDL5M74cJ6/a/c70DmT5iF/mz6AHOkXDkBg/Br
bYYmANcYfxdx63ZFgGlfPakKxLLLsRu014WksqZCFuwuexMHz1Y1dtdIgV/rbYBx
VseLDGjLuwpqy9KkRA2cAyHv9W+cW+oJLA2dweXgc7MZpo/FC7mz8h1xQW7/G2DR
/MNCYGcuieSkSrjdLTVsDAnxvzGXA+JqdWEHqw/FBDDWgoYsBg3PpbCxoOyORc2v
ImVoB9bS3R3cFcfHNfAsWHfdhfFCVm5ZNGpXz55WbPvg0aLEVskwN3gA/1VSwCFP
fFx36zpfWz/+6iXVXhHPpIwKYFLsHAgmSeUEgn0WOFczBSewTHG7FM/HibZdvtaZ
s2v8X3KRiKbNG66TIAqDT7mKk9F/w68d9oB6+AvhIEwoYSXG6kFOpQ4P0DqJRqwc
X7xPUKkAY9N6YN8DGrFuWRxGcyzEYfNUcK3pDRQTSZfciAuEI+w8ORaqGu6HQjNM
to+pS8Ja2nHXxNpOjmrT3Cboz/74YBs6mNvWoY+v5BpnVCTQxYL/n7eyONU83MEF
HNX4H0jXpe3xSobATRmsln6VLDb7dIblrNZS6L35ZBR11QI6CewiBGN5DaaH0Wab
EH1Qw5KGFPNvdeBKEXssEE+BbLf/jE2mvxHvoq06Az74eVA6uTZDrYz8uGSmey0P
/hdXdFD1DGKKtv/p1SotX35zH5P+mkPc8FsnJ+LYLZuMauWld/VQSqkXjFMzoCCV
AoTNiFimGMK40r1/fljkiw7nxtwwuB4Uf0upKmqRVTs4+mHOXkom0OkgYY26EJLe
kKOYf+DqkGf6Dh4vQ6pSBtZ51YxGRMW6h+pkLRdCfZammusYSSNkn/mAupjZaZkc
7k3dNECPkUCAYkmD/rQmeXLuEO5Q91E+y3gGWq4NFL2Qyx+hGKWBncdt9Z5VDeyP
Wxju/1Dsr5JVin9+I8Sye0s+tP079GJEBBPEoQl7IVJBrWqSJe6R82MRIrx//9JO
KjRKUD9H4grDC2Nmy+vSOlGsUiMw7vP4dHu1ltuxnbz87sCtk0RQKuxXISyLZ87N
LllCbhKpuZoCUeHdDiUWaN/M+0hmI/YWKig9CH0ymo698oWPDVb/OAHrpoVj1zdc
3daPA6wH1ggbtHtS5vTjvWCbC89Mxka7ndm1q0jGijYdLFgEEEtcEJIdOCfzudPW
cyD9Vj9m02UdI9aT63XRpr8/l+QsEbRuckKKfUTtOJbchR+xWBlT8Ld1gNlTTHvf
YykFihPA7qvl3rbZmjclILNa/p85p140dCAAyqAHt3NvF0UYlwSC04K/5D9Leeoo
10kY6ecnjRAyzZgeA2EtN4lY5JiYhoL3QJE/U+b4HQYzVbWiQB9aQrK9aiAq0Rgm
3zbuFycoeCfB2XHG9S6k3XU1WCClbUU0KXTwsq5vazFG3/oRcEAnTd0Sp5QWNAiE
DkaBTFpT3LnNdRXLjL6Wyob0CttBOY2dNO7YPcuvOJAiKKK4L7zO8GQb5p2qI3RQ
iSRTYcfaWF2LVPUoJrIgFiZf/6rTa8WuIvBQGMK0pD28A9R9GWlmKJ9SyrS/xTG0
HVxk1AS4vC0/0W0AJNLBKo7+pFkppg3KZSsPVdCbD2ZLiutD0qLW484xOdf9okTb
5/XaUCbnPn0eqacdA2cLnOFvB92CrqWV3BLN4YXTmd+a56bzJcz+2TKf+TfJnbEt
Z/own+XJ+Ajf6JT1fUIuNrxBj6TVtkHPa0DwzRoTF6hI7jziuQmUndXnNH7I3Ur3
whZ3rrOT6Y0OlMcKQuZrNKLAxHEI7pnbD5XpGVHaz/yZDx/GNjQ/4HKzss09bAYc
OSctB8za1aHJdlkI4qMGibdyLH8vpej0rnEZvbpvZ67YwmuJgEAGZo/1+ze54rF0
uko/DN4TYgRzaOUnhd8PyPvcW3P/Rwv5uHhZWhMx4q+c6JhLB3RsDeoFXwXDhpaw
5hKN/sy4EHp1JCdR7T/IWaZjJaQ8ZdK3QbBQKNnDq08ZjjK/23Skzg/ZM0MrztfT
O1vZkM0YO97JnHiBLRidNsbxm6AsRI8Gx60me0+NCW1VCJYJg8QMfMGE2gVKrtZz
5ceAKUOAaG9xn6KLmG3tACewr/QbjavpgcLslWIQnv0XotII8/uh+FEHhWYAz11X
PymGybXfiR1Xqqv105JOwB9qDJcoFDiGZ+LGPzFiwe35fex45eIjKn906hFOBPOC
T9BGh74XqLHmNlBzXh9bABHFYm/RrAKDImtrV1vhz3gv47QYnGMyXhybg7uPZxqc
twlx+sdtxlS9ZjsRPgygvPRgLzfbvLDzeZX97qgyRwsYy89gswekCbzQAzQH0N6k
tMsrYVWvHBuIS1IyYmbOaRSHMJLahmJTATBpl3OOnKRWG3XnMHMMzP4rwuJmSfm1
MZTjz7F2mpGnhv6R8W9OTROSsuk+5FEaeHzq4Ww0/wX8XzM0hGlBrPBkYSstWgnw
xJqy+P1EFqUc2n5AVXgskRz+RJdfXP+i8T/dLsNVSoc2qtpyDmKIbNKwJcV/HIwq
rH2Yagv8LWVcBD/K7RPH5Hg8XQYLNzxTYAo6HwWIxh8b68/DOU+80oNGErnBEQrb
lYBFNhyMS+JYcMyyaWyW91A2tuqXcAgNekfdawzmeBsv9nFtjujNcN1BfV6Lag87
7MzMpmFK56g7lMhRNEg7EDUk29WfCdKseipPjn9DnQjgIMMVQw6xr/eirfcZTIC6
KIQQvEJBqCyaUM7z5lG2drORbEJnZAV++4V7Wn4+h0fbwVYTgwlCbVTYCQrxVbYl
fcrbS0FHzjvX1Ab0Im1BikeW5DIfzB+eQkmMfGnV0LnxVs8i0FEskeiQC94GQVLL
uiG/+X8+U7UmDENIwCPHxjU8uOFZn70NEX78+ex+vBHGfwKzMTCitROXCZZ3mrJq
gtrRkpulVrVp+CEIXX7Ovsx8Age2+WPWk73RATCC6fR6mAU1919Q/w4D55MXIzfa
UAoxfwsMAy6Khv3nj6/BjB+0ex7i2tlfbiHFz+jt0N3aoGMW0yp1SX4LAsleiF20
MbRMnoXzBjZID68psxE6ZpVyggwRf7OJ0zx5w2wpiJqfL2MWsJ/NItq9sTDeqYgs
ikONIzESvwCrR53zxTQk3Chpp+dm/pckpoxTXic/D2YalRWkYNpvsg9NZ62E+6Vv
OZ1ZKcycBuNfJmKB9+rwZ5F+0v+JdXa4fdA6FLcw6LCE9eFYHzbN9PlpyGH+VjiF
JPJKh5/LeicI8DmYmgQzm+WulEcYNpT023gl2+kMmWj1KFU2sA749rG9HteHGfh+
J7LXCzMWctyOTidRm8kFMKR6g2TKkw4kP81bJk9buwfL9LuSQE3Mg5dA4oEMvyzs
XB7qCgBWmq2ruv/Gv5ssJU80nwBEmEUrh56w+3Kmj4BpvE7uUoR+PLc6YExZeaEj
ShihKKm0m3XIErsjZ8X7UXeDJiIvwczSoxnwudtnJxqztrRTuSadPgoZf+X+NWRd
MR2QxVR+C3rlzUGtV4w8VV7ApdrdDhQnDRHLfnG9D73I1uZYsXne07AtMpFv4nV6
rP+47c62fsr9IvMtWUfnoNNr+Ge+crSxpIHujaQfCH56G7BP4DEC5i5CH5cW6RMv
iFrXxirKodJQE3KMxQqziQZ6cf3oxnPBZ3spWxx/0BLFP7O9GjIvuZnSmGNYqXOu
p7E6gZ1ViUp7kuMXWc7UaNRivygxlzmJaVXrjZN6000S+PoMf/qODvw9pdzidtaR
YkjDtcr8YHTV4ESKcfCquEvVibk1NdfbQ5S+RhhfIgyi1q3i8liRUKG7ZPlspoNW
VMIVWTbVqsSIh59CrEJD5AbFabOhqY5QI33cDNgKVHgW2THotNGIvWzY5nFzW7sj
Qad2ZO3+G5OMkNokkrp6qsYdUvm/VacgqPEuekTCGNYT+cyxoOoT7s2//zfVbE2J
tde+5dj5OEUDdYqEtgIg8pqoppPTDcDIrSY9c95NBB/e/zCdgg0tyrG4ei9eoCjD
iFNBBCmBFRWZbjoxg9CIk5kOOxSV/NCSr6oyLJlgxi0rdjQmzFFTqMyi2IDI9zs7
y+RIqBFZmZ7DE199cLs/Rwzm6CuN9fOeQr6n3LzsQq5EfKpLA60azwR27O+IZJRM
Nh9HZnDeLih9nnk3DecEi3QNplm7XoNHlZ+uK4rk+nWxdT/mXZWm8g1ji56LzRVJ
3a5uD+7QuH3TT342DymXjfFw6hfjO3efi+W4yy6uC+YQQTQ9j0LcASHbcXxxlQ6u
BgtWyTXMnoo3II8DFnomiXIikvcIoTtcIQoUCT5NK/s3vFChiPlNFQjacw+gsrmQ
yc7xe+q/tOgT4FhES0nrL/UU0FD9TKVC6TnvOhZ41seiA6HJiLrGfGxl9on40sKa
Canun5qNYTQb46ZRHRjJ0WYMAyb9FmWtIvIes6EMylprZr0yhMNK8m1RXA5iYULe
V/aYVmZ2v2Wz3LNQ6t8/ASOpi+g9aUtg5xMwY2ZhOJX7VgTwAE1DxM7afHYwDpnc
8APAdR0fX+BvsxvjbaZjVWLc8jGxYM+7FEf0pyCebKsrW7AeUiRg4PAI9ji1booc
44FJMafmflU2Rdk+l2tEpZtE850RffGTQa/k4J5OoZF+VatBFGF+/PT8ajb/L3dJ
u9ZJAua2hf3v+BXNZNt49XdfDN3hEepyxssJKGcJpz5/7IC8gM65lDYZnKDmC3K+
vGfWv89LjaQVwIERfLTKYtAVU+0Q5rP/xsARiPR3IppHiuMnh78mNa81DdCetKI1
Var4o2Bzw/emr6w7fzEJ08aLoUkJGVbsbVBW+tm5Nnvyycbdtyr/cxv5E6Fn3ors
toZ4g3YQjTaS6w3n+wIjxzeSlfEl1m+D61nvdGyxW1VSb4ZBYZC/2QsIoicZxV7l
hBz1hD4JFWNLIJ6uRyE4jmamTatlTxxC01FkJFB/Cb76vFyOiJwxZCbFT4Fviqgq
zyC3+HuvsNojs9x17EXdFCEBCRgbSKYYmpN/XNVOBe0/9aZX5tFMMu+PtzBv/3sR
TEdCEO2afuFT+7GbDTwQHpLi9ADeAPauTNusXjwGW+GCpy2m+EpzmUKgbSaVnY/f
aHl02Ysp79dX2U+lGWDubx9/n8K2+dF1PXh/H5lxEfmWtoNs1hVDcfOwgQoPofsO
hJv9S/dRxZjvhccvNmJhFyr0vWPiJa09X9VTIkagVmTYbzJ9k+fCbPCGSRP+WmQz
WlN755mIH1DB9ZO9xR4xIX9CWIuniVb91lvvr8teLgarT84vqAELK/IPoh4MWu9m
RM/r7qNYzMrEPl6/fhMz3ttsLC9x4qJgwOZIji0OMa93Js7bZ9xjDvisjzPmW6iT
mqJkpLXzhWebiIk+4GCPYtOO4xCvWXAmb3yaMWp86Y3JZ5DD0LCEq6E1Pruij+am
sQS9LMsdqMOImmjGE8JSEu2EOMqAP/M48jA0CNOaYmZiVTNFQNBpDF+xmwQzfYoX
b10yQ0RkakXQtbFDfOI3B5bhuqEBbes+9/s11GlXbQ0zicB2OHES/LjQH+nxgjQZ
oNXjroC72aHI2l7ujRn6KOUcJO7OFeQ1HD0aO28kPM+NszCBhWuI+DVEEnCKmdLk
c/0UoLHFkR+irBJkAiXnM6nvWk52tC1LcbtKI3sQDL5ny2K52Bi3/n0ZHlwti0U7
vcXHmuBRLABSRZGiSI8D2csjEPij2/vDJaFKa9A8DzwLPbcXp9apHwR537TDIc1O
1iDCFxZUxbZ0EmJZC7sg58p6RNYe0u1Zd1mXZT6gun/RTRT4MgfE6X/lyeKk3Xw/
QGBhtQSclsbW5IdiQvj2PIps2yyuYk7KvgPaVSCj8z+VcFvTTmRrHDQtc/agJGUx
cZDEP8szyUa8hKzsk1Cj2zVHjh+qa7gQERytZBC9CNCW6PPTUqE4UgSrolpOC7hj
i1fkmhxAQ60feU33kOUn/V/JwMAXZE/NigdAbBAa+hM4G5rAC/w07amCWv1S6ilt
LjTyrJIggWdtGdNwk5c/sWTA1VTuFHcEXyvqauwp2L7XsMwCP1lvfFh9CUqTz/lU
7MIUSCOMrD1dNfX5CDns7tWA8DdTanRWvBUinW6u8rmn9mAB1f6zQGGEt1eCkDas
xXmrUGpDcxFihCrIGFay4d4W1PbM9cxtDpF1Siiw6qLvN+16E0NnjfSEsPjMyrCV
JdNI6ixOnanNWpMNQz57kTnwDGgCVaJGS2u9Lgy5+NkpnciLMnPBUtjGLdZti4cg
pi8i+GJAeO12wSq3MoOKpNMTMiPeLBGxWQVhwLEaLIsFnhvc9/qC9tCKBt8bhsxS
3ccVt092utjlXALt32LF9BFOGjbfjbUy4Ic98W3eGulftXwEJnr4IGtudkCwLXiF
Tqj14yU/H3uFJlfouE8jA3FnZGNdbcEJFfS5ppUYZm0zI2fScTBUv7A3W64etH4R
2s3FTyUhUme8X13ygfbL7wXx7DpKwjI9AbG9xkFTzymhpMOq+yzhhLbaYBQoiRQt
CdZ1J7Wb6Tg/drg9b670ggr5jmel3u1p/g8brsJzwSy024EyFV2dIKD0taj1jvO2
8me+AP2ZS5KcN4EidurOUh8P5fxlvJaLzKj/XJPLRGQOBjRZzas/sCZSLsP209is
dcaZjSZgn0An8+OXyBZDYnHVNkT2sCHPD58+EIJchRcmbeNbVyRoOduBvpFgdeGr
rEWU/sVkC/jQUYh64rCzMMJ/51tBrwN13LiToTHkNIouVSqKSPF4Oenrjdb9pw77
cXyW02VtkjXXcZ8XgyD2ktaMoegNmJhUIjIPmIyfS9OwAqqWfOTaHifHikcPuyaj
WaTafbykLkD3pHspSDDcExXXp8SmpdlerI7W79Vz01ncV6YPMbqKzosD3LIhFryA
nZMwa2WOtfn4Jt2x+YXjdV6UXIY31OuakO/FioBR2H2aYN+oo6Gf2iVns4ZmkzBJ
DVY2Lfo6xhHn0dSvIoIuJO3Sveyr1mhXnKRQeU+Ybl/YCr08cVqKDlzoUuuBUWod
EWUj4eiMxON4Q7Sj4dBQg2j6Zgd6ZG7yFdYbU8n1dBQcGuqaAi5oshweeCZdRxk1
Ygjc96aAPzRm0MPKq0waQU4JFqkvkb1L3PElSCLpf//28QvPrQH9r1mHNGsLj8gy
L5PVT0awCHci1y54lgWXdgUwlSXvk3xGbP1DB8D+WjcC12EFe/LfTX+/9QWDev3z
8ft7A4fCzQRsegeEeUPZ+dvS5wtcsZudS1AjBDY+p0aP6fPnYqNXQdKRaWw3Vj8S
yZ8Xi0jKyZJQF4G2N1d37ZnvD4PYnJQFScQ2lXOmQLnrK4hGCWhKWpCATq/SwctA
eJTnqbUw85ICxMrlPqhkycG1yhKt2iNaDwXUENobCw0JIvSMI1KkSW4H7hjZTEo0
nQAIztVNIMTfvAuAM0fUmJmjDh5bFQ+pb+7qUzfzvHxms17jlJzyCaLPXy3uFwOy
tVt6UuowoSc/CTkJGfANUzXDgHqOuFrZmPAUlMzCSCTLclK6OL9diDvl6+vIX6PT
T46nQxmSMSnqKosupX1tEmlZq0V8T3cY1JPt8Z91u6ejDUpHoDTTxh6JxgQhg74m
cABXZpiunsT4Pie3SGOMzjAtfMVQnm/FjturmchsU7wwBLhETskyfUrmNLNL4Wyd
iD3qpWWeruaumKJlRJ6Gp2D9+fswstzUPLW/AkaNCX7ThiJ4bH9J3sf43Vg6e1lv
+R7rKnRzDZGY9knDWgIGoJOIG26b6aUmf2clyrSMaODGpC3Toe7MC/gc1/WFUZmC
m5oyn6e5eYAnmza1fKx4qyPsDSiaLLeCE3ZJkRlco2ZlGARGSTJra3jA5AFHiblj
jDEVuni7BZ3RxCXqiibvOjtyU2N7fwxAkW4zy47nHG1YG6HEHu9S/tIghYcW17Ok
KOpVxcGRwUCUP1ABnHToZJxaeiuIa8Ajxx8MCMQEfb3lTMtzpqg2Lp+YgZMmc7eM
oGfVMt2ylid5n7i2ZNEK6600pvknHcd+DYlrvN0jvqfp/3bu9JuG7XaKlQuJtNwD
tKfLqWd8iaqzhlz1+6x1PGEscVWz88jv3HMwdPQF0LdvpABfeGQg3VdmRdKrtWhw
/wQUq6tfIzwUCX4aEbwntYjxQ8z8UseqxJiR4e5sBQlwb+PcjhOuM7rSd5wcbWv/
bMdGI09huXXXr1YkxeQF2Zir8P5AmS+hlRPZRrYYvm+nsJa6ykr8a+pujg9UyI5E
XT0qHwho0tVlzpMc+tTu+aqmWcK+hO+djTacToxb/e5NfgNrVz0dTsG7U7cRe3G6
Nl3GJP9x6L8JzaWuW7t42O5xje725YZOoKoMo1AvJ0vAs/iTXq6u3OXt21+Bu6Ez
XCn/20v3x2T2B4Om9kIzw1y50xFXT99V+rjJsCmf2+e27jbAJRD7Aj6Ui25X+UzD
4WiJPxRQ/wDdnEmuGoGO2dYhkE+wVz9s1QAGBwknlfPutLJxlPQVQN+sPs+yw3pf
WWFBn+yTKlVSXmMEdhMQnKmfnRLBSnEfZVyVD0ErEJ7QZmZ29yjKk+/XY7SH54l9
gLuW2FH3WdtNxgeHlW5UD1UR9wIzdFmkEFdwbodYgh/VTtUiZRMmbGAdBSPHQMA1
7YnFdVplDow0riQWR35Fuyfc3tVGCVkr/kY8GfJvZjhjPpbRs5iJIKZNy3Jv7Mm+
AUUuPIpZB38uQ3BC0w6hLxmkjPqlwGuXT7c9RZhsW5PvTjbyItcMA6L4XOwwiWZp
8d1Fmof+aIVNeQRWPSPTvTY78oySaJFyziKDoPQ7Fyn3uoAXllwUGOjmyAqI1Ben
vP/PMJUaYTf0nT6Ev/qxQbQOHiQJreNr+uhAwviYFoOYFBGORHxqGLWg8iA/yl9M
3NKoGvh8otSVGuRrWwZQgCOC4dPOvSehkpX5Yc7Kyg+5HIG+1PVbbPSvFabvsWZN
OiEp4XvymSzPwHwx4WvOeX2ILVYftyHqVS0kfz2FWizunJNKpcZoBkxygES2/k5Y
9CwjNrzLgbb/6rjbtvQuVDR0fplpMBhnUVSEVTArYbD1XispjM5TeXLYwlaZocda
zqVWuMGE0FRAmrVyvYzaxxKzNFT10MgzY4G5v7jEQbihkJ9hULOqFcWGVsvgwyVp
/ZuDUjFFQS0JVh8nKhnNIcGQjRazUtdsNjbTX5zmjmGX/eA6cV9agnMQeUbZqwOL
O1l+TK8AWXhc8a1T8WP+oXxnZ9/vHlzwUJFzasOBJYcTasaiwSyGP0qeFc2C8ZCx
8TquKPtORVkqE6FqamOuXyZ/BrSPA1J+p8IHfoGH7PdKF6Lzb+SnoP+h9sZZ0puC
szjaa+XypZMOqZZo4OuY9wijmDwpbcjVcUjTjX+tEK718oZUKfN6TvbzzFP0Y3TS
I2T4TnjMx1ybyDOz7hgKXW9d7ItN3bXrlSqd8YO/Emd98pqf29n29G99PMliZzpl
MnJ0nbCs+xGBRWp076w1UtH4OMe4Y6jYLh6nxMZGgZIfRkARz4I+65pKiGeSesAB
uveejJBsqKyOyYc9wmu+FxrxS7DozREOpgiuP+fF/1OU/vFHpwWPltVw0lIUb8h2
bgq14YUPnKAygq/jpa3WKbY4hs7snsYZIHytVW3wQhdNo+gGh03g/jUoia0QkYwR
YriAoSji0m/uBQuFRRoeKpJlVEy9BvhTLi8tnsFpGp9w3s4UWW6lrdAWC6K6UoA4
Gn0a2jJIl7FJ6UFo0c/MwUceCi165JHgOjQSozCsJnbEY1RpBo7DRN8J9P9aAsZw
Mxno560ekNF9dP3QO5mGEuCMFIoQgDqpthQfw6RH6XaEKyAAdMxjs42+p3ijr7fU
0gxSHewG8sqz0CoXajf7QF7eloZ/EjMoTPwd09cQ8Bxq/qldo9OcbC+83yoW9smH
yZ30BP7hieg1JL7JDgnMuSqFnp3sKNFRdIhICjy3f1AjcRLgb+PyIkQJm1/wDheP
zhdiZqs4wi5FmG3SZNRejDsFwAHQYsiuNBLboA0tfkCijlfpCVYYJ/TgdPrLsdvr
VFqc9Lvn+QRj3EFU6JSRP0twCp4tVETgLfaMUJSbGSWJfyYDy2d2iYXN1jILGWmA
GHqVGaRR/sXEr4vWZrczTR2Iqh50DmZwtA0BzQ9AQEb7uKk+rsgFB4N031VEh0AH
yG0cHepmMyT6MfwiaUfdqEEXjcyyR9rwbawwSN35HuF/TByr/B/4soC5Q+UT1/YJ
y2Vre/AvJJRx/x+GNbwZ8VjaXzNsqdbbx3ZbRX9nFKd37OUsI2zXANPMM9NXxpQS
u4Lf1FROqIWnDNf00g68girMo9JxFgsOGVNs/3MXZbeSwXScovKTh3s8UznWtiJH
kcX38C/KG23HukQ0eWZht85eNFUiyeXetqG1sL2wU+A6cufaR5bWYXBbJd4tkusx
PU3Uyfpu147Mw3U7i+qKO77qGjrzARzXOWfTZjEb81VJuGnz4nhcuJG3EhvAWrih
W+fn0Dbu7Qa186T8PYnbJT266CaMbLH+kmdGhCv8fg4ufBBgu5trJq8LBELglr7D
giYvlozt9yUc10txacADvF++1ut1rDqILONQsLH8JCpI8AAPOCvq45dGf2Oz2e1N
M7TSgRx7GVwjFBEieSuBfRYgCxwkpHTtkgCNc7abJ2+SeBf9wYmVEWLklq7s0xZx
h0GsGPwtBmMjvDEAZFHvqrpcPmWY565T04nVbfxnIISjSxBSNCLm3ik4JRRfpnRX
EjJhoYvzqgvpc5EP8cXAdHEFjhDA98bv2Mvkqfvls9PvCE2WHeGzhvPoqEXSEq+T
15/eqZchAXCTqGRmmQL/8L/CtbgrlRSDfXm0P4OxPpxo1j3XuykrL9vox9DAw/kH
6U+quxbgCbPpPDZjGTWJ11n1plKKZfIpy1LAxttUur1FS03VXxPEsLa+PdRdUCLC
73xStsZrV4Dh84R2Z6x8+excqKA7UN6lNoMh5m7Mk2raWpbLv9coV9cWqDX2c9Kj
QJlKjwTs7NiGW6FsD6E4QzzUa0bge3eOPK1d8veUxkkBuAFKNhKTi82p694AvGMC
7ECGVnD0L6uWn4vjNekA9Cc6a7WCru0i+ceHcWxQxu6il5IZ3qtHTcd8RgCq8QtR
rAxvjKJYyQcafMiIG+oPu4Eh+4mX4e3QPWUoKkSTMElnrqk1jnmH6Wq83/oGbvB+
aWd0z6ey4xjhbitseaum1odW8Ctn+PDc1ITi85C5RCwSF6D7QhUxD298jO4voCCb
0/KRZ+tyNipy/mFb3yiguZRPxrwAvZv05CwHpJD3BgOjFXMfI0fSnRTDyEs0AnV3
WZaxQ8GUS2tC69y3KDrWMMpqLxMSS9JcDkbv3cppPnD4C6w1Q7T9IovZyvMRAQys
mXnA0pDTN6aEIAgX1EvytRbwV4tuumzAGPZuZ6iabJRPk43IxRDvyxhc1X/m/6l0
H+VURCg2NoKl9S/MGGakSmdz9CX5kIuGctXbffmOxh7vSdPuHK5UGN/RkD3kMYMy
rIe8rauzZB/gSVb4xRRbkpESgTnMQUqT8x6njbYHcL1lWVd0QTn5g1YJUQJnkRbv
ZdcJvE5w+NhUeVqs4xe6ZpCadoWG0nFegSMRNjsn7TL/A5wtvwb0tEGkaELlO1Jb
GFzmYazcS9VM4UbMKGBSqIXtIFc2+PTxDk/bZYmlHsMinj4M00faH9ZkyspLCqFK
W+yEEFxmw5pOUnOIOJ8RBtdQDUY+HsJTBRnQPmQp8pHvYc5jnO/rdRsZDsrGDYRm
PXs/XiLf4L3ogGvSsRFOb4tcNPnwbrWNcYBoTCaUDciRCndW19I9Ws4WvoWXfyhz
D3wCa8rA0RLxEZ5+6hx9uIHDoG5qwO5BioXlm05G/iNzpGPRUtVQW+kq4urkVxLC
eE4UV0QttlHovh+InLMUykHj9ZW0r2OIlfabrWSW9Cyoo3CAcWb9TJXeY/3DAQ66
enuvPhBv9OQTPLDKgztKtx1cWSg+rfKFxttj5+FNGJ+IqspjrHJ/I7W0ULRjxepI
KpDBi7gensuKcOQRPj9sBqsljGvotA9j1Lgb4o21BCuCxPPpzxYGPh5ntlrXUWyD
2RkoSfJrrQvKpT5xbwGcCnYKwbmsBGFyP+JeEibUdMPMSibyUvXF6A0V6cBOeOr7
x28xBExJKsg1+5jjCllm3/y85oZpAgI+QwpUeUvp5SiyA1zS7s3UjAjsjeV6L7t+
QHVcdBR/fd2bZim/91GWozqluowuTIIQ4woxO61vWTfMQAZ+8q0nU0TAS6zp2xOu
9f4HbXPli6wPxd2CXfH/8l74Z3vq3JKILAw7KVFcbpOVecyVQXRgz7o80TVKHvux
1flUyPKDwezRBerNYPFYn+9Med8DErBE0ftHOZQOGJvFC8m5UuEzucYqLzxy/FmP
azpgvOjVZDsTdEKtlkQh/pDRyiKzjZgTPspvjoYMgO96Otdpvsrv/nbaVWAuCHF9
3ZMacsVHgHphEDPl5fNg0h+vf6z2MWrSjvvztngs9Wg9gXBj6eq70FCPyC+AqVIG
Rg6FL5rJCshHmxOu3z+TkHM/GVKuLJBsyx/JAz7iOH4D81totygUUEwOjC4Kv1sZ
xAyuMXfQeOi42VGlmIDIUAj0lVfILZlcjO5TlbRoiQ7riV9gdM+Up7WQh3Os5VJu
uJZO1DZex94L70yQRplEoGFKI0zGFvt565ZaiA8Y8Ckb3qBNFBeYB/HM0pVTvLPz
hmIKoF/zQW5OOhRfWE6vYR2+Ltuv1II6dkqwGjzFn4SZjMf1zqTrQJM5/CrdC8Wb
l/yAYZ2rV9DNgm/tPQFHUorYUAveLmrRQd1iRVIw+FUBU2dPWIZRQnp6OfA1f0PT
BZJPL8JSS0nVfwM0s/YSCAko9o++xB9IT6DXk5tOP1SOEfEf8OFuSZOSdXOOucJd
lK7Jt98N1yh1UiZkDFnnAA/KuyrFyazQqU9u1WHvFD+Jyz7/6oeWJzPdaUpgmg0e
76ez6jetTg2hDp4kwCH0LO7tSVegGBC5kIcdLQRp9KunQ010RTFOb/PPduo+UCgB
vyJtcDRqbF1U/FIzmQPdeDQfhunyTl/TyVjt1dA33jYfcxmTpIWGDyEQ0glRXq9V
ovTGk/etQ1zq+gBtnmgyqRWLtnVGN9fGCz503qkeWgNTxqkU79+5SpDwHc7q6rWY
zKTX9J1z6s/8VHsrUj87bT9tg23v9KmVehJQoGe6Zx1IS7vP2/owviWw8N5/TctV
uexzzimyB8yZ6kKYC/+4S5coKW/s7EhI9M8r7zbNSauMlmlS/6nLXGW0Iic+RzSk
pX/Jsm6PKBya13u/3K1GqNDM5AnquwBwN3cWlDJW7y+6030FPZPvYjH41McMCWO9
mit5xdKatUAyfTYWfOOsIL8XYJPiTdNk773y41sMDV0/MiRauvHsYZMvXgO7otb8
PAOw9ZX5VmdKOPFHCoDNfAUrSML+Ik0gbgQsCr5DitC6DTocVOsMP58gdlwwysMt
dXMvNDotgrR4VXZW/n9+aoZGzNqiWUNYSm+IqFJ9mDpdLBW8fx1bO00n9+pKPCyr
jeAzzUaTHoigP2n0NGrQDE9JwLQjtPydYlrNoPaS3wzGxiFwmiBoNGS4uHNqsTeF
IrbBzEl7ns1TNJJPYy2HGYtZs5R0kF0o7H7bQsbzQTJRUb7eVpBRPQiJDEPcWApO
2dynANjaCCJdkdie7C4d0EsbXkX9uyR1DLNL7ZVdhD6bDWO5CzM+BmKZhnkh6Ipp
Yix5/y0t8zn1Z98iKlm1HQyt5UcH+CsicaUz0R8Pa2b2qkpDXOj0PFXsLuqtkI+k
vfcXHsrqIvgY9aZrMI4SXk2hkWmJ9k5hpzhibtli23cBXz40Ee93Ez8c3w5WrYGz
FT7sHEssjGyWUvG6rwDygqx5eyQOeuvT12WyLuWpZvWFJxa3hBJVdgl+8/0z2MV2
9uTaymWNtApHil9/UZVJr/E8MMZRpNmhZf6JFxKqFZSvIBH2Fy/STmK66FS/IdD4
f9vfyI8xH7L/umgF8EPNP2ZJRkayyQxPnB4VpeUAAcDmfLRbR/8er1QqGiOCQL5s
kvKOUcvA0YoC+ng/XpBK3jNvT5rFEkQpAI05RfTBDhS+CRn53IWBortxUZSEzOG6
jvEz8nmnF0WWjsNafe4s/1f244o5cWG8c9jL8K0oByAFhEZ68TyTnAAURGPUoWMC
Y3MepGTX3kHWNGNO48b15IKLKFqt1wS4Nio4Asj4+bYdGJDJCLwr3j72vHdR1vTu
Kk1ntkfBRMtKrI7q7634HPaxvQlKSFmOs3CnhBgrAtUEbd1IdAAjI4JoMzM6k/c/
yeQUhnwo0R2EjsGZ2xGi8D4pfO93eF53jXSs2YI+g9ll3ic8v5mSulyJoMTIHCDK
lw3r+n9Pi4kOE9XQHK+MhO0ilwxu5weyV7VSQyHEC3XTKr5AewNZUoNVQ6APhgsL
EurU1S7D/z7SFdMRRyTdS+RVomreHIIU0O0gfSkSFMtaaViEtrels8RYNB/OAhzn
5CM/PyX6eXabu8sfc5VFTh39uY+prI+A0mO5yhXWc6Ur+zc03RV4sd4ThsF0gCe4
5d7XEF7gnTxIUy5ceW8Hlf+x2p0MBIE/zImpH1/h9E6PdOZO4/4VOMBZBhMOM8ok
jVv8hDQMe+Ys2Q3cCG4bdIuGlTPQqbRSclgsEHIBWX+GLdlURa7q72+2mShXrKZ7
o/mHS7Nk0I5rzppENbMyh1uNCOcgzIkzdb1ctKzGXvT7AlCSGcXsIHYo0iUFys8h
JaqiDparg49eTjcUMM8N2yOYnCmx+IhXWB7aCOtL3To7+ZrGFbz5W1xcDqCLZwWO
FjVeOnAZgJG5B8GR9rQF8nKdUAYU0YCW6xzqBhgAaqOstMjZUrgW63tmT+UtdWyy
UBXcJFT6PNBGWj6D8mznu+mIshMVj9vjebCSoTuxe1YcW8it+zh3o1RTWJ1VyC+R
C9MvbC0UfKmJ2/yviiYJLqXKVoBZUIcWnDqZh/tye51iXAY6EsKYpIhTJ54Eeb14
dah3FNcKV+7cQNsysobWRjGGXaJgpdU0JZB/O1BY1qtXbc82fTkF//uEKXkM/hoM
Eprd0FYKGDsQk6g6NT4ZptFMMb2uhDWlHq62Jih2jFCoUjv2hbkQAWE7z3/DF8zc
TaflqeHsFJf/3lxLgBam+susgnpe7h5A/dPNTf8tj84HxLUfE7tPQolIz9/TdUGg
7AYxgOpDrGRklSCcl5fexXcH7G+HXat34U4WV2QWq2NY0z2yQydUVR6teqRJeqrT
DbhhPVvw7veYeCn8W245B3AfiMwtuTu2Go7J3ViTBDCBvl+7uLnixGTi+hGzlcn3
rV3nKtD8/tRAwOvqqe0jEUr9/Nl0ignlnXpsUBuSFsfU9P/Svjbsw1El6avYLkGc
nrcIfHJHaaJU64BDFLJYKtHb/M4rNsoiSaXjypMN2X2mOl0lmFNEAvvDInvH3VEi
Cmecu4UzICXex09xfs5WtnKbrMsqiZMSaLUsB4FI2DgjyrjUAUpnZm5ifgzTz0MT
JaQ27PscqpTjvFZ5k1lMEvRKE0YMgxpEHIrO5DJTkjXCGt9eI+xlhOLtBLx2tYp3
KlW7x6bVAtSMhlwxNGcv5CIzP1jo66PAGujfz9rLIdBzllUQBk+iZt/fZquzb5qn
qbipHPc96fTNXhrUGCkaUBC+l6NehKsc7hJ6pI9cDySD3nTG71C3v6l7hZgJdVUB
bAP0pkFwWXtgMKAw1z0QvKFzwpCdtXShhFPbt8nwZNHvjCokfXz5pDspnpbdehtf
1QOR3R4N1ahkYZagrWok4fRspYMJKix8heCCF6vvmxBUcvTovN6M7YsN4of85lbi
VLw2K2S6Ae59D2/DUGU6Y+rqczSdCoCZGim0Vc9OQLQ/HwTwJXGaVvqVFpqcNGqO
9lC1cjX9zWkcYx882PCI+0RzPCHpy9HYLexMhDz8gpL/XhqP1zDka9W0Ac/6/ReA
xGNs3hrqo9l1LKgecWk1BFxtYggGpvo9Y8pOaO8hg1AVfY1lrEcrDebas2EVCsTY
PUB+8dC+SdjSS84SM17a2OQCQVlkFMvD2NraHU3rLXJOF04Sel+/8gGhpZzheGRi
K95V8Vlz+mJ18a4ZcxzqWoKhRFyw3lssFnLmAVIYImX/lKYC5MJQ5/Or0WKu3J/H
1RFmKeiyPduiFENCeVhNY57R2Z26DwEWSIDlgmwo4cUytHRpQ/cke7PxVlkAUDx/
DRVpih/RtQLX1tFxFN3L8Kl08AQZQeG//mrC3pSXmxse6U1kBxDa2+fOFz443nXF
WxPhbI+Qmf2PyRyOCT0GhWJpAm9Jn8yUFY6lXQQ197nsHbopySiDqxJpE+zFY5ef
NZIS+dWzzOuqKKgOlYPULsAxCHOLSSpi/7zFfRj2hs2OBF82m6QJtKh7p/N9QpML
EjCASMb55RctgK7RRjQ7yVGcJmIeyHhiJrPmorKa18lIq7b4QbZ5CAtk3xGalZkn
xnMSAAxylJTvDY40cSLCSWZrs7Bu1k8z2QFFy3qg/WA1fX7aUQGBmiiTZl3KVj9C
LtN8JLiqLSm03SU/C6E7R0Bal+dmVt5jRHvOJcHKCNqlZvTWO6g+W3NQzD5PE/4T
DoyAke5jrXimYJ7br7FMVhmpFNTSu8BWNx3CQsPzC2VExQqetKOJQ5xS+8sehZi+
fIyoZQhcGrN+7TwFPMKSTlAhWe+Ku9t+tjlFUI4o2QBi4ZYtbAy2tzAPa/VKSaru
Dn/9ErzbGiFxDpJQVQHtMuTGooaxzsoTIz/mv2RE6EFEASuFlMhV0MqvI/3GhQyM
i9aXOkbS1m9GkITLv1ygsnaLqj0eCfyhyZZ61VKP7kXMKkpTUZ0qNTN9tIzI2qUt
0J6viWFgaQ6grWJbrdyfkt+Yau+q4txQGpsW+ktotFWPPvfaBshzxUTrtWYc2hbN
ZFR5BuMhAFw3Hr1JlMFBq06vFpPEC8rEXw+jVf7ojaUyAzvSO+avFQF4gKPC7HX/
SamHCM9/JqstPruiUxhqjm39uQGLtS7/et+SVsUZ0t2/1cEm21sef39XnQF4ruKm
3FDSZEUsr0x1pv5s2GV1j5/U7RhNeKXvFbO+gUlgTDuJ+ZI3fjtq5AJ5Ehx+S/Uh
ZGojiWT1vdtPQ2lAhh6wFb700t+FXvHTWo0dF/1ZyQt38FHBi3ai45Llgkk5h1Fd
8m1E1JOOmBws+CQDKDO3AjUHl39mkcntRo7gSkR1xrlvMDJP0gfMlviDXGgLnhIO
4MdctNADRUoLP/038CWdejE5bI9JYiYkNT0vK4Ku3GSu3ZTFMImcPQfE1EsdpOSz
nHPUAftP9c1dkcADiDatTBCwaq/BBtqucxEpSHQa4PshKnaOgCfXWxpxhBh2ReEI
N0UP+Wc6oEzuBYYyVM9H5sgQqGMf0wnKKy7suZDN0XaklxMGE3zePbEqsUOupYNI
rIKcraAKFdto5n0DhCPLLPnB33Qlygt/PrsWqhm40zY5SUieM6yq5afo0nhOvLrE
6KggA5lAoXofGwtxu3tBf4pDAeyQ6gUfSMakHBs/4zvLAK4ZpxG7JEf3zMJWY9YP
q8fXUNkzFmbxz5wLdou/QKyoP7WIzTrTpOWpKuk72D6HbnP7quiK7dg0JFNrPBnF
N4ECzzfdU5PeScto5719+e6AVeexRRevJTNedM28jgUuhes5zCUUhi/QNwcMbTz3
w5ZNWRvM2TojJlcczmhWRf6tD/NzqN5xCh90bYxufnZe+EQZZVkyA6ceF/dKxL4f
OkEFLyY5y92mbqmzQ3uNzD059re+OzaFcSp5r+7AaT6nNswCOURmfwDIlPwl7Pgz
3PvttKBBbugMjCXs0EKXuwirrCX+1+SEGKBSqNKTKtyqOMFDK47yuIISlyRc5ZNt
hKk3mQIDIYPLFpI+ZohSKLCDTOVD8MJda0jzgaJUsWjICPrak9UU7MV6j2Wm5TEp
I7k4t8dYnwqJFNh4OAMLcFvrL8ce+DKe3G1G/9qUZffPC13HeRd4uOoY8BL6CRAq
W+9hVVwVNSwii4zigS0PSH+CkIriXw2BG9fD/qRCzDgVVVHJKdvOFiy2BYjgWJK1
AdKZMuywoCI8tNLroIXVSjwVl4R1M0gbgETe9+IkVK6Nnid4vT/wuHH3n25k3H+v
WcQekDEBKmQ04qt3M/QhMwazynQtr7BFO52F+NxQj8KpqhQyf6GAZePBq1B30dRc
i9hyJR7WSEJ5J3hYDHMmrYTt9UowvQc7ukS/cIpl4I70yetg1AISSm/5mRc1kOMH
TAZsdd7zW8wAXUwAU5qBpNcUmuTTg7xafLmPWFfNQpTbmK/Nm7sGa4x+RqdB0h7H
9OGVLZKr5thYR/GlBLuQHf815RracAl/0F0bekQL8VfpLWX20SWvnmAi7aAEcDyQ
HnLLh9h3MQEfnXtA/G524fsBo34OVRV2MLo5JGnFm0FzCIkoujILSlTN+GPz8/Nj
H7TTAco244NpSGQepJifvGJqSQn7P1A1Rx1EwDEmJjAKzyV1pb9Q4FSFJcdr6cqZ
x8rMe+bXUOs3JkB4DKf+pjiIdIPAhjeXlAOOcyD+W5/Sm7n7wNpmtOHCWzVrZMBC
cu8GZL4dYc0Uz8dstQ28Xl3DNN3n1m5RnE6avQM+kFxKJD81SbASkid2AIWSQbP5
UtH2oW3b+wFnqm1RyXym/BHq0pmXHx7KbTBcLI4XVFkWkPUdjMQ6ry3dRa2LmmY7
Mv3QUITHozXr2rKWPQ9cUJpGt9xZMrunOOvZ3AuAtxYN6vmxPKpSdiqlmGYwHCgP
M+M9qLKPc+sxpejD+1boP4z0EhTDHxWOVaptctFkghdz9Yv5CbuUMqL73GT5D5xD
vLEGLtYoV6ZW1p9RTe2tdurvMpHoYlG8/FPv8psP1/yWYQx51G1EXle+nGTfJYPQ
zEVUE9yZoiD379QuSCP/YV/sAai53HJwTGXYO7KD45RZiuFdWzGkAis1JEqEqKM7
x3aA3puDEdq9/GcAgS5/qR4WehbkjnKGiktaZk4xwkgwhFzexGeRsZgDw2hJa9zC
Zykpe6sHTs+x5R6OSDF2XlEUWW7JfPQbS2ypLwR0dGSIJkX8X3I6twWx1WOgonFn
9cNrhnGAP7w3jQeQZU6jT2Dvjj/yCHpvZB6zMrcOXMQsQfnjFz2iKx+pj4Arh5MP
QGDSB2iMeBEXFlF47QBchhsqk54cT5eAcfrf7Asn6yu1zFujlufDLkXZ9VMV97Sz
IIqvhsMkgsH62F2cWIirvk3dr3+ZM2PlvK0XO+/fcDVsN79964D5CYpD4ib14LUT
MRnlqljXj2KlZF0axlD/VLuASKESLloTcn1p7CUz5Cb86OfUM0VOEd6dRQdiu/cZ
OhgYu77s2Iv50TjszvlTKqSVlxngp3bB503D/dyhJqU3MYyM/3ftqGlaW9L29Y6z
vDN21FRJEgbf2YKOrvS5VWRJCGgqDRmgEwC4/9w1uxgPvLxBuMI1dlT9KNs3ZY4e
vwxZr16vdN3uZ8C4tu+KiPRYvojR8SjKrS0+3PF8Sh+IhYby4nowR0qJSUdV063O
mLUB/pKwtV0lMdJEwoKrsg6LFheB6snWoQe726sExAjjSAJ6BcllXwikden85ut5
Wmi3fl0b5+NKaYJApvVV8CSDbtL6mgnpV/zBISBrUKAVBIwmYXjn1kDDppTe7Fp5
3E4uDixTiCDMyM6U8VkrVurpoSqiVgA1tpLImO1uEwb8pMZSXw5HvaiHKgW7e5eh
emDyiObWVjAtMkYllAPioS2xmr+Q0kdcUlm/oPUEMaHd4Oxn4NzMNlfG1tH+t7Ym
t3TU8+BpRUvFeZTJ4tDqoKpYlzxwv6JrfLvKrRAADjE3zI2zVvFD53cvGGdyH45p
+wutgVoBOKULm81dg1BGro/TrbPo1z0I7scexrBbSTqiAjldK3GGl7l1OdHyEodI
H3gHkCqfL5hujkwzwJDYIRYEr1mJcF8wCzUdssQ9NSRR8JYoMdqc0Dktf4WVwqNW
eFrYSkGVycuEpB8ZAzFmQvi78U5mEeWuHCO8fvcg4KFxfaO11X1hGDaFMuhzKkCd
Y4epJcBGrI5xR5f8owI/3JZKZSCSc95j25OrJd+v+zGihtxv2m/pYHYw0FdMHZkC
F/QN8+u7orkVWjkTtxUQw5EIbaG1W9DynAx6KH77CawvHVSAYVuv1KrwqPF/vlJ5
R+UQVSbY6e8jx1+0OXUcZgWNCuL3CZAYyV61aqKoLyPtBHXR6+2ESYN5SXEQomG4
kftoOPbyh+EX90JH5anzSowIZw7JB+JzdQaSK8DU1PIYJihhARnAKpVL2/uSCbgd
6fWyUkXRVw8wY5PsFW23R0L1+nZhTlYsvddLwx5t7uISqBd03y7W1KMYihJ1p/sz
YBvhsmN6krQwbTPSLs2O2K7c79aR+PRCygKh8rH90iZCUkav450nyBJqXMH8veVA
UaxeFIV6oDY9gnaVYCfplMmkHJpxta6rsixSIc8S9ASDmE1fNtcpe4zISMG4WBpz
yol+7p52ZXvlOOJTYkyZbHxMbIIQVqGIPHPTNoQHlu1T0sQa5QOqzJphk3eg9wZD
Ym9o9MFT/b8FNMsIpR8Hv7A9xBw9qGbfy/BZG88TiwoDu8i2DrlAY5qh5YZjilsU
Q/kzh1gcAWB9783rcWpkiI/Zdxz0fbMdX0RyPKhKUGiNGwb2X2d/fK10drSbhnwz
sM887KgGl/ECmnZSmyI2p9BQpp1+94TuMOF77Y0dHiqKFNuwkpnMX6O2ePIYSjiJ
dvkDLdvsG6vDzHzn+l6EQ9Z4I1IRmJsuWHqTARmPHv3ycztJN7Rrbaqz7k9j9EcQ
L2PVx3jhIV0P1omYXIe2eDLoJuvFR31vD/C1tsD3WP8fg07aaNwaf/vLymhsKX6r
6EW5PInRBHdFAaLf6aYjUFAzDl9o1b6ubDVoj5D12yOFkFSjmgaibuAHMdZJinx7
Pj64oVHmn1aE1nGre9CsMNfI/+yh61aNklC+7/1br4TsLZlgtqY7RJG9j83pZRPu
WoteixJp/QqSrroHBYLJBlb8WnSFNk2uiVnLmSj9jAaKyMLLZHwAlKLcyTF1vy9T
OsipnFZwYSJDplS69wMNMMkVQEjbUna2o6iPYJ9Jftw/oXOLn42QB7fzQ1JwbW0Y
o7BAvAGFMgLlErV9BdqI8RRy+OvNeLMsJ/FgbpOuvxFs7gTKVeKuCs59/ZStFbED
fq/vRPVh0CEpg4GFYl++7tvngQybidb7/qIHd7mn8a4ezlICNTjsnUol5gDw4MnK
HNWmuHea8dKv7k6h5oDczQ7i0nLR+vX5BRP/selomUFOEOgAGtJVXPD/VBroOIDs
KdklJ44y0q8L/BMSEDxBdRZuug2Dz7pe8O51qUZ2b3b1Lzsspfcr96jcx2tisvfe
y9NGGduz+OVBCWXd1HE+SCXv34OKeA1z+pirnFYPKaaNHIb+ZwHrlHddAQeZ/XXG
527MExPlCcMnhe6G5kb51rBRKviN6YTykSuZbX55FbOvmHEsUskpOR5QU7b73LYs
todWItsp9FLMkRcgF44NOFIGaoHETovgjIkYFGckgUGOkQ/s7O8xlDVuUumeNC+3
oO9Z7uplD30G9ogKGzuhVbTDTDV6SS9ZfjSANowtAC6P6H3FZFZfUwGo3zgCGOpb
MZJlmlEaL8i/EAtVzwt1/kD9dxQhLd43VhP+wY5rn6B8Tp2X3xoi+cSLiLZPYwdk
v8vuIm4DT7JVHWKqHAwFVhkTtvSvjaKAWrgDx+tLPt+UGHNcc9xrpaapKcNFkbld
HpZhK8lVSbog3trsgUdI986dUQmkDA1NjdKPeiwEIhzgRuUzXBY5Bd7zk4D94n/X
mSLANCwLuBt8spsjAfMmdTqs7tZj5tOspih+VoCFe9s40SPgdHjcaYT0kVZKhnxI
ylwVcyCAuMaeA9c/fsqMD1ZYq2VB5EKrtL5dyPzod3K6trmKTslD/7tL1HfcyBoe
/eckn3TV2O7WoNxewP3uLNOhclkQtY618XeJn/KRYqo+9tngSW0k4IXE8w3osID0
S7ZWhLBrcxgiacF29NXr2Xvw95T8V9mjwRx7uaAuK+GAQXVjs5b7230XvM8EQ9oG
lw79/qFPehb+X8lVFlCPMTZOzZvQ35n/WhsgBPcfMnBMSkA6qHgFy8AUqVrbWDUx
++G4577hC9snm9CxT0JNeVnvyUO+uFISjk3CmmO6NmNml3Md6JEYv35pmTXWCGhi
O5SdMK+rP6Yf2N75sXQlgpDpYSt9mb2e1NdqCc3YKr9f3+sei50AuN8wFk+l852i
pHJi5kO8bw0v5TjgpvN02p8QXJP7007aXWmU2li2PKA5YDtniXdUSSYAxoGZ6Z/w
zd93z6yqHy46Vr6dA6aUOFd+EejNmnlLd46W9q6NYkJ5vqeZZNkhYM27RUYHimZ6
5xZ2mtu1KuiZMTtp+nbfeS8saMwND/ZS5KRfwidCY/cNTprpBQ6+qL8l1hmtIQr/
fZYeKs65lUkEouKmpcCKjdCGFUqda6QUNm3n7jbPimUERDhJB9+6lRiZEUnxvOC1
T5YGePHZC3KtAJPrcSKBponRQRdu2Sb/TJ792ul9xwlLZCeNpGI2fzHyzxAii2Ko
RAa4M3b0vZ8InXt1GLmUOmmz6DPbCZqZh7t7jU3B8arGZ5FhD1yU4BcgtkFpudN+
BRIJ6P6kn6eTNngaF+O6wrxbzhWzcBQWwFrY2vTAYFzGIRu4UneATlXJ8X/5NC7Y
vpl+Ep2kE+b1qa95wlIX1hh5Zra8043zlKWnDVl5oT4hKXUiCInkX6ATT7zm1XyP
gMtV8PYo1U/Q5G6/hFpLlqyWrgm+P6BS0x1XxzvRhUGkUtrvpvR483GG9VBkYXCp
FfHRt8z1JDp3VRH0kERnrLp7R+cY3dAm6ECAba3kGeS1UqWEUuGvStk+Nw6jspN9
nYAJLT45Eh2PXUpw/kTZMfZSC4VhyCGRPe7sVSSO2C8WyN92TgbKJzosdyDiikpO
wC3340A+PFvqD8n1m6xmc8GvyxgWEWk6d1Dx6KP2ima3hUxgHKSsFqov1Ju6fFh0
6UvoH/9ux9OZFfSwyOZYZYc0I00qlIfxzpVWQXycZZ8cKuDLFVcSarvhvxnWEMOv
AAcNwvHvqWT8klcZ6/Z8Pbe2J+ZMeyLDsvosW4Us2DLty+ftkG/1jaN+bAA7wegE
JLF2pW1UQ4O9DMWORwog4o0MGcaHKUcXqK2V0Yw9JFsVFyGlhQUI44E3Sk0iLjiH
cVjeqN/gKmCteOIvE9MEjIzBk/fnM8/AVd7EoeSd9VwRMt5X6AOV73JfFF6hxW9j
EBHjT6bZRynkZadtESW9geqJB2p/derYGAeTxzU5nKUOpkrLxvUjJCwn7dgJOCl3
BzCxYXzTYbJUccRvCXoUYo/EzlR138KC6P2xqasRDLwAASan/bf9aR/q3535VRZg
22xallTyyuInZKYKxZuYO3qGy0BCch1ffSphhRbBw9iu40ydls1gYGYP2r+fxsW3
dMkk82FgZ3N9DAmygZSXNFZZy8YfYLeig9sMu5mZA4ZNu4uXDQBaLwCz7guYX8ba
VYREwuMpK5+jQmpBdQaOQBURmEqBE9aWfqOS12/NJo+mpg2Py0pz+OHeXXKRJHo0
6sEM7t/WCV0enXlgp9HNpl5rHQGMiIaYZ5zffCi36fq5CDsGZi3nYppLflJXGYCs
pl0ct0RXJv9BM9BUzOnh1wKAXK4uVhOvos4R1h8cCEOAv58CwdfelhBF+tb3VwtM
wvTfohyWWte3Q4kD947VssTYwSmQCh06Z5p5QoSCKHCBU9+nOwlkW370kZy1ee+P
VA8dk2xNK2wTSaT8T5axQOjS4ARt3828TqbidcnxZwq+eAfRfpAyL6CJ4yInLIti
XzktL4/4qUFOFK9HrnAP7qHn+mtB7fdNoEjM5Ugm8FbuzXFl/R0UUVFv4jBPnJXd
e5Soo8wmIlM90HGEldJ0vtjGDPEuN+oD0ibd3C8wMW0RAmkENK7HvkpG9MXXHvwi
Ksm7Pk4TjIMLQE7B4AJajFCJ1Tjth7yt9IEREQtw39ZNx+FerZQzOyBRtjv8IMTH
9OpA/oc0lVu1nswwZG3izGCvWS9Ndet3IQW3YaE+DUnFll9V/UzOVS9AOgpNBC8H
NuQAzfC37cu36jI8ALejJMbqaz/09z6UkvKrlucZtjq4u6Fu++UiEb3IILJvUQEq
9eL/4LVKZ9t+MvZoloV9QkVwB/fCv/XnJzCVOJZ3qAgUZY1KlsqHBiHPRoSOvu+6
+oo0y5TYUYVEKyRHPeMrf4o+IWTNC/zLU+RDoWmOKSc+SG7/13EtR7+xH9Dvku/B
eXYv+wXK2M1dibyPkmoU3epghYe69hNzFO/HirmlcguM7KqNWXJxZ4/FLypWjLsh
E/NgMcP9P2UkoDvReYQ5hzZyX/lRfihfBnXtiv6hMS2Usqlxwf4eLP3v6UE/CmsV
BebIJprO6r4la4evbo/kWyOg2LDJ5GSDRYPjmRbjWV5pXw9dchsdg8xrGIQAjqTT
ta2b2SUJe01600jBykvLFoxj4MB9ovv1pnZ7KMql1QIh+WSHAnIdy50Qae8mKXgB
YdHShhLVYGWyK9rxI2aCRAafTHAfP4w7s8mzCwK8ieygWSyUuQKYErGc7FDnVjwW
K6Hsw9Af7eFT0D0nCVzeytabMs9TXw9l2sHvlF8ilSL4n1aCI5eFSL83uSrMuAfM
vTfBmop1TsHEQF1khn6dFL+pfyGGZ+RE+Y6xVO2LQvIn6RZnMgcP9vKz1MvELWwb
gEcCVyJUWiQZsLRhnj+AAiUshbPjPZx9onmLFmnSUNL2CpaNV893CMO86E3qtXve
6U5Rmu2QTM2g+V3mRZcI3k8HVLv7HRrC3QwMSHonGgbalOJrCa3IP+KTy2YAnSRT
hP64lVBu6SynI4CM/TU/OPFmfgXEsKjgzWZ2dM8KT1tsn4pmAyLxZaaSP1BhUk1W
/NyJdywAxpx6nmZPlE2ARRAaxQAFD0oOYVQzOcV38bF0Qe8+kw6SdSNLiwvjgdkm
woC3GmhQ/iK5Qltk/TsMZUEywexhleTwO3BlU+BcEFii5JBkicRmuCjK+3zd9wO2
fjHqKARe6xx1TO1wk8apl+ebrMPJAggKgJHErkXxQMfXksUzsqS3H3XnDj/FjgdQ
Zs89h+j3LXA8OxgY4+XQzJ41mFLAMPcQL2D0rGYmMn/ts66hE8RLDHP27f1DEBr7
4UvESIq2kyUyqGa19fJUKw4/ohzbd9ED0Vo7GyG9wVzReMkcFxPhE1iH/LtW/KsZ
WY83fX18g+GEd8yqZlCvC6tx+3/23AIkzHCX6p8jnI2HgcVORf0ql3iy0kAp0vLN
w4G6IpHDP+4GaojCu3s6E/hOsGjNd3wLWg7GYE/2i+67qlngCMfbkuiLOICrPlX7
K89FIhGA3EKe3ofqeAUD/9UIQ5C4MaS42Ms9W4lEwgPUQdiT7ks+2t2aM7nI75Nn
riTOiKFw+OfRK0CglqHIzxf11O0WdIthDH9gLwfU3TV4TIeNtgRSx6pqDOicvKmx
tJqXxv28nnfIFevW93CgZnV4bky4nrboOAesSN0xyGxepqGMkBY2Q3ILkeD2A7tx
RiKNUdzElbqNYq65mce+RQnkfcYzbDlFn183fmWmRJHocl+hlWCm/TGnqhDqyDIC
ce6FlSMCky7GThMUnnuRbd+UT76jzyTN2qA5ZIo1A2VbUBbhPwRNGJWfI53OAVOL
rqo3tcQjqp5Dyv5Prt42T7X3avtvjkAMOBH6CYOCvvhDSUmi8EaQ7CKiX7wNnoVW
2Wet+3RhI4JApBgZJZZfxJxUk9vt3hqJ7rrESUbdtnyW9s5hZgXgyChVjtFogaxo
GakIYMXo06TuEjEDUeam3xLwfThLWovsenUmmD7x82BPYQ6KQm1rhWx58vlYdLeB
c7QBM6rJ1aKTzTZb2ZAwjvtKG0F+43DIKRl2WsuGo30Xm/JpPmWzZy099XkkbYd6
3O2Fx6RBKgvgiCxsMVmU/XKk13A7VsSi9u0ml88h41Tm2qtJgdoS7wF0rk/PJwVp
CNovF+xf8X4BUEs0iSqC0qGWwBSxWLwi9275JdXOil8OCRoFTdsQt+QOcaxm2NFT
EBq4RHQGSEp00xV5LRZUxKXepJRTv5dCAVlbraEQ1VqmJV7tu/w5rCJ5R6xB6MSw
iOlfBvN2VYfPRjbbsXF+j6UbCAyy6S3BgLwBbBdLmwRr7rpSbiDLsd63c6SI4L+P
2P262Mhjf/bBf0xWaX0RJ04uy0O8oKE5lkpIlpQbmGTqsMiPZnY13a0oSjYB7ICJ
4n0ZabKmp0Tz23q3HMN3oTF3sKT9mwBntOGB/hQyn8dlpteRwa0wtkRQUYH0e0Wb
aX+C6UTViKm50FI0aQ672l0DNcYd1zcuybgtEQcgkdy5PGdqEAIoChIve6bPHzE9
sHysEG0zKi6W9HwilNAV2sniDzDGiabRZ0Wo29RboIm4Y05/ewBoJxnTGTNQo1l7
8+cylHJ8aX3NPa9/k/2l/T3IfiCPkc3mNDMLjtj9rWq0vENJO/M0pXY7wzZQfDim
Y+4K/eKxMvehbIb8K0c9or5iLagFHziXvs+IPEp69Q43VR/xLmiC1vH+j094M5AD
OPGaTNU3yfOTporz5xlNIdlOLi5SbfkiukDZRROc+2p5L/o56dwe7YTSTdiQ65u+
KF2GTo5e/qBJgRm1XyIv0+sEy20qypC4ogKgjKONHQcFDWM459AJzN612RIyB6Fx
CLbnOSCmOE2qrJOYQKV5iAc3N7cpUl/8hgXzqeze5ZCM+YA3hy4FMxGhuubIrza5
ZGI4znKAfkY3uAVZDe90L8QG0XIpxBMKHTz8yuVmmFZo7UqzJ6qbL59EKsZGnMVq
zW81kI0LH1vfgkCPbQ+Cwz7Jocb5AoIxvqP1cVqutFJTI69uY/QAqcrPsYhw75Fk
9S8rTSyPvmO6BFAnkdyvQ+EZpHfIZzEJ152HAd1u/WIoBXieQkIOo2B6IAP9MZ09
OQtYHRk3N9NfE2PQ/Y/uv844KCUBSnrh/YwdFQj29pa06CYNKeiRUEyEamrgCcLh
tdPNc6cza5cMwC8RuAdvUq72rGyso0sDPNz+tJQ43UUYS/sRxPqFqS+4WwangUmf
NxOhsw6aHDx7+g2n9aWpxWICcC2nKqeSW+VvWNvAeUVVkhPpGecqyPJq0B5YBv74
hpvkgmPGH6Kd4K6tibSmBvbvWx1mDaKSRwPzFYnS6AkQ98Jbwp57iPjwLoxZX/AS
LRqtQztTv3H2l8xuA7XJpsW3MmMqNjIRXwZsGvHlTDXAvMeA14yTd3YYM+saSzui
hLkSwi17yuaLHLzj4A7sRJgfFLq56pQPKS+648sSzQLKp1Pym9KkzCPVnlETyXPu
fN7IOYFpJHFr7pY+jH4UZ8WXTSuBjpb3C7OuX9MLcxxBZXOHIROpJaPrfWTHWS8O
anqEptxJiKRC2/cvNoXOOSKXvDxS2hhrJimp/MLpdf6cfQgyVEHn6RK5nHlUCEyl
ObwCjW1h6nxwr6XqtDKuUq+51qUuCTkEK6y1NnxCKlQGn1FC4FOLTuqlvASK2LJA
C25Kce2iD7c9CGg4ZFnX5dEyiMTJsOO9i6weG6S3h4Rif+3r2fYRtiB4TEhFT8RF
zs/bLuqXSG9DwiweTvqM0Ngn4wCUOtzfH42VXiGD+b61frZrzNElmgH3JLHW+4cu
zd8MvOrSriKEoX8OJpHF4DEMl6w8GHKn/kgNvOyvjF1Z4a3YFGitLYHUaBCF2UHp
v7d4zwGEY7gYiWzZtqEBl297rVw4g7hBWbuOoZkjlQIRezGwhnba7zjf4QMfUfmI
IxDqMZv8SwFstbKZGFz39m41KriKozuz/ZheC7E/zulM7Ggt171MHeJR6Z9R7hx/
BOCoVpKt3yna6XfhY5ESJkyOhLhNuqDkPcbRGoQrBMzQKV1Txbr6CjqFtYlFz+gE
xJmmtUvwKcUN3XXuCUU+aJb4i0tLXrRaBZmg6UHkBJZYTK9plolUAhPRs5QgB2/W
iUgyvK4UTS4bHmwLrN+2iBopV2rlekwOsEOKpkTVucSb2CbMPxO7xFmfTRZ7/+kU
dkwGl+HgBeRLhkxuyq+zDVEqc14E+EcRTORH//7CWT9ufCX4UFdijwCnD66ngljK
uOp7aDyaCqBp7VwwTpJcJP383LUVM8w0V3yO5pSPBJ/eXByl6iw6TR3mqEIEhcE1
KQIyARn/jiMUGwWwuvz14Fwl4nLv/q4rkhuX8J+C8/dExtFlBLkKQM2DTzPzUjrA
8WdRevYL/oKzR+tHv+M3B4SP8kZPf6sCSyHjYPW2lYUWseqRP++67wvRSOmuNZc+
se+fJ1CXj+juBHG7dQJOtSENATkkWnD3NuqjMLk+/U32HiM/w6X8kG0tFF/MEC05
DoKhQvqYGMIxZ82eEO1Fje7uR7hjPlxHZ0RY/yv+EUcXwDBfTrENMrZgJHrlqeAE
n6l+X7Lh3hgvRgY4U6AfuE+vo2+cq1uxqiZuIf+iKYjnxF8itOS9YcAT//ZH56Db
pOmdVN5NJQnfvaE0rXH3aiOt+NoCd8ZfBWTh+xbFgX/AKUbOrxvj5oBovfZU6EHg
xhqtvn7vDFbUsXmOpYMCVhbvIS5/hxkwY2s42jVvl4RcFnN/CEfHf1H8C5pEC2Kx
aBSTRA390FOp9rkrlvIvXPaAbwX758D/BIXT3Heqv5iTeCL5Ixn3Wbbo6+TDkSdE
XpWrjLTJJUSfuciZ6C1cPdx9wa8Mzbvh1BeLNlo2rmG4qhKpXvN2m9JF9HzAYWWc
Df5pRmJ6TpFpN1jHoayjbHXwrddU2dDkzj7NdXBKHyPeR73U0lb9+csqgCV7UKJ2
GIJlJf2LpljHa9/yyo2lmMUUqQUlTeXzRu4RGe9pPamnfKEq1Wu6GEOVVAJRdza2
S8avI1honwtJxTFTwOn7QPxeeD3n9dqjwWw/wwk+zQrpC6oiBo6dEOlhRSQVhD0I
cGg1icnoDn/YCusMLS0LsTqncHJ2bE6sVOHVQWpevBek94QGxlyz5AVwS80aWcEK
UypvyVuvXrvP7ILdHrnwGG6rUsDma5JSLWBSJR7ZxZ/NGDwQB5N2K8S8Jwdqrhni
gxFeDyHNyypfpfMRSYvDe2yljevp8gskyywK9GeD3Km8dm6PuTElNjEvxGsv3SNW
EphKUzK0QcqvU1miT9aLZ9+446jlW7GYt43LUhrhYk6h0Isr5yDKOinEYu8bDX1O
YtKoGfWwfI7jTNksi57ijiAaH7zwMKOlqnsRFUZ0fW2ulRDHwc8mW+E90xL/wEjG
w5jAdizIoMz4fEdIHFyRP5HEUiaR3Vn/PWEN8J8yjMYBy9DCoDCP6arplcgLUxcN
pJCbJkhmAWy3FCUIGxSYvs2qpMKLHKEoHhuu28DBrJ/dRtIpnMpz0fBdFesU2+2T
ThAZE8VkBLdSLjVctC+X9INr5GDUpBTvn3i6yDZH/8ZleaEUthGZPENv05Hhk/Yg
Gg+LSohgDQfrwT6cJzdpbZs6saJ1cpWI07bA6tNir1u2eq40h+xOehJfS2bUkuXd
qEkBDvcayu98B2tRvszMJPRrtFFsuRnGTr9OAowYLZ+VOYuAzKZCajmIQAwklklP
/Mbu4zptWhF2Nc++YhfFXaQUzHtg6SMnDUFmLsnaQQNOJwq/P2zCIytrSe7DyBwM
Grw94K6aKYEwBZNX74t1it+eaDIbg4yq5OyC8Wn8Sn9HpqDFWwQiJSWT5YGACrWd
p9EaQQBR0DpFQH49XkgOftVRaC3FI+yMdMA40NTpOZys9KwRDk0ANJfrnBh5K5Kn
bMJGgShZw/cw5e8DxDN84g6VCd2bmK175BsUSN4ioVbnHF7M1vZQ0Xpq3vvSCRbT
dRaGInP9k4lfJ8r5jn3DmMLNfiiLIQ6TArNfIvgSyYWICNjoehOneGhdReXqOqr+
laRrURHd2TMvXuDcX8WzpInJTJhuFMTvRrjN7a5eDj0Pwj/DXwHB9dt4j/x83z1V
fZZrHTGvGuGoYX1x7rUvdQkSTYSiKYhBzKMa3f8hWxG2Inw4TALU5Z41YN9nQD7x
upItAJ3uQNKoJiGcJPtDFi8PHjB5tjMUfffnF/JTe9DYfOx50hU6hrKXvMBM+1lW
vn7AJzISeQnnQ3kJDCE/6r3FXXCeRrAfR1DO3xRryUvRk8F6f4VV1p5hbqfYy8pS
agIKnRBHQUKg4FkXmURGvQXUU5ATpH5QihyJz5QU3VdsE8PgY2LDsr6XLahjTCaO
LRe0YBDlUw1tG0pID3HWYTQOuXUsby/Yi/CM+YnQ4bkxMaSmfgrmCMt95nYOiLwU
xgRReRpzvmfUe9ktK6t66Co+FxOD+yO2xmtDqqJ1IsD8FM63DBbzXBA15bupHhpf
BmLj70cH57c1N9i2duYZvU2R+zIg/dbAuex26fzi+XAD6uRR4Xaz2uZdH1d2wNom
IpBSqXlF+at3REIe1NNfvpFcFR6VfiXKATCHRQc3wKMcrJ/RdJMLnYGCX3u9kAv7
cA/jmFvgOeD8Tos4HTL6L34D3QdZ5VyWkn13qrgXPtFcEQ+13rgqX/W1Jw1zQqj4
BpcC7Rf5yAmnrfvUP85gS4MfBETTxnv3x3TwZKijuH9XJMxgPNA4J1Rh1j416n6D
486KSvrTiSNwJlWpc7TN3olT3h5VhLBPuQJAQcaWhiFzUOGk3BGG9X3YOHvt/bfD
Y2io7Id4ngbq9O5oPms97uszvq06mmKq3Xsd2WYnNU+dbyF5P2Tce7v/4mzg9Met
60YHGNpDwYtLKdvo/oe23Z5lmXbs1byGBO82QYS0ViNo5uQeah8FFSaJRNTmnzcb
gvko+T/KhfwVBFxsi6zTysxJ7TZAFHUG3xhLTG6K9Fb6anU6mn7gPdf7fCW8EvmL
pLU9XTMLILfDXCVvBPkdWLe3Hd/3ad0n/d5urilb+KT8K6Pk5aM+8xastAwcFK6V
8gVKlFtzk4vkgriOOW4QsxHBj1zoisB3FBOYu0O5/BQ4XDDAgk1puav7GvMk5l8F
hXSN58oNNF6r3yaBlFpLhCYzJFG8hmR4bWWbDpZsI6UMR8Ma1buX0vI9zGZ6u4GE
zUnv7dmPZK6sjwXBC6L5Qkc6IBxb/nlr107kAapqnt1N9NgPUTY1q6H5I0CRQsG5
KyQrXC/YhK3yVMbFq3czyFF81aHtsBxB8LH1Midlg07LfV/K2i6PupzwV1XEp9uX
xGrHvcD3mDb6ebyu23H/qpYsUatOQ8hS5Z9gTzbf4zavgfmwTbHvbmqSsRQB6nuY
X3akkiu51s8RxpNmGotBr16tWo9PfgyWi9HC+fskOoge1LxC6K6n5sV7PO84RqE+
GN40yFSMEj/sdhxzkXFUQkvQjmdGZtIOMLAvPhime01QjXHAgmQ4q+iErJ7tnFiE
pr6JMMYUoDHosWf122Zby/UDHzHpYrdGyajrRwPNAERXvQTzxQkPtzjK3J+MWus5
zebTtJB8e0x2DIkv3754tJyXC/zkJamrZimY8vRzWEQCz6fqjo9ywqaOwvfr5EDU
GVyOk3wWDx9kQ7Vvx2PCs1imj29VACdydAxiAwklCq5RM38kgbkH//FQn4gyCBQp
eib24K4h/ZbMhVDuD/9qta0zxddLoK7wCfZQeclXn8WUhXGPkimdwcf8YvOR1HJC
zfeOLa1t+qnKzvMqdKIGrp3h5VroNi4ojNJRFW7S/ZMuR+SQ8G8TWkzTikH4/v6+
W7ppvzOSC0+gmpBQUefrLBqIczxTFQTFH8cu3J/DDXbsYmaIaNk5nbpEoZrg7D/D
qdBCNNvKLRDvg3Hc7FjbPi3dlEUAnx7rtOj4FIzrZ07QQ9okEmATG23mdIRJvCEk
1nGknrTBFKaph8Riis7N/1LudOAMeiWE8lzAfveWNgqgg2IrBqxXJgcYmzeZhAZJ
18kEx4vD6Q4wxhhKUge3Fp9sN/0gjt6ODgYPSBwi5ai9rlv0wvnYcAmEgNeVOAe2
xzclE2wr9j8f2bHJ8Id0KBoxsZ0QxWtzSjASkeS/NhoIeLreiZOqEOpe4qxTMYVb
TKlnpC2RDeeZoHL+bmX14Ps/doCLJVjoyWAxa22zU4QjXq+k5L941rIj2deWRkip
Xqoa5/CJEcl9q4WjS/4tmHUhHF7Y7MvYQ1VQN6QqvEGFy/QBzh8hWW9KQ3/hS13J
O42CaHKeyOG2ylz1astJ/t7dXnMKtUxBK2hHaGs9YoJHHRHcmHsP7SZ3yB3MDxH5
ILWdOM30qVSXlxFCO/a1WM5Svo3trPQn57nCt2cPcNAN27iIt+mOqX8h1e0modzl
i0WRLwxCfP4seyQUbH4Lb1F672Wd5yKn2GFJBT0/hBu5tVgLlfpuNm6ZNdnWwm96
ncALmQTo9ZrjDFqDhgNwcBxFpLmp1pJEjp5Esjwl61SiJOoPQ3VfNsnEkaQaESl2
5v5Y8YMUS/Dqanqx5um1qJzQYeNNwNJd92X1SK6khWQCazo4XKtozMmgiiLCVI8x
yRXIJD/SIII427FawIhkWtCjmC3OHu5MmpC3e21o+AQdriVrzpLb+OT+iW1CMQza
3LOaRZKvS4Mi08KcQSe8iynH4SrrI0MI8Pnj+eNHv5BVy2lXN7YHF0fPYZHtc5Su
nfm8AyGud9KP/Ca3Vw6m6/woV6jlMIJBZxaMmUqC79MBCVdcnogH7nl7Sy4Os3/7
TbLibHWUF1ffcTvPddWW7Df7LbeOHSOH2ZNvwsBOuc3tLJUiB0FRKXYUET8tSr7p
6pVuUIpJjcnAY0NtighJ6HdY2Jvlevdq3E7MNgI3BxYbMnrKgCTkUY/304awmrXF
RSIoMpRH5Rrjnps3fsrSPEcccgJjT74zrWgbGs5hgr4CCA/btzOI8jECH8J9L+Ig
1MoVDBi1NfTBhssDt+p9w+SJ4y+qTt2p2jg17wNG4vJ7mro8haRn4myEqPC/B+eK
ZoSvyB0UCGm9iW5COXX5fdCuRBTlVYwzvbOpWfjz822SJobC4MFTEHYdgBjq5YHN
c4oBuiWpI3eidYN/9X0ssmP//Q6nH4BNjKT37dygX4J/U2TcVMj/ZBuYPQqcxbhS
HrVBfIUnoDoKFw3oU1gcughiC+3M6JEWmNDRpa9HWck7uF+MyeBd+JkwxB/lEiq4
djYv+n+vpvagpt2StEGWhvExpTOG/f9T+XJ1eXsw6m2yeUEixaxGOokxA5xk727d
32lqA+yHU9pDqCA4NXzWWjiaOoR5iszspwEO2WLhzfujtfv/35gFM62Zzb8jWcJd
kyoxOJ3goqDIRDCQGMeC0nDV2NwVD2AOz1z9ZrcR/7vg+anWCFBCjtdqcb9O5NRH
I1Py8AkxTKLXYzInCtvIu0AgJggf3cO0yyJ3j9CtOy8HGHEe5vvEZGpyFCE7kBDq
MD7WTN/1tgtIXf9GI64ONmYIOGjjgtMu5t2QDP2B3jyXXCeBMZFlbm+hEfJ/Lase
RArFbcGmoe/XWi7aNK9WliNqYJVxRILWRzwoSGQfsOf3FHwz6Ys4QpsBUmuJ6o86
dip8sabfsXwnhwPAdRYEpu5BBrt0h1xovo+uw1h9CDgFjGgW7CjLJhzAvSYNXxoR
8BV8sghwt8AQgv7LsaPi1rqvIL5zxxk5jzNy/Vk+mPUJSB0agXs4zb9Oe8TVoqOw
LgeNiHZeXpW8J7L9WXrA8Sd7h2W6S7unNPLP/ZfESf4VMhAjWlOZNC7mLohggqFF
Ff5sn4ClJ9J25uytS06aspqbn8hWDEXvELtAm7eNmFHq2IAI+jx719Qlua2RvyIJ
jZJMIHg4MRSKN1GTJi9PnjXsSmd365PptBuqFBYU0lpewM39scnh5JrdWMUx8aOG
/J7F5Oi0hXw5pU+wqroWFC96g9igWO/fgJdS6RNQC/BBVV45l66AdIcd0EJuQ1p/
nLjWo2hP2PnUusivk9Tw7bXf3QYHA3ufiTh/nzKFnUcJs23MsaJ4WAfD6Oupzqxu
+nlGewi5jawKz8RKRtqROn9MYuM5NmvGDNhekPCAmj/8/rGOVUNeonu1Mi7j5GMw
rYEcZOcReOO8c5N/r4086zKlQmWIRd2mY/5pkACui5DlshjN3sJdVuIgM8psYYYl
PnnpVzwZYLGSWztTG+GMy24bSYQ368U8MajoWS3KKK2wX7wA90GLH7p2ANY5kCmw
ZQj6hi5QPpp1yE3EQdg2TU0UypNsO8Id6hyuK+a1W/XjsRofElfRVLWd+CIF0EQ3
JcYvoirjOJOuSf2TFlguj9qhl6MHLUjZXDIwaLJhj03gUn/heRtEiRQDATT9XJqM
J2b+J0YrrQZutH3IDnOP1ftee+uHnyX1dSZWffOU2T39f4Xp6vjM3CGiiLvA9YYX
bfoIjhvdEOZP7W0Ft/8stR6/eZpO8sQuGmuf6wOAKcdp5Q9cu6mTBAsvijZkXrIy
7+0qZAa5FJVwY+cfYN0XeuyBUDwc+sOuw4AYJS4f//PJUSTjYfkL+r2+5Suf3rBo
iJqw66EpXXMi8Svt/LdA2uyoZCZ1wABb66wR3y765jLl0Mu+jzuGXUDTcw1p+TKt
DM51BBPLUYvDHdajvWuuZAM8eBoJbbpGOAANnYZ4M7/mYlHeWs+kkMSKE0wQ2dcX
Qu+aVUlXsucb5PlvO7NMW+nlY0j6EkHTnaJtOwdOUTMk1kKf8CBXTbqi7V8JQ9UU
ssGLekw0r+QpLeVymaLW7PAFNH7nVMmQ9HlbDgTUqtQXDBmwiebkLxivfDlyYpej
JSFDl5huMIMiUkPSrHeeBJRJhG5xx4I7W+tVP3NYZ53PmMivwDsImB3oKQ2sbA7M
HTG+pFodt6OI89NennQ9VX+goQUJQD+mWCd3v28hQ/7jF7Xq3M72JcW99yyDyxrP
t8v3V8uhcu6Rh5UcMdhNA/9QVeDxe34Hka5NIWD6YpCfsWQBgkCFQlYIiE3idD5p
QxLGg5e9VVXEz90t5knuYFfLGkdBGSfZjCWXep+b4qpoVTLBvk3BR77z/B1y+k7c
zpgCrrvbmiRJlptS9XPshciTUfUZBVUvHdULBtdwhr8q+YpYuRLXF0Ny56/4Wak6
4l2oJ92B9zj+emjoZJOB5vlaGu2/Iz9lkK1JAsIWPMS0KJdpdpybr8lxzUGuomIm
aootEP9K1G/VnRfyadCdbiWMdGGIjto8jQg3uBzy1IQMU8W4ggQM8BJi81Bu3WTf
wx3Ez2RreZR7Reg24tt3ftdLJfszUlzFVjZeysE/jXR89xRdjZv3rCjVmRFRx70i
dVvW4lC67ma44ZW+szYQ3OhzDdduI6+Tx8r1T/x4bhOIrYUh5o5lUgu5/KKR3ssQ
A97/f3dDgcpQGvtpLqNyzMx+9Va4FgjLX+4tudnKv9ctr4r648LslBAsJL5rHENb
W+E9xuxsPmdnlqvJXG+6vrLeHhmAEA/AgMxYRklLQnQqxI0tMm1DS4JOQFSBLbh8
F8eYML1zTVNeNnENJuKjIKMwE/+9c5L7mTzvBNSFpg1E1Q+6NRmP0LDsnYnsq6xC
tyT2qG2J0EdAitpLtE4mtmnegbxqA0EqdXHoOEdi15hko5p+ZNyPSpja3BFgBrWx
0slY3NtfFQkLmSwzlBar4huwyLaIX+JkpRhI3AoWCYALzX/Kk/DKuHB08dOTM0lE
vceni6pYt98AqcxRELLnnhLp8Iqh41eBx95OW2gugIww2iEX1RTNGiXobuZE8/hl
OzE0ydVQO+GMNJ7if5zMFQ9wPuChuttwFMzO+M/GpxwaO1C/GOHwAoyZnay5HpWC
0HoMR0oz31GHosgSsa6MxjoElqJBJ4oPDr1eRK6HTXxwkw70QHHgKMw3wL/YRnEN
KEHbZZ3PI0udhn3mA+70lv0aQHQ2gX7YyhKy/aDNSOmUN2BHMukb6JISePzmdyrC
s8hEGgIIUvai3bIwW4vwCDUGBnHiSI5oY4/jYk/muajIy3UdjshaQoC4Snlv3Yjz
2EuoCtc5/JOfOjb9jvLI7o6XF0lne/yVC0AL0FlM8Y6DYQxxWr4rj0GFobXuZdj0
SVx3S85r71uqt9Pm7xKVCKgvCD7bZaNlQx0Vx/nzsI4NUjHbdar5y6BiIwJMqsFo
dHb/5r+9WIYNa97iY+POEYYFituCCvlO/lIAf821sZIZAHtqcBbmVjIPhVfJX5mz
zPLs1VPE4kfcknYUxStBrktqRoRaegCcNsazW1UmwdmkcIj/jLRmv2u6i0+KX91b
/RPY0vhq7I0tvGgPU7HcxehswZpWEvbXmMEjksvp+Ds9nwJcIxDaofTIonOL0kd9
NxBTKZro1HF0rQ0jwl6cjzQxeFOrzFcZlIqU/aya43/HJJs/byeCj3ZFAqYM3DEK
7yMPliPzWa8msH7JWCyCFsj0EunRlmh5mbMY+Vx293XjxXS3kgiBbEosDcLipgfy
BYJxif1Dq/3ThGd+alGIkVcm8bRb9pBck31H5wZtZP/qCNTFbPULYsdVXkIxQ9jF
nZZQwLn3hQcMKDEOl807y6+9+L+FZ5GqDjw326gVH5eZq45Fu6oNI+izk0VNlSck
iDxvAQ1BHWDTm+2TV2H0XQGa39SNHC8Xz/QQAMmfTFWw1xDKJ336gGiaR6SOI9xS
oVkkH53Lvy+qnRQDHaVdkA9zuXOpjsoDsSwXN1hNiOPt+2pz9pzohOzlX1D60ppl
vOW0/Qz2ka/hTlTkK7d66le7this8N5p2BlEDuwgnJY7EZl6n5PvPccRciGbG/4U
xBrpQ2CLuOaV1ZUgMf0h4hqkHObhAb5cjhd6sd6UF0Zh58Cb56ZNPRWHqhtx2ABU
ehD36Qqoztu3ZI+tgOyjNTMb7GZ+bjSC7p9VtKQYAIRt1HjeKma1LYOQTAO2r88Y
7Hdx/Sn3kFWPlMqSisAqBae/Ncy3rsQwxPel1wk6B41ANRty7Zkar1s6rEE65vN3
Z+klyfU2KW+3DPpw5if5RPF3dWfbae1mkdMf8jogibeF+3rFdc/aQBIluunJttjh
uwhQ62H98cB820BdpchEaGAVHLctl0WwFOWHM2T/tClBM/9S8BJp/fSEnU8d7g4r
acpqtY6ikuMh6omwOY8f74u+NftcZC5zmWv01GoYY9FpJascxgUiL43R64wA3yWp
itgbglw4DQ/5cuE9+UbKB3Z3w1fUMDMGolZn9EfVb5d5t+3usDaweYlGsuHg6Frc
jZ/T7BMU9r7yiET2RfgoXQg7BjNGmOEOcycJjatX/N21hmKdxSD7nnEqRzRUBusg
yO+OSBc5vLWsW3eQAJUihTbQCNwt7P3XWDFgH9WIh0B1EjttLKrimwktJZ6A69jV
Noagfh8Uw62R685YynVMC9u5kRyOz4N6V2RP1rFKwr1jMyT5Atrg42acHXH0q3Gy
0JVXf248yqtc+lic8TdO4bIQVXR54BzmcuLHMHbRLzSKBCCDyBcXzbZLsWf2wgsL
sizpV1Nl1SXG5x2it00JsX+nsZcaPMvoIN6ermOMtSCSID5NW47eMYVdXy7GXxP2
NJ0ozhw11Zo/goN1Qn5mUwleYFK0n6FZ/aVc7mv5f4eT1iGUDL1YtIsKesKLx0Df
XsvP2ZzbOKH/pvzWtfluoVl3ikyuU6SAWRpQXQBEv/RAssMYldOuRcHy3uc1jgoX
/fESaNDYdFE6e7Woz/uVL+hKAC2Lzz9WNisud/9jVXu1Qt95GXsAK/LUtDYJ1WJ9
AhfA9JbzbHShBTX9C6nCzyC4OBJJpPGAgvQq960nQt/WtjAIAzhoKukbVjNUgnYC
0yI6iL14DbExkZmpvSzcQf+vnqlD+ZZ1QymEIoIaOzses5++eMMv34anVfHyazQQ
sp4gJCnEOQJDBv6cf8oHiYEqmEM/tb/ZkhxV3SAY4l2t8jEhFIMOwOeTPQaJcXil
5UvcSmZNSp8bPVYSnFatK2e0ulw5MMJMH5MoF6Em6OQMNfAWqettHVT0Rdxoz7Tp
b2amyd7voX3K5X8M00HNmLaYAlinNiJVf9yKD7vA4nHub5s/3+YY6clHhA0irwmb
iaaWMmYTEBxhgSq0R8Msox5gmWRuHaYwhvEuOd8qjSKV7QPu22W7zGqjr2bzpimZ
bwMWaxUypLBuxDZO0EfQIGPhbKirg26oVp28gOv8wpG3KoOS13tL95KRJMDTwpHs
hSXetmHRhMLOcWy0FU77t1dg3iU83HFH9wvZYZ2DLdHHYCXJ5gspqk3+cAhlissm
QQEewpLYm/1xJrx7KJjq58FU+CS9sUNweNBxa1Kkozr2LswXeVuN4jvbWuAxLqKv
u1NiIoj2/E/4nYfmMe6JSkKkM8lAWIbPwDudykV9Av6fDR2o58tDWVIvqdinXabn
XTq1nNHYbYRaXA4F7gLAGML7fHItPYFEQGFP2f5Qp4hr77o0WqrCF6kT6LaSBh99
2kiYIuj81020An+W32zVRcc38l2sOOLpMeAKjJ4Ik3HcIBMpMYy0CFszn/V+hQIL
8lCXTlQMFQ19VTS28hlZADz4NiacyiCJMNMI2f6GdHu+rpHgbF80Ssz5wLBR6xpI
U4zOOelorWrpfB3YevxRP7Mc1wjEoQXmIg4VyPigtpl0hirM4u1iVCkBxTuJBSrZ
8XdbFpwKoAqTiCXsTciH4Rh3Ca+WzvBDLUXFH/2PQ63MKEA048Q6ROpvzixwDBZB
le+uur3aaXmCgrIjP2bzQd7hrImyeexxMqsRuF/GL0ykWi0aTvw6qpwOw46EpaOS
/Pnd3Xz8/yFBOuY2OCs1OHsMn4XVc+VGEf6Z0AfJttg5TDC7Z3nS1lcrstt/TPDs
RScuIjzf7cnAWtO1FSCMwZk1oRzp20R9KzwU7Y1kb6PqnKY793+7b1cf/XALZcxO
+BEdVX0hsZ8WfCrEzL9yPo0fKtG5mYLK46kycp4yWJDaqjxvuk0fLZmbI1bsAOE3
QhQwXVj5rcQ+xvtok488PM5lkYBRciYqEsnbCHvgt/gR1oErNQf7iinTOEt5EEwi
b8R9eVwd2ActPjJ98cdRIbCwD1ZPaeGqW0dSISJLGejYgc5VjPKaXSwIQwyMTPUG
yICagmRYv6sjISUllrSnaBqXy7OO1B7dePoPP7W11ygy42zm88IVabhmjMC7UYoq
aDAV40xiy/oA3winmH8ftstvny1EzXub93kRUyFLBZ+PJ364OJCUpJbEVj8eiIfi
2I2i2A1EZoUVmDfo6q+Iqbh5iBZ15v+g3MwFKxfl3O4TFL/0k4sq1V9GmfPMvAh8
HOJv0JCTQTUDT6+QOqdYRkvqi1/U2gga5cJZxZPsdNgXeCat/yr0S6vL3NLTw/ia
wOpnjYYzwaGRMq/bIuobfLFHyp8id5Qh8FeDrMuYgHqrJPS7ZYzOguYRtT3Xqbnz
5isbQNDqjAzLd4FvAtXq8MBN9QJDqod3EywxpHHzHnnCVLLhCEaQJ9Vhb8kniCHM
lMWrxI0xPntWBFKPVMLtgfe8rSDKVT+84OMdCdP+2yLzDk3hNuNz3xKpkJXcAqqs
MEjjQd5RqaEZdLDHVXGlNKm6p37dVXpqB1v7QMHTWzk7CqhX2uFCwsdFawPotgwF
6NmBtI0Ck8aGOdpSXqPuUXZpqUj+zmjXyb02byBixgSG6IJgR1yo5lJPqHlXh+Sh
bgPTY9mOrlWP3yUSu/AaIQfDb9n7yoZubeKwMtf4TH0R3FH/yRTRwn22Q493f9eP
gaWC2Pj8u9vJHBG3Ci9Vd3zlvcsfgrQhmK51vU/W8oeWc0QPNgnUI6c0uUPLMHeL
tolsJzpnuuolEKGZLMk14h/MXbYUpvF/IskVQ1i2UxsmLAOIMdhsQIL36dHdYEFV
IxIBkZvNVMyy+bHGE0rnuEUh99dAwsFX49cOjS8FjvbcdpIGvsLshfWFgwY0qI80
NiWvR/45n31G7wg23Igwb1ldj+yKFLehSMR9VXZxHJfjgknDcrJ1Wo+oM3zTr7Hp
pStff5KEhErENQ+jx8CqGf+f8vhIQy+UKbtCuHYCTXpeDLQcOjKLNHOHCGIJUZfy
TOIctGuT7srB4Afz7AtQCYYwkVoY4c+tdysbE/LjUJr7CXRY+R9lUH1Lc0wjLB6l
Mu82Y+SjrQ5B4DK8dhwZD+ZaGSYVJmH1aPdXCFPrU5XqS0rUPkpdZmu4sXf8Fj9h
pb1DBe292xmXZsLDIJleuu6WvJpbTrYnpC5aalBQNHS9N6DPZeSEQ3HcPfat9hfI
kpVJVQspG83pfqHIOqQ1Vc+AygkrpuwlLSjG2j7IzPO63aK5in7t7SyRLnoidavL
aehacjkGNW0HauZ6k9iUYi2P1feAP7K8iHFDO2m0PI6WS1Sz3LXoktMnDIRki86H
naax8ezfk5Ff4hG1n4mrDBU3Cyn8tP0g0yo8lMVDl8pwXh1Ku3/3CWC5wqVTyVzl
pUPWlx/LLbcppCANDxdikdywT5ZMR+zEF3pnYXSgnMgTkpJlnavOlqqkxDn8y4Oo
Lz4JM/FmU8YBew0f1f9+odwXLV8ZollGrVCdby6zf/nmwsQ4WMcwkVe4NP9WigmD
WX1yIJUZrZNAqqPhXu2fwF2dQXa/4yFIJnTQ/Cjavk+BMrr4gFWivPXxlMGwi4oq
UtlCCP6Pw3JIaQ2m1Mg7Evtn73c3BWe0I7/FYJTWyoImdu7fCJuPgeo3RkghDQOK
DVT+jj5/kSlKPa/kqWqH/8dD2ezBtNS38E75PxKg4pOwTOAoqfpbCQygN6XUNreD
7e6WYlcs370qNcTqjKOs/pA3WPd561VEZlCa7sgfNxvPoPWqrXUOo6SgwTJvgBrh
dbK7mlfZ/r7mLWpjNkTkN1CwiBvopPWnmo1SeEIxX9gkTD8mhH/MGCkxkFuWtQ1i
cFTyyQQQ1bgDVa8EMRGJCI0fwT3lb7bHtePALLgnYrtuRWJPc369nZSLEw3HgEqT
tbxnHKEVZVVqnY/JMNg3v9cz12UoAW1ZEjjnmnMebpngmlV9fYMJ/GEZGqwByQvG
DeSp35yjsRP/rPyJy5qIv2uxnfdtzjfr1RuUjlL2j7YyxKzt+U2Z3FHid1XJAzyJ
xlrpGk32nLM93vYVfF/5Sd9RgVOuOpmEz2kyMnue8QmrSYQwPXYlQe4uFWLPuAOZ
2gxsveDp2VfkcEAJkdg13uL3A50tPQxiSYYun+csABycdyeng1pd5YzUHSLAv6qD
74yWrrVUEyoSRo9ttxE2FMxLG16WcGK4yGlMZooetsdDUgjtRW/eXIGXI7+y9hBh
eyP6AvMuUZ1UepAZl7g3mV4sWJS36F9HXqDO+G/qTzWHpzN4YpkWRA0myWMmxRCZ
SA5zD1Vp9TuKLGAbqqyutsRhejp1/gD3spxVMwtkCodk9syqYbScgImi54hPSyun
/CBmmKE8jh29vTtI2dqbYkT7poYAzaHCdwftQBHp1YP8PWSWL6XYbZYYRnBYuBjQ
DyrXkoNiIeYHUAfOz9erXH5G1ZfMcL1i6QzAxaeWJvToLeVCUasf2COlmgEJuMcR
xETF1z8/vQJjV0jM6Ot6s8hXm1kxkfRW689eS0mjCFGHJJLMUgOiYcdFDsymbIV8
Nd0vDoyMoBmdI0ysptAXFAcpnNbG+FCzcaR47w818UhoyF4ZAAPjSUmfC0k5eph3
CNrSv5mlVu7MvGbVXCL5u7UftHECq3S3o6yDfkBxRVNVxt6OPvSo/i3AJuitdwGg
KndhecyO4nH4zXuAYCSAG1I+En+G0yQT0mDDhltD8MPa2POT2KHWbax1ExVYo/Xn
LbmoyfIhwMspal1CnYg3k4cz5HVNYPTsuWYktvzM7UHPqJCUVq6Po3bx8lqhR12y
Iyc3qPas1ykE9Ka8FBGmtAwOm52bZDUlKCUbXFI2uj/Wi5MrZpDRzgI0+pRqcBs1
qJSl+MPWW3lC4t8BatHajCS+HDoJ26Lso9PowUNgKH22nIUO6yPN2oZantx0HeFK
9Hcz7/Wwl4ivSI71jMlDvPjGFECerNoHpOR+CeXfsM4bK/iX96X9QfGfzN2I8rNs
6YkxG24gaYd/da/Uri6AVqgYU9NoVnT86v0MR3bcTSO1sJesa6sXAdvk04DKmqmZ
NC91uT7vINvBtWNCQaqKgijwHdZQSr4xdif2s0hx9xjPc7y4rQrbBbjICrJwZcH6
7JK5RYlQWMpgzM+gjSFBJMwL2hgWWLTdDoYK+tm4SbwcEo9dZbizCA0sEnYOs942
QHkIt8LJsCHI5yTgD/gzCbeKSkNI0SeHg4vrj5vHh5IDLDg7wcMLlhICP83TtLZd
xGS6rexgXYo8NbEAOMDotIvAr7cYMpcNQ11KhKmrU0oIwWTDFt2MzUFjwNL6IGzj
0XmSmnkDtt0b1WEsh9xiiBJzSZbxn2KbWuxCuB+6W2p+LSjItadrZw3JLEDIQnyS
/XSy/2re0tWIbPVtUapFra1ZwvtREzH+e/jt5GZUCrkFlQdDZJvbkaU53m2ouEg0
maSkJpgqxtUh4149x1ubVQLU+zJ5DeJ8EugqKKfUPEL5HIJEDuuvU2RnnvrMUyWu
uAHoEx+O2s3xHOdR9vE+Mcm1NHcNSGOtSZMfJwH7CV7Jq5wZWuK/RmdJmKeySNv5
1QdP9UUDmxPiZjVzQIYy4ICXO7lQvFi/Wy3njnf8fTld2nT/Ep1bQH0d697GdY8S
PNYqTsmlG6rc49679jovMxKjtsXCf/LA73qeyekPe78P8foN41P2pR9pCPlNwS1M
SxEr57mo9U5YyE2fV6Wsr+ovbIl3TUVNBJUmAm8WM6O3IRHrhzTigOtn0Fk1AmMy
biJheooBoRIheXM/tQCw77de0SnjIdjpTzQtwYaD/AUUvpGxSKQCQQOocNW1e0Qt
WRICnr4EsG7dMdU98RySTQ+edzdoEeKyps6o5mBGbtFr3XUkLq4v8xLfecaCZM2K
/q4Of7hpMlybJFn6xTBN69PLfV7U1i4eCa1WfSnv1UMvxU2og36XX0px0B6siHa8
dPYcVjDVo459FVGed1gHWi0pSYhTiOaOEUr/iD+w74mOAjY+utiO6cnj/287oMkg
rjv+/A1jPCXSYMse9QBCgP84qh3A7hhriTnbXslGSvJsYxKv1JW94PgyZxrdKicy
tO4tEnAF3Mwsj2q1hdVIJZi3IHWTUUpkNns+MUGaORWWwPX5UZFoPbj16K3aNJ4j
JYMK7+yNzNBFHh262MTRt6UGUrlsSX2O01n4a+t5qJyQuKyfouIr7C4FKB5nmDKf
uwAh4kVWlZbCa4C4HMY1572DZXbwIIcO0Jv3DcyyReyLyybcjcYnpS8h5MrEHqxk
GNGkCALeXCdlmKROJLnddkIgk1BaOgZev6yzIxEUsgAXnQOT65wj4mY2muqJD4b+
KNLBx3KKJ4ErN9Pdoq+flkIGufKcJmp7DGaC8ZXHVz+4eelZVErsY7htk6oujQ6x
OczRvnatN+/xGPh/DTRFVsToznL/M2P9PHBtYrtauAl7Qsp7E5RrsLJ4KwDnS9Kd
Y9UURiD7mGekmTuAKRrNJhFWrZySw+yUr9Ktr2mpwFitPJ1O9lQxhFS2EldEqPOO
H1kSkE+yWBbqjJ+moSohdM3G45OeFncNb/UWBxjmziyTX5yW6wj7mKOr97BM2gHC
939NISWj4mqcSADJM06ELpD5G0uVUvJJwwR2uTbcKlaltyjJgfFjF9k7WEDMN4fy
WMX3OJEcpxJAauDikLThrBuWGjL7Hv9ZIMD6nnpG05MvXiH7TKzWC34IkrVJZc8d
8OamtauADbem6xTefBIB+iSCiucgV93nRjnFVYUL0I5Mzs34slLGb42sYgsn6PUy
8FO2LVi2++vIhCyKHCdSIWauk23GL2/NGnWDUF+9KiMYjFR/BdmkCg5Zj9gPwnS8
AgUEU9k8HaHbgfe3cuqEPujzR+mxxKaD7gFZOdvaCfkKQpR3gfcizFuXZGqlrdXN
B0CpiF0+XENheumeYlcyycVhXkPR6q7lF4itwfaMfA2QMLmbJqJaIjacKSEUXWz1
hmchYdfYusg52y6Dk8qxDDq7yLyOZHtpBYBXTekQS/doBTeXgERhVSIplcCMpNvh
I11chEQ0ZGWNSn2O4YmILjgDmKk+I/wmK3a8bKBUK9fzLA1GjD4SUa3u2Whkk6Tz
08ybaoBD6q0K1bpRYDDTuhm4yA9ayshTBo46f/TBUdECPqyhEPT5710JDoK34igH
mLY1XIqqL8DBluTustIOJ0egZoBT56CRLazRNdbdwRmkDN/jxWyaw6AGou28WqdU
iSLMk0XuoTwz29FhnaUqV60ve6c8qzOVLM9X3Jj0ivLGjbRwbsaO2mR0FhzyCGt7
eysc4qvtLBC70YU/1rPLICZL0/61Vj1ZSSeKPxft5Tb/KWGLMb7MypG/FrF7DmNr
j8qkfF2PRGQAcTv67hjaNFUVsCi1/17nloElVz5QOivG3J/6U9g5UGhEWHcjtyBQ
BShYYsnGGAWs5umlXzkutgRsdSQCF5pmdaQvGn+P8VAjQATyAJuktfIbBvm7kci1
gg4k2bGTlhrPXU2CRojggjSWljep67NQuGeniECJBAcHSsHuoL8UTCS6l/OVM7w9
uqa792TyK7XDh+gxKpItEKR4Dc4nIsPOuiPgBJUS131d2N5cT3hDTyRkoEA/f1B7
LpOD25yP33XCsSrrOe/w92wot9qAi+8cdnojcfweBD4TcLrVaM0DsZ32xGICCSFA
Q+fwd7qcIEremGmBRqoX4U5Bj3IKe6ViiAZIy9exLr2h/qKef0iYI2BxT/sfzYzq
uTyO0ynDI+mgyLuiCFfqFucGIQPqGU2H1tMDqOXXts1Pb68/Y75/HxlPR5r8KFCN
447UU6Ex+LNAyZwHET7rZjC+fqQP2Zulm8Su9a19BnMn2uz1vGrniFtpJ4jREJoS
2DsVRmyVSDRb8wDTO81r1Ihis5s2+wIvDnI8V3/Lwbqr/HD4jj9lJVWhBMy/Q7yI
vW0ApG7xcL/Ba+jHdQc7mA0Xlb/mYpw1O1HCho+MuMWCaFNoj3Po8XdXmEmtI+au
1wAFIrJpdM0/f3JZGl8OVJMa8KHdGoIhDFVYIQJUpf5mnhKLx9l//wVr5e4FUsgt
gnXDM4fKK2RMTNNV7T0mCVaahsE9wZdmROsomEEiiDI7i/j4nyS4Wgc86p5nb9gA
7dce2EU/cn751MMCGmH1hFIWXV8IgsOaJHZk4FzIg3O8kVsjG3l5gSvtvKT0YMQ3
eOIIfMoQkygJy/Vt5WGIIpM5KXvrSjAAsd9eIOWRAResWKtsOy5Q2vWjFEwxVfCJ
ry0CegmNWzMkLTsMcKbXX94gPNvUvbnLmRDAu0QLChzcS0wwCXuW5BscnUf3i7FK
RXYhAzOv6j/zvLLCLOqopREtiJwT/IdiCXZZgwNe81XrGJL/AvZuZESamiPQTTTo
7pG+74J0V3a/aiaetKkf0s+c8aBbh4hIX1G6DQ1TbH1giAIC5xdJIH/nGYYSXNgg
PvG6s69E70fkBwLNRcvi3ziXEuVYTN9aFTsOQFD+7YJhAkTdmebci7o2auacKlZY
bwKrJQ7HlxAFADvtpIRFISP4jiNxPbZk9VSenS4u2jtVHUHuBa2wEf10fl1+fbU4
Ia9iesCdRGgonxhBGxAwfuRhF0yuLtDxiSaLTSTeHCwHsJ9h5W+NLWXZcrP7vkp1
fGryA8mBMDAUz/dEVioWNPeeaV/ZrQ5Gi9ZGIMiRSKXEv2beZkX2wVNkN5iGXIgh
4Yu0+8qkYgHOsMkU6ZPu935Cuh1s1M/5SncpwBa2Q2nFcaE6jN2lRWK4Z8LM2Ogj
GOF3iRtcGK0eKJE2Ucf69TdMkz1nBSXYsXgLqxN930gMPrnTuzLjw15ll8H3kDgR
iipm1zTzOCsYPsJOqhrSpH0KFz27RQh/J7ZbiFa8rkeR+2M/kM6VH/VwToVvwA0Y
Rp6fk1Ef4kPKjqeMlAaaDuPReG/jYq9xBVY/FW6MDqSBXVa62GIefrU4jmlMhWVl
ZUV/id/QpCxszLdv90pFr7Ud4SbdixdzwKAsnN90iOCgxbfc7PEcjqPTSc+z+Q1X
sggdHmZsiFpErIkuQY8de35ryxasAGGcUnCx8RtK/A2GfGv6+gDNDBCS8Oo0u5kg
QO5hTz3NKZCFadMwAP4uqU3tjFHCp6rLmCJ72WCqGFpBDVm56fEBYARbUwJ8HAV4
k2XV55LAedO2redYW3uy4okCL8+x4Jr8sf8BLQ4p4HzzRNwaIbHC10Ve8oIDDEJX
INTLn6BWYgg87n/Xtn9Fb4sufASx9nJwy5C9Iwg1lTM56rxxT90oKwmdmQjf72Fa
EoOwuQWsqforCGkpgaiZ0Pble6UsN7y7u8zQotvO7xJ9oqIj8oIa4MwROdJhKfMK
9ZNrRX7av5Fq4viIDg3+/EVaWLOdtFvcy/7QIj+WzI5dOch8/Jzgdi/a/CYmOe9v
QN+pJeCfRKZfC1MicgFccHMNLD+UkfBOWCH/cncL2wJr3gN5o5ACff75GR7eAQ/m
qSZzjum30VKOj+296PVR4sd0doBMlFsMQiliOjrboj0xqCJyF1I68GlfEXIpd+1E
Ze7hLXaFU05NQWKtAFP3kw48YD6qjJ1N7ebMO1fZn435aMrS8vGklLpu/gb4e2xZ
/EH7puz16vGIMNDZpFm16tkNOb0O7mY/3en1q+veh32WeGo3by5NrGEQgv2FEolo
KjRxvRNGdAP5nb3cshsbt5kQy4Y6rOEdtabl5h7JI2gwJ5qTRRPetxos+BOnc+DG
22BRKau/G7+Pl7FrB9mdxE4kS5nVlNYMXjtQs90tyASOUtZlQuMrNxHoVQqbwxvs
IvF10HrW9fXwGdEZPyph40CWVX0lEh/0yGW6gnLcpwdCWyeYn4+bwfFVC952aThO
H63h27vW2ZisiFjJSJDJIfcsupi7QmhDoTvzVWO9cmKYK7IJtUVSRbzAKXO9xp64
f1rw3+UmmDk8UueIlEFnnzDvxDasfIXZ1TXweQI9nKxpWzeNcU9u0iyANgPEgXPK
6JvLM8OYKgpHzJ+czaDot7w9IGZ/rO50qTBvJO097XYcVV1RBywTpohmV30AKeWv
tjeT8/aWQlX9VuNxnD0C/sp3Rfo49Udn+A/6De/5cQjlDNCVO0e44MqRkpKuCx7x
adVSsNcN0No9t0h/a+iTfMGLurrB5zCuv7SszYzPrrZlXPSmTUIS99BrpFHZ4zUA
LH0z8HjtQdrr98wIq9P+MA6gkDPZR6zDzgzFPv8PoTH+K0U05VBfG4ja05X+VxcJ
g/yAoWBC//EK37A1rf3OFXnzdUuPBfLHX1sR79JnkggmHemR54pbsOUloHzC29WQ
eJKGdOyeM06fN1f7vXF5u2Js82YX1lBG8urlD32evhlN0qEACyr9tUmWfPtdpGRo
3WHjJPqguOaqoPyZb9CpIzeBO4eJTeIMk+9cjswGZmg7tqb6akRTQQYw/fkvYNmm
9/Rv0MM1xUpm0ImJIgjqSVLMD4lDNm+6iJnNYMo1fDY/ayD509tP4E/MmlSLdNuo
zdskIcKfQJPavBawr6czmLqNTDDxRfJyln7b3caF0K/fSeKxYIYOvQbM45iATpob
HQCovlPqFtvcDxYvEO7OiSxt0Ztohi6RpBT4SevAYY3ThDnsoTRABkTcL14uDFEl
uSUTvkczqg/GPOIFojsMAsu5HyqNdWsDdkIiTaD9s07RJK3X4UAXeqVUaUaoWs4r
BZ9znSk93FtOotctKNFuEtULF97HuPYEWP6mrBwVjguXOSVvdxU+jpm5RgNd7F6e
7v7CAZ2VFP/zN4AbGGJY8poPA7CA/+O/k2Pn4hdF/mnn41/YssLg++t26V5zGUZD
BczXw7CW4DSyTsyupu2V5lX5WHe0gFTHplX8FkVitVflDkGdLy7+qriCm9Zi7l7D
RdNtBI4JiPz6JBycCs08EjA/nDnohvclsWGJRTNHptmpyFQCI7uC9nRqpDGnlnae
sj28kOPo6C7gyCY6D8+UMGt155ammc1fNE1KiF0aTE5VIzgIiCkv0akl2MtbgN+s
RVTra2+7kQJvQHbfy28mJn8zSSjEd7blZasgt7BOkc008g6lSTUE2BftmTIlMQW8
Z8TTxkWIBCgxxFjFHJcBkNOSZxLNKLyYgcVM6VYGSYXqjL7VkVU4d3mprbKbLo9C
fqKE6hZnbra5Il5cZ+GhdhpcxcVq6i0YIesqJILUYmxzIVwSNWHbuXKmZWLoJo0H
lPgjZPwGH/a3ZyOqQCowPL6P4k93NH4eT2QhzULkNS+Yi7JAo60P+a2Y8xBbM7Tk
6bBXXB8UR8/YsXwljy6Cx7BhZWt50WHOd0tc8bhoVrwkwOqgGbKEWP+2s7os99s5
nORRlP9rLNwPWcT3BFk0HbyUtCshU8m6M77W0PxsfyMyD+GthVMCurtlfCSUSMV/
txazDCPMHD/8JMa/G4VgGm8v9aUW2AI3kHK2Ye+AM5CjvmZGwtTDBbVju2MhRhkr
tEqIqk8ui80YsF8mYB2AAtbiRAwBLDq9hOlPt59kiJz9OqbxmWQ/zvIDBxt238Jt
7NmYUocRwylQdPpphah1HlNHn1mjJ/WldeNY8lUNAaYSbItXHRfL+30ZujF6IVj7
ULu8kuJ/usoJNW0ipVUTvtUCO6KmISqoWRGLo/i6a1sKwQOny6DdsnuO7gwHtavW
TaFApj1O5yr2lukTSBzPvnJahO5xUM0TVrwaCacH+pVgIibv51Fgsd2ur73fwGG3
NVaackOHYDf8HT1jyAvryDQtlMoo6hElNJEHCW9eOo91jhbEDAV7b5vIANPwps/g
jjspxVKnUO1FNJ1/8iDf94SMeFn6mkDI5Rt3Gww8V5uDA+dvuACrW1AsKP+CcwQZ
jCiQ5ZcJp6U0Js/w2XLKbAxmH6Se2KU47oM+69VgoFTdgvJG/NsrpgoZjoKO9+AQ
8cD2VLIki1lGFSLQSnBdUb1lWv7CUGGyMoGMHYNxz4W3lMAOajRx9KDy25ErZU2z
dlEK0M+z3DajhrPfzxFk9PERSn/rs4u6aRI950qb0oPOv4aO2VOG/nM/jT1qOYmO
7JnPmZd3ccShTRDIurxhjMehF5IZCSVbOIPc3POoh29dtfOJXAxJj0OvY9/Q1ukI
SxQLLclag1xM+factdimD0Mqx91paDGMQVWBDNvcFpWTOQxL3kMfAbizgqsTvPJz
gqkxr+J+r4hvnc8Fja11Luo3xxrbPAgZWZt8Tn6eMlC2Q/EbW+EhKcCnsPo+vqiy
qmyZcCwbXFONcyuoGbxHiPKwgC5TJ+zuojcION5FreYI/kRShvJauzlnHNszqceg
/plcI0m3NkL8PVwwSnz7YmmLTDlLYmcrNzzWwgXcwVu3F0pMapq74G8awrIqnqcE
8O8pmn6B4UODiJzzYw7tKyN6PcefIlKFVjyprRxWvItLGfTH92pAq6lEnPyp8Xdl
SkGCsOxs33iDK1Egeh941rZqF6z30TS3EUmoIqOfsxIV6ezEDsQk677effyhn+mu
1iX7PI1J1XyYxoZEHbstQ4P6S70fBe33dAeSV5RmiXAGr/f5Jg4V3Wli3zQ0PX2R
mysq0K9t52FeNFhey2R7q8xK4bIV6r66nnX6lMIWvkRtpLYbPZVoT8LNRVMgp0s4
cPhxKg5Vgk8T4u1rXq1piRlJoRfdF6apOKSghvs9/Oii5yErF4EVc0elsUQA2rgk
fCyZR9CgpLt60XyBu6Ug+ugaTod/18U5HLZFHdzCEzvuOH+BRL2reWmPaeVAqypj
t9oG4L03lQv9cSUGegyFRMdorwrORnPG/9ks1W3FI6uE6IWwfMr1wy7Kpif8NrEX
Cvio4P9ruhsgE53nUKHqU0iduEoFF9bujDBFOVCupnyXlYg8mnFagy6fojz7CSLK
ka/BCCOOovuRQlIRgjsY4fGorzVDi6LVNaLPMrxAw92d7DbBV224VXK8f8h+lti/
dk6qweLmuJTQryTxQpuHwQzT2BReUfEBmZvbYVvdYnXpvse/GN72byttGe4L5Mcm
oB4tyMKjEg5jKHPtJ1BBZeVh/w+j2Cmgwg8iS4SrRBITrvstYEf2OBZTuNljzovr
fxzOx1k3uEDk/+8OQN6r7RMlZfr3yFc9kPRM7P7hYBrZdJ5tBcgeWui499MZU6eU
/JSTuI0Y0HfqlNcH4h9QR24nXNRn5YC+9OmP2a7ZiaaAPr//NXpx1V5rhRIngNgD
KJotMWxSIRpzGZscpSwaBjD7xk9f6F1yg0u4sptKd4eL9SSOgNfQoQfOEYJ2VrZD
9jQ9XER478ALTou1Mqjb+gIT5O8E+8VZ9S8aEKcVRA/rTzVcsCPYQ1sayfHBfCQT
WH7tfnd5ljM0HWUhjwt4QTulJtr4P8QhQ9B/+UyTLXjnqTY+TXnN+gsSN/YQqFOf
WagaZldsZcXKXSaWENXssq4/8RJyzPyJELcwVTfMBqaxFa85DkrYo4pkt/NIIfWe
T9TQnQj04h5T3knSV9Dm+t66td9X3pz2qW5y7oPahLijpSplAl3fVa8xep0tacbM
Pi6Kvx/9wn9ttieCLmOkaWs6Lzj+zely6V3yoXbZL/T8JgYBjkxKBND+jSltROS2
YTsdmVlYG9Lq4rW9+JMHcg8G0rC7MM83OtOktosQhQx6/dd8YlJk+SmJeNENk5WW
C5qUv3VrOrlJ/xgIsaaV/hm6wtY6q780QVwIHKnNem78f5Xe/tPdQelmocEmiUpc
Q/YsBxKJ4+LU89IiXPca8LqD7MdEZ9G226OeOUgiIba8+hwGrK1x0tCJrJlr71Kq
Z30gMiZF+zRrEhjsF+PK8CcHHlSR3/+SV88cPPbj7ELKbzgkHhdhzsUnbR5/C6jY
bxINYyh7P0eL9wUhyEXGjePzWEdOntyFlSFiZPcXZtEGyxMdB2xjd2m7q+kOcXVC
IOTK9LrISgkusvlu7SXSQnap649GDHXwggZXjzbIx/1TOz9dvJhbsVu03nVerhfk
qWksXyojfwtCAnM6RWaC682GEnoxAj6g9tJQ5XHbXyxrRNKM1jLva8wHKkk0YtXj
ePH9f82e1sEOUWIqKLhhEVBY05OGb9PXToZx6LfHNSfR07MCIhih/2/BYkio6HAl
lEDSaOLMQI7Lf0I5wgTE+S8K/MsMZIFhhDiBm22TM10eCzpK8d38S81um+tsofdc
8onuTIQ7p3Ye3uoGKPOXo4yIHhu9ERHn91IfZEBkhKZJGpUxphqSm7lAaGBs2K0H
j7V1dGc5k2i1k5QhwXd9/Z/ClsB/Ii4KPX2vF2OwXQcHqiGetPbhOcid+mnKsQpQ
SuPt2df1u/08xIqgJmYRjy5d4seSJ1L6WGR/+wp4JRQI+KW/Q/g1DzuUcy2d4Lpb
aUKVvIY7UZt3mSZLQFr98dY9PxwxNucS5ayqdGNpGKdS8/gO0Oh3TzkPNsOD+gp5
pxuPJ7MT5zz/UV45Vxo+5Hi3iH3womiPsuXFyBEraea1V3V9Kgd70vGue7oWqgCd
zYKaPbypnJC5GPT/CPk9Xb9KuO3hbV/3ydPI5plWBckQ1L4GIbjSto+riyuATC1g
2D5bzvFCFwD2d69uW1e+qU344g60uxrui9ZnJE42fcO/uLyWyuYG/gV32V/N+cPo
+8V1EnG+CXf0dl5VRgJDdsEBLuusjt44cxZyIEWFTdnjXtym8pbdZvL5cW9yr1zh
HP/HWz8dNLiaHeOzlxZURCVT/6qVj108+SxLNMBDFgoJXHJoi6K4x+9sZdjM6rWs
bmlGKJTVf+d2qYZO2qiZXhw7R/1HDtT+x0ZG3RCAuNEzlmhb9YBcfy27YzGltd80
Uf3PbP/rn2mV7ihxzGKaom7V++l39S8gphc6lGn9hDkvgwNKcL1sjmDlJQKhuQJ8
1A9l/S2NsRuLNkwGvyn/8eXCKCQCJH1VRHolXeNvvK4cc+9GoT9f5lp8ojBX36j+
kGXK453+SR6B+L5alIbgfFaStJvKbO35sKXMNbri/TVeNY54+X1aN9w6wjIHf5dD
UcaX9Ja0jmODODOhKTa79s+OFT1do4mFEo3F6WR3yTzjZU1jW/lTIbjaJZQpRKNy
hwjswn+AZfCIwR7CjLttWIb2smR5dZyPMT6PloszTET/yo/Y7blZN/1gyRLJ2H7Q
rvikEV2YHGFcJ4j9CFxWJxNR4bnQx6LHmlwwwh8S8ck+bkOlK1skY3rC3lZeQ7Au
9eJm94HONF9E4Wevc6AcCj4Czj+OK3SViSyoGBvqe/m4M9BrN/3wuk5PE9hVxVA4
5W+JPduUvO1cYF39dYmCBzSxrhC479RmvpDGYOMdHsB8VtPAGv+D8JI4AmMYjqgU
kndQmooiSWvSigwDOAwxqEW9+5VzJanuBXcxZLmLOn68dQ4NbQvq5bJnP6lCN6KI
DQNdqbDfqDnBvYdSawQGGoMbO+F5PZ6yBj1oQfUEG3Ho03Plk1haomzUf1D4e0Gt
mU99DhpFrZyZXOvg0oukuTa5Jl/NfECqnjNx2+Ik7ThRjN7SBv70FGyIGgsFY9sw
Onirjwv/DT5HaeymT4C/sju0Nq4wciesGjnKv0WkaOLunQkipoNU9tFUXFxOXXqs
iZibuNpnZV0gAcsC8p3mOb8gWLnn5aZXgWG/DBpC6yf5Ux5RyKojSV/mSZ6Y+exQ
GwPe51CEI9kNliZi+F+07TL662ZfXjbuF9OZgMiB+dV21KMybQMduD//VL2Umzw/
Y1yJgEMQY/QhyZEcq2gFQhYAwDclNCmH/+xJBB6MIUyq5Byj/2yCXjWNL6R+65zB
sioSbetSssRRbobs9S0VQa+UvHLmW5jHnDT5HRakhd41KK6SzsZsVHWMDdqMZ09g
g0RLwqXmA1DF8MHbiUdJ7Jff2640ZMh3FrR5vRLkG2evvjUdcVNmYqadYCecJspi
Q48tJCqJbRXaAcLnBialtV0/c1bJDcKKIKXRnBWE1b5DjVs4NgzmqRkO9Hevy/4d
6+XI9JNh5Tt1YCbOv9Elo607h6yK2kZMDzU+pw20YTDUfZqsLlWZ6x/pO6+seJo9
BaZYz4irath4r5OyYCLBgqlvKBhYzVdIw7NpyYJzaxtYkv+8Vrd2uOc+UWSuNTe8
+LDk730xFDPvrGjguWob61g9tzeDFlLOLanunNXCPjWdMnnqOy906aPgCELeKByC
BozxU76f5t17YGrAOW6OOI+lXDGPZjlVbuLjlMcNqNqt659lGLHKWDZHdt4gq0IL
oBqnkZiCc2TGvDkHRnyLX+m3PTAkNpK8GLKBCeR6vxwNZ5+jPOuXToC7tJA3l/rS
bHbs49C18o6j1m7Y4cuoHp0noQdfi5SHxRA940iGYcdahW/wbV8cUy2yCosIjdM8
/VoHF7AOPOsmk5piuSjP1uHmiKx7iD7l5FPhYDIML9m4ueqQ/zN9+g5sFojj7RyQ
ssjy4AyOdfroxxnozh/8quEXoqPciazwDg6P7LqVTYxiUtXdiB9a+cZMI09FEbMf
tAYkM1YdRIA8fE/xA3VtLZiOfOQdSlTn9OMXvySBaumk4eNYyl9hVoV8jV0nras0
UJcFbz32ihAWDFW9vjyR6UBhQJsAlEmPOORwl9xeEYNSKl4w2GxYKTiI7+eMPbFR
pdlUt+J8AOspvyAclSrpIlZcHnWeThzqHHA9xaA5VAIB9V1qKJBn+WOu40CJvhwd
nDRqXYaqU+wkRit8i0ygFcoi4Hx3n9uBQidzseRXkVKM7NOkaYrtPwglD2XxcOZa
7iPZz1DLsymICWlXOcnJeYCMhATK8vSrW2/nIDieVBcVMuiW6jp6Kz4xN0HZIeC9
45xZPx6wYft7bwDBeQyoDR8+ZFo6rf83uL2sbZ+ltHjWjl5v9vcSkOZFuJV6UJpL
pUjV/rmceQXsk8YsRXYkgKSHD9dgs7X/Yqcj2S+Z+jvwu82bX/iy6JS7r3d8i2fC
NUzoeApWDDPhSKdYMi2cQK4CLkL9qCvJiiMgb1+Mj/UQfA9Bi0Gc/5xvjOo5He76
hKo5Xmxfmd1jDwPEhyC+B/VlLikaQEVt8VEmZLmvsQyqIxoUWJDdFZt3dcAq8U6h
kAH8baQekncr1his7CGPxndovE45gobYtVWBBsojjoft/y8bJ3Acjh+dWwK/neVH
3Pe9rj9V4Bugil2CcOlpwvW1GbFOCvSt4VClohmOhEoV53udX+6ehn7GL4p5BEy4
Pj0mIJAltrYG0OX2F9HbucwClFyG7fG+95uTU6+3LCIJb03QfMN0pCuqF/E/RGFc
Fq9+8oh2+NKNSGYPl1cImadOk7/DsfzsRxrBsmZgQp3yOsC6V2bSha/NIV18SrRl
sV4PxvSEvpKSt49hMxG0yj/nDYJ8FITjPxvymDOZgqNMYQbSoELFsVQPHincJN8q
8vKNpVlnCJdEM6RQb1uymdyVdo5sr6eYC760T/s2MOcCn/nTe/4v3oE6A3uftgU5
WQEUqLkf3dk+cdsGvQ0L5XBmij31/AmRiWdU54kVUds5PWZedGj+MjAYROdf+qXe
Qfz+2KHJre/Q2QzKOsLJEmjTkMBT+v8JPWFnxktXPhEvf6SOaxVHLKyU08sa9J/8
frInVQMfoLllhcw5dUpkLj2OL2h9fEIzP7AlicLhjP2NiGbbiUiccpB5Bxd2ptDO
IgfGr+59ds4T5a15tEXz6Af0U4wquso1MPMr9+HdxKUg1Sk7o1UgLP6s7KS+GXkb
1r5qToH3Hw25iaqK70D9xvH9YCf4H5nA4nIvAbgdmZk69WbYnBefHgVyrxSPhR0v
OIVzIsAinS6+ImyYXS8/Ct1jshLKcOVb38Jc11Xz8IOJ582vVYbg8z4T0+cHTCKG
iBCBpIz3Vv7BgSuWI+eyfPPqZSjA8aq3KsX8PotHALiZUisDF6zImZBqWtI8VRzh
X7O8XVe0d5XHcMf0Nq0lHrdOFCLnCEq1B47zU2sYDwYnMhqbCt2fu6RM1hE3f6F2
kiRw4k8Ad/EZ6WLtlIz59XtNbFSEHiEQc6KNO5FCHhcKzRx8FHi23EFALzjUYZuQ
KTNwcEcQjxNbdB2hUQdmeEVRhPfPYRmUocfeY+zSeg700B7O//wROKRe9is6nlSJ
oW/4eazYf/qa+jHVQIBV6Fiuaiq8rohaGbKLCc9Tt/EWV8WFT/V0jNKZ6egr1zCd
1yzhuH5s42tL0F5xlwo80uE/Wh2EtPLKIV1v167SRwhaunWCPZjBOFLfsH2iieNZ
MAluXkBycBKpTM27bM/Jzuf8kkbcNbz+Jz63kdBSD8VH2B5kSZfvzy5yL+VgE5kB
5HJYr4/JzMqbGVKScNlQV7OfT/x0Eyglc4swnT0GURDi8iLAoA2gTOMy2F1Kdikt
214ekeoWkVljJwwo0ysGi1ylK9nzRgTp5dMd6bQ4F0gBYFj7FLF/W48VAaTlnxEg
LuNtUSdyLr6Lsndt9LtUnUZGUnHTCSeYNkWW2oIINXUYfiN2Tp1ih5aXmKiiMZVb
iCJC3iy60JaYMMnBNAgx4E+BuZfCvA/0Sl/l4+uTmKFoGtEvHXXpBl/nqm/31NZg
hsa6XgW88bkZXS8av4DAr+QtNlm0JmDa5l1Zfa0ebc/q1414CaAgLEkQXUHRaeAb
a/7I/bL1oKyeUApGBkb/eo3z3uiWMHxn949UqLZCQsonQyrdNAlfyWVMaq7bmOl0
uUKnxbTUgmUiPvYQQupTwP1SKJWaAMUy6tYYJf9lQ9xisLQ/bGFtVLaGpxGz3kTH
wi0WlwNgWnGOqqSVR0t2CI+KgyhByPTwxownjUoqzY6kI+VknSvIp2mw/tAuHH/a
GD0bZbgOAwS97UFxeCBZjl3ZdzhZi2qpMOoln2jvthLN4LDjqMKeFQ7TFVLx5pg/
WMNNmxei3AAxLNC+2WknzDsL30llzqS3RZlbCEJW5SkIMBkDfQIJQ8NvF/keef5f
ObA1JvpXqiLRIzyJM0NKyx2yRAfTNGgNC6g/Cv3WiI9+ud2XyJbTu3YF5garLXEU
CCO+eZ3SFRNu9iR4qx5+CfZei70wFO6nGKIk2tO3862CbczwN/DF4KAJQEsF1S/c
LPeuLU1BMt22z4Wr1m6NRFiEv6NPbTrJKEAokHOj6DZGL4nYPLR7fSEBaK7sqbD7
QWnwDOerUNlU7I5x/P7w26pfVFey1UEmcugtBZFGn0mc4FiX/VGMGHdNt7GFNo7b
ImcXtoOdF8+Lod/8co/igssNAclioBH4dYpcD0BiDcdr+hPZKyEBoDPfy+2hqq6S
vG+OiI4E9E8cy2jSOMnQmIRatQO9bxGYlrHlEaWau2TFPQLQXhUQYmYvXP6Ym908
TnU7LEIAmrb8ZdvSe+NWnYthBKM416dbr20iaBHKgmvIE9kis9AHm9TNtZkLeGUx
mcN4efr2voCOKiR4oonAumaozYyo0i+Kz8hJ3mWClL7UJabSa6MbvC+ihkn32pMq
Y7m9dFwVF/aiIz/e9jrtCCGI8B193cYJtLC3/EA0NdJW3vLMjymN0v7tJvh+Jd7d
lyBGkCXzWEf9J9gLQbp4TROSNs54659kk8vId9U7NYxSYD0UILxwViInLnG8t33y
A3PbxPe5V8bLg12NxC6LrvJ9oX0YNRUphHKwrUVW8tV1/tbrAojwsvt7odtH48PF
ZUXuuev3dF9stzHk+3ygNXM84IVpOGreVQWVVrMoRBX18WaI/RezY7BC0EP24K+0
SIk8CuFYV6bpxBT+qdSlATPqyGlUAiuf0i3nVdvaaB0rVVf1L7CwZ0I5sxX7D3XS
wgkiTIHxdv3dT/1aPLKdesddhWU0VNL2TjXSJLVvlhsqDTNZYpIBvt+d3tbwRZ5w
KKYiwliw+7BX8lsLQ3BkgpOqOJzvoXCscYPb15aJKi/dpN9UYwP4bfS0SMnqMClN
VNkTUydRwuK9YpZHFh+TGBYR6dEOj2j+NRVejkd23PXbw9adOSQjWdHuA1/E1qWO
2QDFdhxg3PsYxxWcQ4MECanS65/SP/6i29yDZxjFJjgoC4EbifedQcQd2LbnuCuO
5xiol1JN9fBWHosNfYW++hbtnE/g2oyTpLjYgszUsU7aJcDhKO2gKzpoi/U9mWMs
JGEmOz6PkIATGr6whNUlE3FGTKG02wz0vtx6XLS9VfEr5EeUiS68pAK1p4GC2EnH
pZD91mm6J1UdgAtO1nJvmFhhgXNH2wAdRJB+KJOP+CQqeGHSt0KXEHdParCroRtk
WqmYCsLUbrpkQ5T1XS7HeDYRkJpSlxv0bCNJQcDhyu6Fl9dKzzpUDMt7nhAQb3bF
jZBV65Z699StlVEMQlkCMLHnjoMEOGgQGqXuSRsKgkmPs3QETYNOpnoayU8j+Uhk
jsGBVAdoKKNRu4W9fpkgfe/Ry8IfXOqPZwvwYVt4ME4G0Evqf191vAfruQ5VyMMj
BWRKrTtn7O7PIxmqRhFMuUVATINmiT7rvCswRuV0yBkqkciGRybdGvQvBI0C6fvd
/iT4/V5Fc6hYhN356oIsyuU14hCIOvnq821hU7umYIs6HmB3tHi2HqsI4rVLibj0
0k+LCthSf8aAQAOsEpbPzLYzq32OzDM2FrmEwALRQEUtorzMBc8DZaOx0Sm5oOAK
oNTz/dYUB4AclWw/cAQvtSRa4EisTJutLM2HE11L0p6gf0BAZiYQgeimi/fb1T0L
6XG4eMJYSv/i7I1ExXtg7NdZSaE7aTiGplrpJMz7Lexv9WF/sXdNOpwvRluePezo
SHP1MLsdH49MZYgO969xgDANw00eOdgHx2dLaTLEmFqr/BJ0fOoszNT2ii2fdoYu
nScd8cUOBvizAs6Ooz0V0swT1Th9MKo3nbjih2lBCRlguavmklgPetCI+rb73Nhy
SUG1wI92kmBa/RDfuQLNCwrnpPzx2sRGWhaLy6qY0zTmi6QciC54T1+KEIRpdmFL
1UIFRb4e6GS76U+vauDe9c7KXOAcXN2ObUQBxXl5Pdje3hSsJeh/0EhRTvDmSB6i
8BKzEM3CMLDLZju+CzxovzP8jWlz3G46m9VlLZV1mTJSpQgx0u15TN926ywEA+gM
pHkuvG4de/xBkKcq7splFOH/47hMHkc6qMYTspWA4LbGaku/9mAFnbm1iChDAagh
0rmxx32fa0ByrEUaXzm4xZy5j2BjZ4orSfNNBqb00moNFM4QyIpi23+o/KeplyCv
ZLTDru0HaY7U9WbTdEDpoRJFd5fdYPk6Pk/BFwRiy5O/ukIFj3Z9nmhyyueE/gpe
TbCmZDLfewT8hQph1MeX7qN2MuWecedMQ5UcOcBksgqJff7qxb28m0qgElpSw1zz
YskXuBD2qwxcBHBosY5qO0LLf9fBGaV6Xz939PspqD59t3aLfIG+SdLghA3or1SQ
7VHiCB4DAF45gLsEjzdY+yv4cVifBynne3Vyg33vH2Op0ojEpDjJCDqZIWkOz8CI
a0+seimtXxBOi9nwaJnnNKiIIG1vfdOay4dBtyMPNGVvO8uWmLQ0EcCdxi8dedeS
rnf+oxV+5cpdqDn/ch2+sP3BfI5B7gUujeyBXCl7jLWPA66p9I7/N2nmqIKyFZRE
1fLzIqh6zHtKZMMDI0v0wZnzIZyR+WhN4KRJSTxfhkCrip4Im6bIWDqa5Zf/EHbT
QCEkiR8c3jmSVzBQ5LwkY5ZkudtbPnpAQjSYa3B67N1hn6VBnKxQT9UChzslwlMf
i1QGochLQph7YC311HTwtleKosQMj9DA8omD2L9QNuLjVWg3sHd2p3P/A0Xcop37
pqeBJWDTcWib5f6rpd09cvkO5fO3n3nlfxJdw3uh4l9hvzJ4mLzXnrxb6ugemcR7
h2+QSBlBcypfSi5q54xSwURLZRAzN9xENh3XhJnz7o4YnA9kayibJfW2sbBXCJW/
OcFVJO2uEXYyM11fbu/Fsd7PTIIzopTfiZ+UsU/mZlayssXOrSFAbj5prN9aECZI
KK+nTjyPD1a9OopmWeO1D9QbSVCU9i9T1XNsR3BFeqSm1C7Nazn2kW/KtTTDxrlx
zefsSDAq9PCK2Fglhs8rPyxn6YbM1VBgvQFC66H4iccmb17BEDphcHt9EdFJLCjL
U3/VJHg++XXHpsHszQON3+2tEL45pne8JiAmSpQCgmNAF7Ehp5uwwSujZwCixgtO
ZqX2Rw37gGTRgfPmNz72b4zTM6Aww1eP8Daa4DzrwYbnswnlDxTv2+NWoeyr96sL
mMUhxwn5fx/fT59VK6hJ9BtNDuIU4Rez1lXEKjw+5cTZvJfY6n/HptDDgx+vqiNw
/hu+Eve1gEcsqK/PSYbEMfzi434b77JW8IkQT0slyYYSB59eDCMtriPTJIiYZp4w
wlFp90xXJLDKOTnjb/1tcOQsRtpbt9wXJe4v/kHXUBcNBXiR7BEEKJydq9lTVNO7
bMGN549dToQiQSjyHmX+Wbtt7/XTOwN2Olj7VFEBfu1iXn1CTjvTT9JDpG5+QzjQ
un0mLxbnjmbASoHq1Ig4lnZop5wG8mO1YJ3oaBZ4L2izvSpX8rLJf3mnNkwVazQg
ZfAZG1XG0MNTlN+EWnIa5DtM8Z5cZFu+uqoo/MLfH/+l8l4KA7VWUgI3WumZn4Kw
rCzMBkxNIb8+8RRCUWnXtjAG2ER4x6PUi3kwUXnt06AK8/DdIFe57hLMat3sBuGq
b+XunTLZK4skP0hI4DHE/z7/SMnvymvyKeagf0qkqsAEOu3Usl+lugqa+KFND1oU
Re3VzqGNj3a2f4NeMakTb5k2x3v21cE8Rj8KN5elCV5Li5lYcQueShGddQ1Dx09S
RI8JT6Dp1vGKGSJP2qivHZfcdE9q5GofDP2EyMct8ZazJg/2m3Vv5p8ODg37wi2l
sX63X9OBTaewGIznH6T2dwsN8ZB6jjTvTVvpSQpH9QSA39qOp9SRnt0UNVJc6wcD
UdfWFrpFLeROWkgBITFsocUN40TOEnU85Dp8EWLhzHn9T2XFMeN3rrkzsFZW+1Qw
Et0YnOjbuEZDu6UrkRz0aK2Rc0K8mmm6wR9SjoLcwPpYBiFRodn74XQBUO3W6Bea
kf9ESWoHHcDdgcVruk0ku7JCPch/WJIOPmLRUbyE+PQG9z4cTa2MVZMCeMjt1aBO
6elIVZ2oLbHWGU1hZhMTWA2Qg6ObLY7y9eFvHHtQg2ODiM+s2JU96Xq5NVdLg6tF
PBnvaf0jHT2N+qNMQe8rUia3e4V0DoSHiM/nH4M7gf3Uak01l4r3mtZ/SY3x/N+Q
WSEqeZ8ZnmxikyHoKaXeBjbbmf61+A/nL0w/dg0R0u8QrhuI9WHBw8FWeiZiiUCC
eoF4LOZDlTdMyNQuOHDNL1XO/n3PMwbY12TuWVPE+E+prEMpzLLcQqEXl5zBIAxO
FQz+W4A5inpyB+bSlZB6fSJYvVWS9Fw96kdvEdJQmmeHX7vKJpHk5rFVr19ONK9u
1ShmoOjPcPVJPAN7YFAiJfqdpHvYkFqakCwmuA/8fAUAr464faZPAoGKlWC9YUW+
CqY1yizSgM9KqBE9gyfxMRiaXgtpjhTkXTBucSaxlLAK+yMrhEjJPA3Al4w0AfMG
tjNsbd2PmgyNePDMHvyUumTSoIH5aeFKrC0XvgFSHVJ1xqVCYXQfrtKLD14QlqFo
fpcq/6raeFkdkrPJAervMyAfe+nskmVSQRfgetRCoHgaTyjseHMmgeJWm0g0Nbpn
59xAcKxNr70dZ4E6rM97aFJtmYqplR9KtgcCxofPyQ/vw46UKaKPVtQBcBVFa+/f
9p8jmIF8kfnm3wRjXEKGDS6zpzK5iuTVaNMA+o8farkHYMutphYtIEtsUqdE0r6d
9TZPr5Fd6qXFW9tkiMhYBet55ZS57wcNp9uwMYLAifYuTSUDulrE6oRyDphrnxVn
r4XLgn1WzBAmVnOaIlB+bFsC2oeuHBNl24YoVsvaIcP1BTI3ogE6iKnbTVJ9U/TP
ajiIJ3yDiffWmYt3XX3seWtMbQ5CIXzq5PmyHAYi3AN1tKN5MpMc4zr7DraUQGA7
D3Y7hkFMWd/jLWgFzJ77zX2nHRGOTVznVa7phTeyaPlRyjeaGaTnMIJcjrKOt/0T
4niiv8C8OPQ80tkOnxsEfmfWBi/OGLY5HrmG+FRjDpusekOfG9Xu+BvfokMxBd1Q
Ye4hZVyb9YruPQDqM1bjycBiXlsJ7evd0UOlmMua7PjGrHQvNBgQOD6sQtmtX3am
0bUWhuJaAAx02JBapdCLYQGPKYjZpVe0epCNvWkvrqbLLE4VygX+aOyguE7U9IUr
Ok6nvXsCvGrW0+cqP0gclVjRpgpcTbo2Rf+iQ7ntpQ4YRRXDcGWyOtD/WGedCKMA
Pnxztd0BthWv5ZaPoGViEeOjQhJmEzY7ICC2ANKa28LCs9+FUur0gRt0YXZMFAoF
4kv6booEOxtRauEP0oBR6EBFQtulAtxn+p84W/BPuaMWLorZEYDUyH9Jy7JNXNNo
2w6kEYQgSuL0lVIc9rw6BNdh+CghrKVHRQrffpYUESPf5mOFNry/XYyQBbzI8PBz
q7Zr7rd/FVS38fElcsbYPACrr/gDGbcmMqO0pzVxJIMtGWGkRkobgFhYb0JGDApS
/TjbZ/bilVyspuoPyPlaiA2h18h7f+mt+LUF5/+MLfFNkNvaYdneeeFaB6ogzMan
poAvvMskTmLqd9sI4HwwIR+4UdWAVJdkdh50lqVlxrARGa3y8lZicFvoz1+fnXbZ
kQpIaffW0dQzLdc8rQtB6OqPgreV+BebQXiScpXFENCNfLlAVDlmPjS0Gsnu5qw8
9G+R+KkNH5JbM3Cp8vx/Eet5JGEsscC6gA64b3W+EJQcf1tuMSRFnNLMsu40Iynn
DnFRz2I3FL2G/LPbWaK1KBZO5rEM6KMEC95DBLJd9aKYDwwXdNpJwkwcOsBqD0o3
SOAl1akOmIU9VpkoffACCnw8dVXf1f3IpI8kN/gPaTEQOCaQOE3bfycZ4F6ANZ/r
oXOwpMsTKcrfH7TVIHKVnWB/7xemumaFc+j5s0SeN/BCpLpsVhXN6mpZ5jW8gZef
1MkQqSxzoyNBO+UvDUx7W6B2Fx5MJsJzC2I86kSMQkTpYc5zM2lgS7e+hurASOfw
lGd1gz+ixTyHawV7UxPDm9DafvyBVA2L5t0+y6SU3+7GNE66BnALTwfXTG85+pF6
+YmrHPDhMYAXYPQsgo9SM+magBb55WOwzSBk2LTEjaTZu61XStdVdrkP6eTLlX0I
ABvVzJCC8G57tZR263UacCH+PNuDAIQ8BZ7edHEAdE3wzprvbw5oHORWoL3kKZxH
nCoANBBN0EOm9oKivBlnekSBlqAAyvG5uoaTrUpBUrr++VNdV9cqcHXdmgGQVhhV
EBa3vNvKZwreMLtBWPGqYzUBesfb0QD/k6XvmRUzAFIEytvA3Lu9H0JPU9KJuGKt
HV8agQ5HKrXTJUIHfy9Ymq3jOEuSqIyfkO9c95VlkiHBPJNcsTlUmf6wMv7ncGmY
CEt4nZVgLtQDJQ91LXMZL9hAgsuaY+c3sNGzZTUyt7AzFpYDW7PzCRIqRBxV2/5K
8uld0CYbCFxMNV/i5FJRGZ5nCvF9uNNPxkgC1PEQGz1PGXB+Ns8J14+y5d/ftNUL
WwTGUAt+jgcQvSDHT7jwXYJPL/qlqfxswrwOep6Ykl36rPQ/z3S8rXVhk+EVgpZa
b0Bwe3bpsoLN8Pn/NgHFVPhAQ/t+F2sdZQN0DRJyyib8GknkVtRUBBxEf4gG6j9M
FjDJG6rJ0DugsqyANc7l+ZnTGhRNGb896Dn7vDhei6CW6vQuVfI52w6wakjNE3tv
9A1SCosHkHXCav88oohCwBbVQ2iBFxeajppSDV6awd0PKiJry9TUy9xeuqG94IBK
yaM2xlt27EKBCeW5rS5H4rPaHn8ONhYhAESjNrAcT9VAE2NEYuzq3ojSkwxmODWY
0FwDiBr8SCTA7RuyKEpzidZ3uo/tSxAeTjSVmaCVufkO/iVnyGsxxLOy3xsEXPx0
+InJ0lMaa13nRBzLUkxaHqMrjMwR1A/ivaIHQi1fkUxSm0s8MlLSiR2Q5gfxZJkH
+h+eCIHdzjC/TrXVovcyhLI55AZzUMKItLaMS5OLfS0YBT0JTH1yv2xT2aVAOQqN
sBXkekPI0CX/667xbu68k9CJVfu+KQj7UK9uiXTqtSqbPKI8V2a4eScz0gw5Fhus
UB6J3AI7xo0lN1qPAjFuFzafgfNDj1xmp+cZKP85si/6eA2qDbHepZRWWMZXbN4H
7VBnSW8lf0jpztddEm/q7dZVb3mc49k05teYu5HbhCiGzYqwUw1ViY+WgzrryHnU
Nw7BHvFa6Iuj4EF2ToUqDoBEP7Q0bq6YSaIGLmsukBB8jo9l8dUBaRN+xX1xbxgr
LsuyJx7U+Ys3c5u/Uq3idcYbizUzWQWhu/i8aTQk/2YfHWMTR6CgAAdZR0TtDk4Z
06uIMEGhC3IzK4tjxo2rItpGvXgoNqzxOiSbBEU9cHg79WLOJf2CRW9D2NsTfa7Q
Pxn8o98ljb+9beBb9Nxqx7KAIT5DGK7pr9RUOjOcg0Zm68DuwGC9eW5aQtkb2yPI
wCRMfQ8lv/fC7e9kX6e0pAZvdMxYt5/vNnAf4ZWa/RPc9ggMNFry8pabZIy8gq6E
GUkq4lKxXEVwj+yPDGEa7iLEEMcAl5wqHCB9L5Ah1JhwfbwdJZq1TDaajgOG++7n
BVRwuTSFCie7wVw10SOFlpcYFKGi8U/UpsUXm/i0NzRfJORH0i3wJII6w+vop0Td
FHA794EJ4ncYqMrHyOq2YicwKnx96o8yGtoE/CPsC/lpTxRnGst9c3D+YU4ukJ+u
Qi/Es0S4uFdKC9kbE+WboIpR8Agl5olT9DKUBvG3iwwN9AIrkE8NTwTSdB+USL1P
SkpcJleZ6cCgdWeBmoJdMSCV7T9XCrfLxXQGoC4c2A5Sc2wNVJ9kQrKkIlV6jmYM
LOFGF9BWT1VA7TtGM7cSZxPqxkHicGVFiUzR1njUUawrVUt+es5wnSGIu720h5bt
zKRxQHkAXqDvqD7nkT00kGIVvQVPIr0+PSy28qT/iBYHe7fJwf++pdgJsI/O29CE
XCqL18FChpT4Kiz3nza8pJMn75J+aw+N5YxrrAFFhI2ctNSC2a+WtWQBnckI66l+
3m+ftL81WL/63bgODl0KzBxeWb/PZ00qnm0vV4al8JTjNitpmgLw3YPqN1tprgFJ
GnrP9I8gfkdm1xmegrN5MtX4lfMJdn0Q/2aKT+gJJ28Nb29Vp3uS/rJAg9y5qjBM
iFXUTCX2qC6vjMmTqW/+VYQBgMETM3J17Pb3AOIY8qIlicHEp2+xGvzRgkj9Dtk7
9jQLIjYtZFf9OJG2i+oxlX3L6mBgPmy5Bmdmj0oeixF7UEylBAWdbg0Fb/nTd2f9
ehlg0GC3CxB6owVPWDFSdbmYjJ+cgu4w+ZqgRIaUTBGmbIcmLrOJFmOOmGZLBcRn
P7BF3Al+YoOTVxTE+ooHLJwN70fUcGChOMgE44w5h9miTXw7Ir6/UMKjTJqt2JiY
rRLvYWPpc1FiIMMhaOZeEgB5W9Tpk2wq7yMzAThdOCxGTJLnWcNNJnz+QerzhI9B
CfcqRZE40Fg7VaWvMUwYHrNPjpBfBAuFUnbTvbJj2AD//0H6MEiCwAi1lAtgQtyx
95jCSfRw3cDh9Cy5z8mkwqCsm3uXCuVHg5zvym3AQ21Arj2OBM0V8oudDLwpYROd
vRTGujaOYLwrEPv8E7bjKSUBzCS8btDdW6s8Vougb/dpNrtHbs9YltWskBuyyvwR
hV3bXYF2YtZItYlLn9PPe7Gq+OsLND7d+VRZyHbw1KeCPuCD8IUMJnmqQXx9+PGD
ii+NKjE9O7Tr02OINAictl8apjjzdgnnIZYWIzaHTfPlaxDUvJJXCU8uefQGA2r5
4MeZ5UPETgdqYS5MA/nWjmuv3CidsEZE+AS/EDab2iuoKSG6ez1DHIC/m6CGIEcn
+shNUg+jXnnEN5mcHYbA6KOhazqdAJkOkm27vug3hgkCgzNl7McylsbdW5/UT8ol
tYFmtEwwUgH+DZNPWZDaHkhWZd7g680H03i69NcJVzo8rdl3aK7HucFMhQQpgHQb
S3XNgAhHHFQvv9flGwRuQAd5wz1+HAexMq6CR/D5DtG+kj5ZLJkDXrvL4J7iC54M
gN0kerF+gIFE5JbdjmEpagioeq8t7plGgXThmq6AG6LFa3xc2AHMX6kYWhExPkZo
v1q0+Jm1fSVikprF52uOXqg1AMGHB2mr8fto7tiL6hmwqNQ7ahfxJ21d9ZnQxbQ8
IVZX8CD2a5lk7C7v2ohyiEWvQb6/LpidZ+/0Dsp+l9Se2N9tJHcin/PZUuXGyXDq
8bT+EjEmvDjFXpMbHQton60stGt5GgofotCiXYQHhB2BRfdK0U0ROVtAiRfYh9/4
OZAj+f57IrmoWQXLLS7c7Fzq5bs7oaH//QjQBzafaeJWs2tM6l0TKJBv6gzEAh5y
ILkkV7jsqN7AmZoU5KEIAsVDi99DGjsAJdqIEhh0S2/t4OOymBG5mWzD09WEe2Qc
f2Dy9vfPe1VWVgwMY7OoZkjGGfeQWu8I4V2c1tf9OZz3B6qEUkwtz/xO/5iXd8qP
WItQsuYiT4tgWqHBmAJ78DVHU04y9PGi8dLLU4L6fKBvUZmprmKI284h1HSQrG5j
wEG6WAA+TFhFEc37htyaAbuwF+sasVtni4iEKUx6jmsTUbOfKm2eLUtyiLM/hZed
2D+QqoLv2YfALnkBMuck26xyWaJeWBqEoSt0tY9L6CA=
`pragma protect end_protected
